module MockArray(
  input         clock,
  input         reset,
  input  [63:0] io_insHorizontal_0_0,
  input  [63:0] io_insHorizontal_0_1,
  input  [63:0] io_insHorizontal_0_2,
  input  [63:0] io_insHorizontal_0_3,
  input  [63:0] io_insHorizontal_0_4,
  input  [63:0] io_insHorizontal_0_5,
  input  [63:0] io_insHorizontal_0_6,
  input  [63:0] io_insHorizontal_0_7,
  input  [63:0] io_insHorizontal_0_8,
  input  [63:0] io_insHorizontal_0_9,
  input  [63:0] io_insHorizontal_0_10,
  input  [63:0] io_insHorizontal_0_11,
  input  [63:0] io_insHorizontal_0_12,
  input  [63:0] io_insHorizontal_0_13,
  input  [63:0] io_insHorizontal_0_14,
  input  [63:0] io_insHorizontal_0_15,
  input  [63:0] io_insHorizontal_0_16,
  input  [63:0] io_insHorizontal_0_17,
  input  [63:0] io_insHorizontal_0_18,
  input  [63:0] io_insHorizontal_0_19,
  input  [63:0] io_insHorizontal_0_20,
  input  [63:0] io_insHorizontal_0_21,
  input  [63:0] io_insHorizontal_0_22,
  input  [63:0] io_insHorizontal_0_23,
  input  [63:0] io_insHorizontal_0_24,
  input  [63:0] io_insHorizontal_0_25,
  input  [63:0] io_insHorizontal_0_26,
  input  [63:0] io_insHorizontal_0_27,
  input  [63:0] io_insHorizontal_0_28,
  input  [63:0] io_insHorizontal_0_29,
  input  [63:0] io_insHorizontal_0_30,
  input  [63:0] io_insHorizontal_0_31,
  input  [63:0] io_insHorizontal_1_0,
  input  [63:0] io_insHorizontal_1_1,
  input  [63:0] io_insHorizontal_1_2,
  input  [63:0] io_insHorizontal_1_3,
  input  [63:0] io_insHorizontal_1_4,
  input  [63:0] io_insHorizontal_1_5,
  input  [63:0] io_insHorizontal_1_6,
  input  [63:0] io_insHorizontal_1_7,
  input  [63:0] io_insHorizontal_1_8,
  input  [63:0] io_insHorizontal_1_9,
  input  [63:0] io_insHorizontal_1_10,
  input  [63:0] io_insHorizontal_1_11,
  input  [63:0] io_insHorizontal_1_12,
  input  [63:0] io_insHorizontal_1_13,
  input  [63:0] io_insHorizontal_1_14,
  input  [63:0] io_insHorizontal_1_15,
  input  [63:0] io_insHorizontal_1_16,
  input  [63:0] io_insHorizontal_1_17,
  input  [63:0] io_insHorizontal_1_18,
  input  [63:0] io_insHorizontal_1_19,
  input  [63:0] io_insHorizontal_1_20,
  input  [63:0] io_insHorizontal_1_21,
  input  [63:0] io_insHorizontal_1_22,
  input  [63:0] io_insHorizontal_1_23,
  input  [63:0] io_insHorizontal_1_24,
  input  [63:0] io_insHorizontal_1_25,
  input  [63:0] io_insHorizontal_1_26,
  input  [63:0] io_insHorizontal_1_27,
  input  [63:0] io_insHorizontal_1_28,
  input  [63:0] io_insHorizontal_1_29,
  input  [63:0] io_insHorizontal_1_30,
  input  [63:0] io_insHorizontal_1_31,
  output [63:0] io_outsHorizontal_0_0,
  output [63:0] io_outsHorizontal_0_1,
  output [63:0] io_outsHorizontal_0_2,
  output [63:0] io_outsHorizontal_0_3,
  output [63:0] io_outsHorizontal_0_4,
  output [63:0] io_outsHorizontal_0_5,
  output [63:0] io_outsHorizontal_0_6,
  output [63:0] io_outsHorizontal_0_7,
  output [63:0] io_outsHorizontal_0_8,
  output [63:0] io_outsHorizontal_0_9,
  output [63:0] io_outsHorizontal_0_10,
  output [63:0] io_outsHorizontal_0_11,
  output [63:0] io_outsHorizontal_0_12,
  output [63:0] io_outsHorizontal_0_13,
  output [63:0] io_outsHorizontal_0_14,
  output [63:0] io_outsHorizontal_0_15,
  output [63:0] io_outsHorizontal_0_16,
  output [63:0] io_outsHorizontal_0_17,
  output [63:0] io_outsHorizontal_0_18,
  output [63:0] io_outsHorizontal_0_19,
  output [63:0] io_outsHorizontal_0_20,
  output [63:0] io_outsHorizontal_0_21,
  output [63:0] io_outsHorizontal_0_22,
  output [63:0] io_outsHorizontal_0_23,
  output [63:0] io_outsHorizontal_0_24,
  output [63:0] io_outsHorizontal_0_25,
  output [63:0] io_outsHorizontal_0_26,
  output [63:0] io_outsHorizontal_0_27,
  output [63:0] io_outsHorizontal_0_28,
  output [63:0] io_outsHorizontal_0_29,
  output [63:0] io_outsHorizontal_0_30,
  output [63:0] io_outsHorizontal_0_31,
  output [63:0] io_outsHorizontal_1_0,
  output [63:0] io_outsHorizontal_1_1,
  output [63:0] io_outsHorizontal_1_2,
  output [63:0] io_outsHorizontal_1_3,
  output [63:0] io_outsHorizontal_1_4,
  output [63:0] io_outsHorizontal_1_5,
  output [63:0] io_outsHorizontal_1_6,
  output [63:0] io_outsHorizontal_1_7,
  output [63:0] io_outsHorizontal_1_8,
  output [63:0] io_outsHorizontal_1_9,
  output [63:0] io_outsHorizontal_1_10,
  output [63:0] io_outsHorizontal_1_11,
  output [63:0] io_outsHorizontal_1_12,
  output [63:0] io_outsHorizontal_1_13,
  output [63:0] io_outsHorizontal_1_14,
  output [63:0] io_outsHorizontal_1_15,
  output [63:0] io_outsHorizontal_1_16,
  output [63:0] io_outsHorizontal_1_17,
  output [63:0] io_outsHorizontal_1_18,
  output [63:0] io_outsHorizontal_1_19,
  output [63:0] io_outsHorizontal_1_20,
  output [63:0] io_outsHorizontal_1_21,
  output [63:0] io_outsHorizontal_1_22,
  output [63:0] io_outsHorizontal_1_23,
  output [63:0] io_outsHorizontal_1_24,
  output [63:0] io_outsHorizontal_1_25,
  output [63:0] io_outsHorizontal_1_26,
  output [63:0] io_outsHorizontal_1_27,
  output [63:0] io_outsHorizontal_1_28,
  output [63:0] io_outsHorizontal_1_29,
  output [63:0] io_outsHorizontal_1_30,
  output [63:0] io_outsHorizontal_1_31,
  input  [63:0] io_insVertical_0_0,
  input  [63:0] io_insVertical_0_1,
  input  [63:0] io_insVertical_0_2,
  input  [63:0] io_insVertical_0_3,
  input  [63:0] io_insVertical_0_4,
  input  [63:0] io_insVertical_0_5,
  input  [63:0] io_insVertical_0_6,
  input  [63:0] io_insVertical_0_7,
  input  [63:0] io_insVertical_0_8,
  input  [63:0] io_insVertical_0_9,
  input  [63:0] io_insVertical_0_10,
  input  [63:0] io_insVertical_0_11,
  input  [63:0] io_insVertical_0_12,
  input  [63:0] io_insVertical_0_13,
  input  [63:0] io_insVertical_0_14,
  input  [63:0] io_insVertical_0_15,
  input  [63:0] io_insVertical_0_16,
  input  [63:0] io_insVertical_0_17,
  input  [63:0] io_insVertical_0_18,
  input  [63:0] io_insVertical_0_19,
  input  [63:0] io_insVertical_0_20,
  input  [63:0] io_insVertical_0_21,
  input  [63:0] io_insVertical_0_22,
  input  [63:0] io_insVertical_0_23,
  input  [63:0] io_insVertical_0_24,
  input  [63:0] io_insVertical_0_25,
  input  [63:0] io_insVertical_0_26,
  input  [63:0] io_insVertical_0_27,
  input  [63:0] io_insVertical_0_28,
  input  [63:0] io_insVertical_0_29,
  input  [63:0] io_insVertical_0_30,
  input  [63:0] io_insVertical_0_31,
  input  [63:0] io_insVertical_1_0,
  input  [63:0] io_insVertical_1_1,
  input  [63:0] io_insVertical_1_2,
  input  [63:0] io_insVertical_1_3,
  input  [63:0] io_insVertical_1_4,
  input  [63:0] io_insVertical_1_5,
  input  [63:0] io_insVertical_1_6,
  input  [63:0] io_insVertical_1_7,
  input  [63:0] io_insVertical_1_8,
  input  [63:0] io_insVertical_1_9,
  input  [63:0] io_insVertical_1_10,
  input  [63:0] io_insVertical_1_11,
  input  [63:0] io_insVertical_1_12,
  input  [63:0] io_insVertical_1_13,
  input  [63:0] io_insVertical_1_14,
  input  [63:0] io_insVertical_1_15,
  input  [63:0] io_insVertical_1_16,
  input  [63:0] io_insVertical_1_17,
  input  [63:0] io_insVertical_1_18,
  input  [63:0] io_insVertical_1_19,
  input  [63:0] io_insVertical_1_20,
  input  [63:0] io_insVertical_1_21,
  input  [63:0] io_insVertical_1_22,
  input  [63:0] io_insVertical_1_23,
  input  [63:0] io_insVertical_1_24,
  input  [63:0] io_insVertical_1_25,
  input  [63:0] io_insVertical_1_26,
  input  [63:0] io_insVertical_1_27,
  input  [63:0] io_insVertical_1_28,
  input  [63:0] io_insVertical_1_29,
  input  [63:0] io_insVertical_1_30,
  input  [63:0] io_insVertical_1_31,
  output [63:0] io_outsVertical_0_0,
  output [63:0] io_outsVertical_0_1,
  output [63:0] io_outsVertical_0_2,
  output [63:0] io_outsVertical_0_3,
  output [63:0] io_outsVertical_0_4,
  output [63:0] io_outsVertical_0_5,
  output [63:0] io_outsVertical_0_6,
  output [63:0] io_outsVertical_0_7,
  output [63:0] io_outsVertical_0_8,
  output [63:0] io_outsVertical_0_9,
  output [63:0] io_outsVertical_0_10,
  output [63:0] io_outsVertical_0_11,
  output [63:0] io_outsVertical_0_12,
  output [63:0] io_outsVertical_0_13,
  output [63:0] io_outsVertical_0_14,
  output [63:0] io_outsVertical_0_15,
  output [63:0] io_outsVertical_0_16,
  output [63:0] io_outsVertical_0_17,
  output [63:0] io_outsVertical_0_18,
  output [63:0] io_outsVertical_0_19,
  output [63:0] io_outsVertical_0_20,
  output [63:0] io_outsVertical_0_21,
  output [63:0] io_outsVertical_0_22,
  output [63:0] io_outsVertical_0_23,
  output [63:0] io_outsVertical_0_24,
  output [63:0] io_outsVertical_0_25,
  output [63:0] io_outsVertical_0_26,
  output [63:0] io_outsVertical_0_27,
  output [63:0] io_outsVertical_0_28,
  output [63:0] io_outsVertical_0_29,
  output [63:0] io_outsVertical_0_30,
  output [63:0] io_outsVertical_0_31,
  output [63:0] io_outsVertical_1_0,
  output [63:0] io_outsVertical_1_1,
  output [63:0] io_outsVertical_1_2,
  output [63:0] io_outsVertical_1_3,
  output [63:0] io_outsVertical_1_4,
  output [63:0] io_outsVertical_1_5,
  output [63:0] io_outsVertical_1_6,
  output [63:0] io_outsVertical_1_7,
  output [63:0] io_outsVertical_1_8,
  output [63:0] io_outsVertical_1_9,
  output [63:0] io_outsVertical_1_10,
  output [63:0] io_outsVertical_1_11,
  output [63:0] io_outsVertical_1_12,
  output [63:0] io_outsVertical_1_13,
  output [63:0] io_outsVertical_1_14,
  output [63:0] io_outsVertical_1_15,
  output [63:0] io_outsVertical_1_16,
  output [63:0] io_outsVertical_1_17,
  output [63:0] io_outsVertical_1_18,
  output [63:0] io_outsVertical_1_19,
  output [63:0] io_outsVertical_1_20,
  output [63:0] io_outsVertical_1_21,
  output [63:0] io_outsVertical_1_22,
  output [63:0] io_outsVertical_1_23,
  output [63:0] io_outsVertical_1_24,
  output [63:0] io_outsVertical_1_25,
  output [63:0] io_outsVertical_1_26,
  output [63:0] io_outsVertical_1_27,
  output [63:0] io_outsVertical_1_28,
  output [63:0] io_outsVertical_1_29,
  output [63:0] io_outsVertical_1_30,
  output [63:0] io_outsVertical_1_31,
  output        io_lsbs_0,
  output        io_lsbs_1,
  output        io_lsbs_2,
  output        io_lsbs_3,
  output        io_lsbs_4,
  output        io_lsbs_5,
  output        io_lsbs_6,
  output        io_lsbs_7,
  output        io_lsbs_8,
  output        io_lsbs_9,
  output        io_lsbs_10,
  output        io_lsbs_11,
  output        io_lsbs_12,
  output        io_lsbs_13,
  output        io_lsbs_14,
  output        io_lsbs_15,
  output        io_lsbs_16,
  output        io_lsbs_17,
  output        io_lsbs_18,
  output        io_lsbs_19,
  output        io_lsbs_20,
  output        io_lsbs_21,
  output        io_lsbs_22,
  output        io_lsbs_23,
  output        io_lsbs_24,
  output        io_lsbs_25,
  output        io_lsbs_26,
  output        io_lsbs_27,
  output        io_lsbs_28,
  output        io_lsbs_29,
  output        io_lsbs_30,
  output        io_lsbs_31,
  output        io_lsbs_32,
  output        io_lsbs_33,
  output        io_lsbs_34,
  output        io_lsbs_35,
  output        io_lsbs_36,
  output        io_lsbs_37,
  output        io_lsbs_38,
  output        io_lsbs_39,
  output        io_lsbs_40,
  output        io_lsbs_41,
  output        io_lsbs_42,
  output        io_lsbs_43,
  output        io_lsbs_44,
  output        io_lsbs_45,
  output        io_lsbs_46,
  output        io_lsbs_47,
  output        io_lsbs_48,
  output        io_lsbs_49,
  output        io_lsbs_50,
  output        io_lsbs_51,
  output        io_lsbs_52,
  output        io_lsbs_53,
  output        io_lsbs_54,
  output        io_lsbs_55,
  output        io_lsbs_56,
  output        io_lsbs_57,
  output        io_lsbs_58,
  output        io_lsbs_59,
  output        io_lsbs_60,
  output        io_lsbs_61,
  output        io_lsbs_62,
  output        io_lsbs_63,
  output        io_lsbs_64,
  output        io_lsbs_65,
  output        io_lsbs_66,
  output        io_lsbs_67,
  output        io_lsbs_68,
  output        io_lsbs_69,
  output        io_lsbs_70,
  output        io_lsbs_71,
  output        io_lsbs_72,
  output        io_lsbs_73,
  output        io_lsbs_74,
  output        io_lsbs_75,
  output        io_lsbs_76,
  output        io_lsbs_77,
  output        io_lsbs_78,
  output        io_lsbs_79,
  output        io_lsbs_80,
  output        io_lsbs_81,
  output        io_lsbs_82,
  output        io_lsbs_83,
  output        io_lsbs_84,
  output        io_lsbs_85,
  output        io_lsbs_86,
  output        io_lsbs_87,
  output        io_lsbs_88,
  output        io_lsbs_89,
  output        io_lsbs_90,
  output        io_lsbs_91,
  output        io_lsbs_92,
  output        io_lsbs_93,
  output        io_lsbs_94,
  output        io_lsbs_95,
  output        io_lsbs_96,
  output        io_lsbs_97,
  output        io_lsbs_98,
  output        io_lsbs_99,
  output        io_lsbs_100,
  output        io_lsbs_101,
  output        io_lsbs_102,
  output        io_lsbs_103,
  output        io_lsbs_104,
  output        io_lsbs_105,
  output        io_lsbs_106,
  output        io_lsbs_107,
  output        io_lsbs_108,
  output        io_lsbs_109,
  output        io_lsbs_110,
  output        io_lsbs_111,
  output        io_lsbs_112,
  output        io_lsbs_113,
  output        io_lsbs_114,
  output        io_lsbs_115,
  output        io_lsbs_116,
  output        io_lsbs_117,
  output        io_lsbs_118,
  output        io_lsbs_119,
  output        io_lsbs_120,
  output        io_lsbs_121,
  output        io_lsbs_122,
  output        io_lsbs_123,
  output        io_lsbs_124,
  output        io_lsbs_125,
  output        io_lsbs_126,
  output        io_lsbs_127,
  output        io_lsbs_128,
  output        io_lsbs_129,
  output        io_lsbs_130,
  output        io_lsbs_131,
  output        io_lsbs_132,
  output        io_lsbs_133,
  output        io_lsbs_134,
  output        io_lsbs_135,
  output        io_lsbs_136,
  output        io_lsbs_137,
  output        io_lsbs_138,
  output        io_lsbs_139,
  output        io_lsbs_140,
  output        io_lsbs_141,
  output        io_lsbs_142,
  output        io_lsbs_143,
  output        io_lsbs_144,
  output        io_lsbs_145,
  output        io_lsbs_146,
  output        io_lsbs_147,
  output        io_lsbs_148,
  output        io_lsbs_149,
  output        io_lsbs_150,
  output        io_lsbs_151,
  output        io_lsbs_152,
  output        io_lsbs_153,
  output        io_lsbs_154,
  output        io_lsbs_155,
  output        io_lsbs_156,
  output        io_lsbs_157,
  output        io_lsbs_158,
  output        io_lsbs_159,
  output        io_lsbs_160,
  output        io_lsbs_161,
  output        io_lsbs_162,
  output        io_lsbs_163,
  output        io_lsbs_164,
  output        io_lsbs_165,
  output        io_lsbs_166,
  output        io_lsbs_167,
  output        io_lsbs_168,
  output        io_lsbs_169,
  output        io_lsbs_170,
  output        io_lsbs_171,
  output        io_lsbs_172,
  output        io_lsbs_173,
  output        io_lsbs_174,
  output        io_lsbs_175,
  output        io_lsbs_176,
  output        io_lsbs_177,
  output        io_lsbs_178,
  output        io_lsbs_179,
  output        io_lsbs_180,
  output        io_lsbs_181,
  output        io_lsbs_182,
  output        io_lsbs_183,
  output        io_lsbs_184,
  output        io_lsbs_185,
  output        io_lsbs_186,
  output        io_lsbs_187,
  output        io_lsbs_188,
  output        io_lsbs_189,
  output        io_lsbs_190,
  output        io_lsbs_191,
  output        io_lsbs_192,
  output        io_lsbs_193,
  output        io_lsbs_194,
  output        io_lsbs_195,
  output        io_lsbs_196,
  output        io_lsbs_197,
  output        io_lsbs_198,
  output        io_lsbs_199,
  output        io_lsbs_200,
  output        io_lsbs_201,
  output        io_lsbs_202,
  output        io_lsbs_203,
  output        io_lsbs_204,
  output        io_lsbs_205,
  output        io_lsbs_206,
  output        io_lsbs_207,
  output        io_lsbs_208,
  output        io_lsbs_209,
  output        io_lsbs_210,
  output        io_lsbs_211,
  output        io_lsbs_212,
  output        io_lsbs_213,
  output        io_lsbs_214,
  output        io_lsbs_215,
  output        io_lsbs_216,
  output        io_lsbs_217,
  output        io_lsbs_218,
  output        io_lsbs_219,
  output        io_lsbs_220,
  output        io_lsbs_221,
  output        io_lsbs_222,
  output        io_lsbs_223,
  output        io_lsbs_224,
  output        io_lsbs_225,
  output        io_lsbs_226,
  output        io_lsbs_227,
  output        io_lsbs_228,
  output        io_lsbs_229,
  output        io_lsbs_230,
  output        io_lsbs_231,
  output        io_lsbs_232,
  output        io_lsbs_233,
  output        io_lsbs_234,
  output        io_lsbs_235,
  output        io_lsbs_236,
  output        io_lsbs_237,
  output        io_lsbs_238,
  output        io_lsbs_239,
  output        io_lsbs_240,
  output        io_lsbs_241,
  output        io_lsbs_242,
  output        io_lsbs_243,
  output        io_lsbs_244,
  output        io_lsbs_245,
  output        io_lsbs_246,
  output        io_lsbs_247,
  output        io_lsbs_248,
  output        io_lsbs_249,
  output        io_lsbs_250,
  output        io_lsbs_251,
  output        io_lsbs_252,
  output        io_lsbs_253,
  output        io_lsbs_254,
  output        io_lsbs_255,
  output        io_lsbs_256,
  output        io_lsbs_257,
  output        io_lsbs_258,
  output        io_lsbs_259,
  output        io_lsbs_260,
  output        io_lsbs_261,
  output        io_lsbs_262,
  output        io_lsbs_263,
  output        io_lsbs_264,
  output        io_lsbs_265,
  output        io_lsbs_266,
  output        io_lsbs_267,
  output        io_lsbs_268,
  output        io_lsbs_269,
  output        io_lsbs_270,
  output        io_lsbs_271,
  output        io_lsbs_272,
  output        io_lsbs_273,
  output        io_lsbs_274,
  output        io_lsbs_275,
  output        io_lsbs_276,
  output        io_lsbs_277,
  output        io_lsbs_278,
  output        io_lsbs_279,
  output        io_lsbs_280,
  output        io_lsbs_281,
  output        io_lsbs_282,
  output        io_lsbs_283,
  output        io_lsbs_284,
  output        io_lsbs_285,
  output        io_lsbs_286,
  output        io_lsbs_287,
  output        io_lsbs_288,
  output        io_lsbs_289,
  output        io_lsbs_290,
  output        io_lsbs_291,
  output        io_lsbs_292,
  output        io_lsbs_293,
  output        io_lsbs_294,
  output        io_lsbs_295,
  output        io_lsbs_296,
  output        io_lsbs_297,
  output        io_lsbs_298,
  output        io_lsbs_299,
  output        io_lsbs_300,
  output        io_lsbs_301,
  output        io_lsbs_302,
  output        io_lsbs_303,
  output        io_lsbs_304,
  output        io_lsbs_305,
  output        io_lsbs_306,
  output        io_lsbs_307,
  output        io_lsbs_308,
  output        io_lsbs_309,
  output        io_lsbs_310,
  output        io_lsbs_311,
  output        io_lsbs_312,
  output        io_lsbs_313,
  output        io_lsbs_314,
  output        io_lsbs_315,
  output        io_lsbs_316,
  output        io_lsbs_317,
  output        io_lsbs_318,
  output        io_lsbs_319,
  output        io_lsbs_320,
  output        io_lsbs_321,
  output        io_lsbs_322,
  output        io_lsbs_323,
  output        io_lsbs_324,
  output        io_lsbs_325,
  output        io_lsbs_326,
  output        io_lsbs_327,
  output        io_lsbs_328,
  output        io_lsbs_329,
  output        io_lsbs_330,
  output        io_lsbs_331,
  output        io_lsbs_332,
  output        io_lsbs_333,
  output        io_lsbs_334,
  output        io_lsbs_335,
  output        io_lsbs_336,
  output        io_lsbs_337,
  output        io_lsbs_338,
  output        io_lsbs_339,
  output        io_lsbs_340,
  output        io_lsbs_341,
  output        io_lsbs_342,
  output        io_lsbs_343,
  output        io_lsbs_344,
  output        io_lsbs_345,
  output        io_lsbs_346,
  output        io_lsbs_347,
  output        io_lsbs_348,
  output        io_lsbs_349,
  output        io_lsbs_350,
  output        io_lsbs_351,
  output        io_lsbs_352,
  output        io_lsbs_353,
  output        io_lsbs_354,
  output        io_lsbs_355,
  output        io_lsbs_356,
  output        io_lsbs_357,
  output        io_lsbs_358,
  output        io_lsbs_359,
  output        io_lsbs_360,
  output        io_lsbs_361,
  output        io_lsbs_362,
  output        io_lsbs_363,
  output        io_lsbs_364,
  output        io_lsbs_365,
  output        io_lsbs_366,
  output        io_lsbs_367,
  output        io_lsbs_368,
  output        io_lsbs_369,
  output        io_lsbs_370,
  output        io_lsbs_371,
  output        io_lsbs_372,
  output        io_lsbs_373,
  output        io_lsbs_374,
  output        io_lsbs_375,
  output        io_lsbs_376,
  output        io_lsbs_377,
  output        io_lsbs_378,
  output        io_lsbs_379,
  output        io_lsbs_380,
  output        io_lsbs_381,
  output        io_lsbs_382,
  output        io_lsbs_383,
  output        io_lsbs_384,
  output        io_lsbs_385,
  output        io_lsbs_386,
  output        io_lsbs_387,
  output        io_lsbs_388,
  output        io_lsbs_389,
  output        io_lsbs_390,
  output        io_lsbs_391,
  output        io_lsbs_392,
  output        io_lsbs_393,
  output        io_lsbs_394,
  output        io_lsbs_395,
  output        io_lsbs_396,
  output        io_lsbs_397,
  output        io_lsbs_398,
  output        io_lsbs_399,
  output        io_lsbs_400,
  output        io_lsbs_401,
  output        io_lsbs_402,
  output        io_lsbs_403,
  output        io_lsbs_404,
  output        io_lsbs_405,
  output        io_lsbs_406,
  output        io_lsbs_407,
  output        io_lsbs_408,
  output        io_lsbs_409,
  output        io_lsbs_410,
  output        io_lsbs_411,
  output        io_lsbs_412,
  output        io_lsbs_413,
  output        io_lsbs_414,
  output        io_lsbs_415,
  output        io_lsbs_416,
  output        io_lsbs_417,
  output        io_lsbs_418,
  output        io_lsbs_419,
  output        io_lsbs_420,
  output        io_lsbs_421,
  output        io_lsbs_422,
  output        io_lsbs_423,
  output        io_lsbs_424,
  output        io_lsbs_425,
  output        io_lsbs_426,
  output        io_lsbs_427,
  output        io_lsbs_428,
  output        io_lsbs_429,
  output        io_lsbs_430,
  output        io_lsbs_431,
  output        io_lsbs_432,
  output        io_lsbs_433,
  output        io_lsbs_434,
  output        io_lsbs_435,
  output        io_lsbs_436,
  output        io_lsbs_437,
  output        io_lsbs_438,
  output        io_lsbs_439,
  output        io_lsbs_440,
  output        io_lsbs_441,
  output        io_lsbs_442,
  output        io_lsbs_443,
  output        io_lsbs_444,
  output        io_lsbs_445,
  output        io_lsbs_446,
  output        io_lsbs_447,
  output        io_lsbs_448,
  output        io_lsbs_449,
  output        io_lsbs_450,
  output        io_lsbs_451,
  output        io_lsbs_452,
  output        io_lsbs_453,
  output        io_lsbs_454,
  output        io_lsbs_455,
  output        io_lsbs_456,
  output        io_lsbs_457,
  output        io_lsbs_458,
  output        io_lsbs_459,
  output        io_lsbs_460,
  output        io_lsbs_461,
  output        io_lsbs_462,
  output        io_lsbs_463,
  output        io_lsbs_464,
  output        io_lsbs_465,
  output        io_lsbs_466,
  output        io_lsbs_467,
  output        io_lsbs_468,
  output        io_lsbs_469,
  output        io_lsbs_470,
  output        io_lsbs_471,
  output        io_lsbs_472,
  output        io_lsbs_473,
  output        io_lsbs_474,
  output        io_lsbs_475,
  output        io_lsbs_476,
  output        io_lsbs_477,
  output        io_lsbs_478,
  output        io_lsbs_479,
  output        io_lsbs_480,
  output        io_lsbs_481,
  output        io_lsbs_482,
  output        io_lsbs_483,
  output        io_lsbs_484,
  output        io_lsbs_485,
  output        io_lsbs_486,
  output        io_lsbs_487,
  output        io_lsbs_488,
  output        io_lsbs_489,
  output        io_lsbs_490,
  output        io_lsbs_491,
  output        io_lsbs_492,
  output        io_lsbs_493,
  output        io_lsbs_494,
  output        io_lsbs_495,
  output        io_lsbs_496,
  output        io_lsbs_497,
  output        io_lsbs_498,
  output        io_lsbs_499,
  output        io_lsbs_500,
  output        io_lsbs_501,
  output        io_lsbs_502,
  output        io_lsbs_503,
  output        io_lsbs_504,
  output        io_lsbs_505,
  output        io_lsbs_506,
  output        io_lsbs_507,
  output        io_lsbs_508,
  output        io_lsbs_509,
  output        io_lsbs_510,
  output        io_lsbs_511,
  output        io_lsbs_512,
  output        io_lsbs_513,
  output        io_lsbs_514,
  output        io_lsbs_515,
  output        io_lsbs_516,
  output        io_lsbs_517,
  output        io_lsbs_518,
  output        io_lsbs_519,
  output        io_lsbs_520,
  output        io_lsbs_521,
  output        io_lsbs_522,
  output        io_lsbs_523,
  output        io_lsbs_524,
  output        io_lsbs_525,
  output        io_lsbs_526,
  output        io_lsbs_527,
  output        io_lsbs_528,
  output        io_lsbs_529,
  output        io_lsbs_530,
  output        io_lsbs_531,
  output        io_lsbs_532,
  output        io_lsbs_533,
  output        io_lsbs_534,
  output        io_lsbs_535,
  output        io_lsbs_536,
  output        io_lsbs_537,
  output        io_lsbs_538,
  output        io_lsbs_539,
  output        io_lsbs_540,
  output        io_lsbs_541,
  output        io_lsbs_542,
  output        io_lsbs_543,
  output        io_lsbs_544,
  output        io_lsbs_545,
  output        io_lsbs_546,
  output        io_lsbs_547,
  output        io_lsbs_548,
  output        io_lsbs_549,
  output        io_lsbs_550,
  output        io_lsbs_551,
  output        io_lsbs_552,
  output        io_lsbs_553,
  output        io_lsbs_554,
  output        io_lsbs_555,
  output        io_lsbs_556,
  output        io_lsbs_557,
  output        io_lsbs_558,
  output        io_lsbs_559,
  output        io_lsbs_560,
  output        io_lsbs_561,
  output        io_lsbs_562,
  output        io_lsbs_563,
  output        io_lsbs_564,
  output        io_lsbs_565,
  output        io_lsbs_566,
  output        io_lsbs_567,
  output        io_lsbs_568,
  output        io_lsbs_569,
  output        io_lsbs_570,
  output        io_lsbs_571,
  output        io_lsbs_572,
  output        io_lsbs_573,
  output        io_lsbs_574,
  output        io_lsbs_575,
  output        io_lsbs_576,
  output        io_lsbs_577,
  output        io_lsbs_578,
  output        io_lsbs_579,
  output        io_lsbs_580,
  output        io_lsbs_581,
  output        io_lsbs_582,
  output        io_lsbs_583,
  output        io_lsbs_584,
  output        io_lsbs_585,
  output        io_lsbs_586,
  output        io_lsbs_587,
  output        io_lsbs_588,
  output        io_lsbs_589,
  output        io_lsbs_590,
  output        io_lsbs_591,
  output        io_lsbs_592,
  output        io_lsbs_593,
  output        io_lsbs_594,
  output        io_lsbs_595,
  output        io_lsbs_596,
  output        io_lsbs_597,
  output        io_lsbs_598,
  output        io_lsbs_599,
  output        io_lsbs_600,
  output        io_lsbs_601,
  output        io_lsbs_602,
  output        io_lsbs_603,
  output        io_lsbs_604,
  output        io_lsbs_605,
  output        io_lsbs_606,
  output        io_lsbs_607,
  output        io_lsbs_608,
  output        io_lsbs_609,
  output        io_lsbs_610,
  output        io_lsbs_611,
  output        io_lsbs_612,
  output        io_lsbs_613,
  output        io_lsbs_614,
  output        io_lsbs_615,
  output        io_lsbs_616,
  output        io_lsbs_617,
  output        io_lsbs_618,
  output        io_lsbs_619,
  output        io_lsbs_620,
  output        io_lsbs_621,
  output        io_lsbs_622,
  output        io_lsbs_623,
  output        io_lsbs_624,
  output        io_lsbs_625,
  output        io_lsbs_626,
  output        io_lsbs_627,
  output        io_lsbs_628,
  output        io_lsbs_629,
  output        io_lsbs_630,
  output        io_lsbs_631,
  output        io_lsbs_632,
  output        io_lsbs_633,
  output        io_lsbs_634,
  output        io_lsbs_635,
  output        io_lsbs_636,
  output        io_lsbs_637,
  output        io_lsbs_638,
  output        io_lsbs_639,
  output        io_lsbs_640,
  output        io_lsbs_641,
  output        io_lsbs_642,
  output        io_lsbs_643,
  output        io_lsbs_644,
  output        io_lsbs_645,
  output        io_lsbs_646,
  output        io_lsbs_647,
  output        io_lsbs_648,
  output        io_lsbs_649,
  output        io_lsbs_650,
  output        io_lsbs_651,
  output        io_lsbs_652,
  output        io_lsbs_653,
  output        io_lsbs_654,
  output        io_lsbs_655,
  output        io_lsbs_656,
  output        io_lsbs_657,
  output        io_lsbs_658,
  output        io_lsbs_659,
  output        io_lsbs_660,
  output        io_lsbs_661,
  output        io_lsbs_662,
  output        io_lsbs_663,
  output        io_lsbs_664,
  output        io_lsbs_665,
  output        io_lsbs_666,
  output        io_lsbs_667,
  output        io_lsbs_668,
  output        io_lsbs_669,
  output        io_lsbs_670,
  output        io_lsbs_671,
  output        io_lsbs_672,
  output        io_lsbs_673,
  output        io_lsbs_674,
  output        io_lsbs_675,
  output        io_lsbs_676,
  output        io_lsbs_677,
  output        io_lsbs_678,
  output        io_lsbs_679,
  output        io_lsbs_680,
  output        io_lsbs_681,
  output        io_lsbs_682,
  output        io_lsbs_683,
  output        io_lsbs_684,
  output        io_lsbs_685,
  output        io_lsbs_686,
  output        io_lsbs_687,
  output        io_lsbs_688,
  output        io_lsbs_689,
  output        io_lsbs_690,
  output        io_lsbs_691,
  output        io_lsbs_692,
  output        io_lsbs_693,
  output        io_lsbs_694,
  output        io_lsbs_695,
  output        io_lsbs_696,
  output        io_lsbs_697,
  output        io_lsbs_698,
  output        io_lsbs_699,
  output        io_lsbs_700,
  output        io_lsbs_701,
  output        io_lsbs_702,
  output        io_lsbs_703,
  output        io_lsbs_704,
  output        io_lsbs_705,
  output        io_lsbs_706,
  output        io_lsbs_707,
  output        io_lsbs_708,
  output        io_lsbs_709,
  output        io_lsbs_710,
  output        io_lsbs_711,
  output        io_lsbs_712,
  output        io_lsbs_713,
  output        io_lsbs_714,
  output        io_lsbs_715,
  output        io_lsbs_716,
  output        io_lsbs_717,
  output        io_lsbs_718,
  output        io_lsbs_719,
  output        io_lsbs_720,
  output        io_lsbs_721,
  output        io_lsbs_722,
  output        io_lsbs_723,
  output        io_lsbs_724,
  output        io_lsbs_725,
  output        io_lsbs_726,
  output        io_lsbs_727,
  output        io_lsbs_728,
  output        io_lsbs_729,
  output        io_lsbs_730,
  output        io_lsbs_731,
  output        io_lsbs_732,
  output        io_lsbs_733,
  output        io_lsbs_734,
  output        io_lsbs_735,
  output        io_lsbs_736,
  output        io_lsbs_737,
  output        io_lsbs_738,
  output        io_lsbs_739,
  output        io_lsbs_740,
  output        io_lsbs_741,
  output        io_lsbs_742,
  output        io_lsbs_743,
  output        io_lsbs_744,
  output        io_lsbs_745,
  output        io_lsbs_746,
  output        io_lsbs_747,
  output        io_lsbs_748,
  output        io_lsbs_749,
  output        io_lsbs_750,
  output        io_lsbs_751,
  output        io_lsbs_752,
  output        io_lsbs_753,
  output        io_lsbs_754,
  output        io_lsbs_755,
  output        io_lsbs_756,
  output        io_lsbs_757,
  output        io_lsbs_758,
  output        io_lsbs_759,
  output        io_lsbs_760,
  output        io_lsbs_761,
  output        io_lsbs_762,
  output        io_lsbs_763,
  output        io_lsbs_764,
  output        io_lsbs_765,
  output        io_lsbs_766,
  output        io_lsbs_767,
  output        io_lsbs_768,
  output        io_lsbs_769,
  output        io_lsbs_770,
  output        io_lsbs_771,
  output        io_lsbs_772,
  output        io_lsbs_773,
  output        io_lsbs_774,
  output        io_lsbs_775,
  output        io_lsbs_776,
  output        io_lsbs_777,
  output        io_lsbs_778,
  output        io_lsbs_779,
  output        io_lsbs_780,
  output        io_lsbs_781,
  output        io_lsbs_782,
  output        io_lsbs_783,
  output        io_lsbs_784,
  output        io_lsbs_785,
  output        io_lsbs_786,
  output        io_lsbs_787,
  output        io_lsbs_788,
  output        io_lsbs_789,
  output        io_lsbs_790,
  output        io_lsbs_791,
  output        io_lsbs_792,
  output        io_lsbs_793,
  output        io_lsbs_794,
  output        io_lsbs_795,
  output        io_lsbs_796,
  output        io_lsbs_797,
  output        io_lsbs_798,
  output        io_lsbs_799,
  output        io_lsbs_800,
  output        io_lsbs_801,
  output        io_lsbs_802,
  output        io_lsbs_803,
  output        io_lsbs_804,
  output        io_lsbs_805,
  output        io_lsbs_806,
  output        io_lsbs_807,
  output        io_lsbs_808,
  output        io_lsbs_809,
  output        io_lsbs_810,
  output        io_lsbs_811,
  output        io_lsbs_812,
  output        io_lsbs_813,
  output        io_lsbs_814,
  output        io_lsbs_815,
  output        io_lsbs_816,
  output        io_lsbs_817,
  output        io_lsbs_818,
  output        io_lsbs_819,
  output        io_lsbs_820,
  output        io_lsbs_821,
  output        io_lsbs_822,
  output        io_lsbs_823,
  output        io_lsbs_824,
  output        io_lsbs_825,
  output        io_lsbs_826,
  output        io_lsbs_827,
  output        io_lsbs_828,
  output        io_lsbs_829,
  output        io_lsbs_830,
  output        io_lsbs_831,
  output        io_lsbs_832,
  output        io_lsbs_833,
  output        io_lsbs_834,
  output        io_lsbs_835,
  output        io_lsbs_836,
  output        io_lsbs_837,
  output        io_lsbs_838,
  output        io_lsbs_839,
  output        io_lsbs_840,
  output        io_lsbs_841,
  output        io_lsbs_842,
  output        io_lsbs_843,
  output        io_lsbs_844,
  output        io_lsbs_845,
  output        io_lsbs_846,
  output        io_lsbs_847,
  output        io_lsbs_848,
  output        io_lsbs_849,
  output        io_lsbs_850,
  output        io_lsbs_851,
  output        io_lsbs_852,
  output        io_lsbs_853,
  output        io_lsbs_854,
  output        io_lsbs_855,
  output        io_lsbs_856,
  output        io_lsbs_857,
  output        io_lsbs_858,
  output        io_lsbs_859,
  output        io_lsbs_860,
  output        io_lsbs_861,
  output        io_lsbs_862,
  output        io_lsbs_863,
  output        io_lsbs_864,
  output        io_lsbs_865,
  output        io_lsbs_866,
  output        io_lsbs_867,
  output        io_lsbs_868,
  output        io_lsbs_869,
  output        io_lsbs_870,
  output        io_lsbs_871,
  output        io_lsbs_872,
  output        io_lsbs_873,
  output        io_lsbs_874,
  output        io_lsbs_875,
  output        io_lsbs_876,
  output        io_lsbs_877,
  output        io_lsbs_878,
  output        io_lsbs_879,
  output        io_lsbs_880,
  output        io_lsbs_881,
  output        io_lsbs_882,
  output        io_lsbs_883,
  output        io_lsbs_884,
  output        io_lsbs_885,
  output        io_lsbs_886,
  output        io_lsbs_887,
  output        io_lsbs_888,
  output        io_lsbs_889,
  output        io_lsbs_890,
  output        io_lsbs_891,
  output        io_lsbs_892,
  output        io_lsbs_893,
  output        io_lsbs_894,
  output        io_lsbs_895,
  output        io_lsbs_896,
  output        io_lsbs_897,
  output        io_lsbs_898,
  output        io_lsbs_899,
  output        io_lsbs_900,
  output        io_lsbs_901,
  output        io_lsbs_902,
  output        io_lsbs_903,
  output        io_lsbs_904,
  output        io_lsbs_905,
  output        io_lsbs_906,
  output        io_lsbs_907,
  output        io_lsbs_908,
  output        io_lsbs_909,
  output        io_lsbs_910,
  output        io_lsbs_911,
  output        io_lsbs_912,
  output        io_lsbs_913,
  output        io_lsbs_914,
  output        io_lsbs_915,
  output        io_lsbs_916,
  output        io_lsbs_917,
  output        io_lsbs_918,
  output        io_lsbs_919,
  output        io_lsbs_920,
  output        io_lsbs_921,
  output        io_lsbs_922,
  output        io_lsbs_923,
  output        io_lsbs_924,
  output        io_lsbs_925,
  output        io_lsbs_926,
  output        io_lsbs_927,
  output        io_lsbs_928,
  output        io_lsbs_929,
  output        io_lsbs_930,
  output        io_lsbs_931,
  output        io_lsbs_932,
  output        io_lsbs_933,
  output        io_lsbs_934,
  output        io_lsbs_935,
  output        io_lsbs_936,
  output        io_lsbs_937,
  output        io_lsbs_938,
  output        io_lsbs_939,
  output        io_lsbs_940,
  output        io_lsbs_941,
  output        io_lsbs_942,
  output        io_lsbs_943,
  output        io_lsbs_944,
  output        io_lsbs_945,
  output        io_lsbs_946,
  output        io_lsbs_947,
  output        io_lsbs_948,
  output        io_lsbs_949,
  output        io_lsbs_950,
  output        io_lsbs_951,
  output        io_lsbs_952,
  output        io_lsbs_953,
  output        io_lsbs_954,
  output        io_lsbs_955,
  output        io_lsbs_956,
  output        io_lsbs_957,
  output        io_lsbs_958,
  output        io_lsbs_959,
  output        io_lsbs_960,
  output        io_lsbs_961,
  output        io_lsbs_962,
  output        io_lsbs_963,
  output        io_lsbs_964,
  output        io_lsbs_965,
  output        io_lsbs_966,
  output        io_lsbs_967,
  output        io_lsbs_968,
  output        io_lsbs_969,
  output        io_lsbs_970,
  output        io_lsbs_971,
  output        io_lsbs_972,
  output        io_lsbs_973,
  output        io_lsbs_974,
  output        io_lsbs_975,
  output        io_lsbs_976,
  output        io_lsbs_977,
  output        io_lsbs_978,
  output        io_lsbs_979,
  output        io_lsbs_980,
  output        io_lsbs_981,
  output        io_lsbs_982,
  output        io_lsbs_983,
  output        io_lsbs_984,
  output        io_lsbs_985,
  output        io_lsbs_986,
  output        io_lsbs_987,
  output        io_lsbs_988,
  output        io_lsbs_989,
  output        io_lsbs_990,
  output        io_lsbs_991,
  output        io_lsbs_992,
  output        io_lsbs_993,
  output        io_lsbs_994,
  output        io_lsbs_995,
  output        io_lsbs_996,
  output        io_lsbs_997,
  output        io_lsbs_998,
  output        io_lsbs_999,
  output        io_lsbs_1000,
  output        io_lsbs_1001,
  output        io_lsbs_1002,
  output        io_lsbs_1003,
  output        io_lsbs_1004,
  output        io_lsbs_1005,
  output        io_lsbs_1006,
  output        io_lsbs_1007,
  output        io_lsbs_1008,
  output        io_lsbs_1009,
  output        io_lsbs_1010,
  output        io_lsbs_1011,
  output        io_lsbs_1012,
  output        io_lsbs_1013,
  output        io_lsbs_1014,
  output        io_lsbs_1015,
  output        io_lsbs_1016,
  output        io_lsbs_1017,
  output        io_lsbs_1018,
  output        io_lsbs_1019,
  output        io_lsbs_1020,
  output        io_lsbs_1021,
  output        io_lsbs_1022,
  output        io_lsbs_1023
);
  wire  ces_0_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_0_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_0_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_1_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_2_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_3_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_4_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_5_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_6_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_7_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_8_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_9_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_10_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_11_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_12_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_13_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_14_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_15_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_16_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_17_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_18_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_19_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_20_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_21_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_22_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_23_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_24_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_25_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_26_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_27_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_28_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_29_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_30_31_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_0_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_1_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_1_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_1_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_1_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_1_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_1_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_1_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_1_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_1_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_2_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_2_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_2_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_2_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_2_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_2_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_2_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_2_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_2_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_3_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_3_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_3_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_3_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_3_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_3_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_3_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_3_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_3_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_4_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_4_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_4_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_4_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_4_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_4_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_4_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_4_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_4_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_5_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_5_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_5_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_5_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_5_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_5_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_5_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_5_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_5_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_6_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_6_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_6_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_6_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_6_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_6_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_6_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_6_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_6_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_7_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_7_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_7_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_7_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_7_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_7_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_7_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_7_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_7_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_8_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_8_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_8_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_8_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_8_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_8_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_8_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_8_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_8_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_9_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_9_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_9_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_9_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_9_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_9_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_9_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_9_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_9_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_10_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_10_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_10_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_10_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_10_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_10_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_10_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_10_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_10_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_11_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_11_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_11_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_11_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_11_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_11_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_11_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_11_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_11_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_12_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_12_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_12_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_12_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_12_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_12_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_12_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_12_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_12_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_13_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_13_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_13_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_13_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_13_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_13_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_13_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_13_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_13_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_14_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_14_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_14_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_14_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_14_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_14_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_14_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_14_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_14_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_15_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_15_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_15_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_15_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_15_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_15_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_15_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_15_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_15_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_16_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_16_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_16_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_16_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_16_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_16_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_16_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_16_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_16_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_17_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_17_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_17_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_17_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_17_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_17_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_17_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_17_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_17_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_18_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_18_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_18_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_18_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_18_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_18_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_18_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_18_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_18_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_19_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_19_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_19_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_19_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_19_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_19_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_19_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_19_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_19_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_20_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_20_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_20_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_20_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_20_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_20_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_20_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_20_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_20_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_21_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_21_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_21_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_21_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_21_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_21_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_21_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_21_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_21_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_22_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_22_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_22_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_22_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_22_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_22_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_22_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_22_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_22_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_23_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_23_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_23_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_23_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_23_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_23_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_23_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_23_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_23_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_24_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_24_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_24_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_24_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_24_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_24_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_24_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_24_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_24_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_25_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_25_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_25_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_25_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_25_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_25_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_25_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_25_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_25_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_26_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_26_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_26_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_26_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_26_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_26_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_26_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_26_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_26_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_27_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_27_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_27_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_27_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_27_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_27_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_27_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_27_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_27_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_28_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_28_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_28_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_28_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_28_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_28_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_28_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_28_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_28_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_29_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_29_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_29_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_29_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_29_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_29_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_29_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_29_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_29_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_30_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_30_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_30_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_30_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_30_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_30_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_30_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_30_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_30_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_31_clock; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_31_io_ins_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_31_io_ins_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_31_io_ins_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_31_io_ins_3; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_31_io_outs_0; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_31_io_outs_1; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_31_io_outs_2; // @[MockArray.scala 36:52]
  wire [63:0] ces_31_31_io_outs_3; // @[MockArray.scala 36:52]
  Element ces_0_0 ( // @[MockArray.scala 36:52]
    .clock(ces_0_0_clock),
    .io_ins_0(ces_0_0_io_ins_0),
    .io_ins_1(ces_0_0_io_ins_1),
    .io_ins_2(ces_0_0_io_ins_2),
    .io_ins_3(ces_0_0_io_ins_3),
    .io_outs_0(ces_0_0_io_outs_0),
    .io_outs_1(ces_0_0_io_outs_1),
    .io_outs_2(ces_0_0_io_outs_2),
    .io_outs_3(ces_0_0_io_outs_3)
  );
  Element ces_0_1 ( // @[MockArray.scala 36:52]
    .clock(ces_0_1_clock),
    .io_ins_0(ces_0_1_io_ins_0),
    .io_ins_1(ces_0_1_io_ins_1),
    .io_ins_2(ces_0_1_io_ins_2),
    .io_ins_3(ces_0_1_io_ins_3),
    .io_outs_0(ces_0_1_io_outs_0),
    .io_outs_1(ces_0_1_io_outs_1),
    .io_outs_2(ces_0_1_io_outs_2),
    .io_outs_3(ces_0_1_io_outs_3)
  );
  Element ces_0_2 ( // @[MockArray.scala 36:52]
    .clock(ces_0_2_clock),
    .io_ins_0(ces_0_2_io_ins_0),
    .io_ins_1(ces_0_2_io_ins_1),
    .io_ins_2(ces_0_2_io_ins_2),
    .io_ins_3(ces_0_2_io_ins_3),
    .io_outs_0(ces_0_2_io_outs_0),
    .io_outs_1(ces_0_2_io_outs_1),
    .io_outs_2(ces_0_2_io_outs_2),
    .io_outs_3(ces_0_2_io_outs_3)
  );
  Element ces_0_3 ( // @[MockArray.scala 36:52]
    .clock(ces_0_3_clock),
    .io_ins_0(ces_0_3_io_ins_0),
    .io_ins_1(ces_0_3_io_ins_1),
    .io_ins_2(ces_0_3_io_ins_2),
    .io_ins_3(ces_0_3_io_ins_3),
    .io_outs_0(ces_0_3_io_outs_0),
    .io_outs_1(ces_0_3_io_outs_1),
    .io_outs_2(ces_0_3_io_outs_2),
    .io_outs_3(ces_0_3_io_outs_3)
  );
  Element ces_0_4 ( // @[MockArray.scala 36:52]
    .clock(ces_0_4_clock),
    .io_ins_0(ces_0_4_io_ins_0),
    .io_ins_1(ces_0_4_io_ins_1),
    .io_ins_2(ces_0_4_io_ins_2),
    .io_ins_3(ces_0_4_io_ins_3),
    .io_outs_0(ces_0_4_io_outs_0),
    .io_outs_1(ces_0_4_io_outs_1),
    .io_outs_2(ces_0_4_io_outs_2),
    .io_outs_3(ces_0_4_io_outs_3)
  );
  Element ces_0_5 ( // @[MockArray.scala 36:52]
    .clock(ces_0_5_clock),
    .io_ins_0(ces_0_5_io_ins_0),
    .io_ins_1(ces_0_5_io_ins_1),
    .io_ins_2(ces_0_5_io_ins_2),
    .io_ins_3(ces_0_5_io_ins_3),
    .io_outs_0(ces_0_5_io_outs_0),
    .io_outs_1(ces_0_5_io_outs_1),
    .io_outs_2(ces_0_5_io_outs_2),
    .io_outs_3(ces_0_5_io_outs_3)
  );
  Element ces_0_6 ( // @[MockArray.scala 36:52]
    .clock(ces_0_6_clock),
    .io_ins_0(ces_0_6_io_ins_0),
    .io_ins_1(ces_0_6_io_ins_1),
    .io_ins_2(ces_0_6_io_ins_2),
    .io_ins_3(ces_0_6_io_ins_3),
    .io_outs_0(ces_0_6_io_outs_0),
    .io_outs_1(ces_0_6_io_outs_1),
    .io_outs_2(ces_0_6_io_outs_2),
    .io_outs_3(ces_0_6_io_outs_3)
  );
  Element ces_0_7 ( // @[MockArray.scala 36:52]
    .clock(ces_0_7_clock),
    .io_ins_0(ces_0_7_io_ins_0),
    .io_ins_1(ces_0_7_io_ins_1),
    .io_ins_2(ces_0_7_io_ins_2),
    .io_ins_3(ces_0_7_io_ins_3),
    .io_outs_0(ces_0_7_io_outs_0),
    .io_outs_1(ces_0_7_io_outs_1),
    .io_outs_2(ces_0_7_io_outs_2),
    .io_outs_3(ces_0_7_io_outs_3)
  );
  Element ces_0_8 ( // @[MockArray.scala 36:52]
    .clock(ces_0_8_clock),
    .io_ins_0(ces_0_8_io_ins_0),
    .io_ins_1(ces_0_8_io_ins_1),
    .io_ins_2(ces_0_8_io_ins_2),
    .io_ins_3(ces_0_8_io_ins_3),
    .io_outs_0(ces_0_8_io_outs_0),
    .io_outs_1(ces_0_8_io_outs_1),
    .io_outs_2(ces_0_8_io_outs_2),
    .io_outs_3(ces_0_8_io_outs_3)
  );
  Element ces_0_9 ( // @[MockArray.scala 36:52]
    .clock(ces_0_9_clock),
    .io_ins_0(ces_0_9_io_ins_0),
    .io_ins_1(ces_0_9_io_ins_1),
    .io_ins_2(ces_0_9_io_ins_2),
    .io_ins_3(ces_0_9_io_ins_3),
    .io_outs_0(ces_0_9_io_outs_0),
    .io_outs_1(ces_0_9_io_outs_1),
    .io_outs_2(ces_0_9_io_outs_2),
    .io_outs_3(ces_0_9_io_outs_3)
  );
  Element ces_0_10 ( // @[MockArray.scala 36:52]
    .clock(ces_0_10_clock),
    .io_ins_0(ces_0_10_io_ins_0),
    .io_ins_1(ces_0_10_io_ins_1),
    .io_ins_2(ces_0_10_io_ins_2),
    .io_ins_3(ces_0_10_io_ins_3),
    .io_outs_0(ces_0_10_io_outs_0),
    .io_outs_1(ces_0_10_io_outs_1),
    .io_outs_2(ces_0_10_io_outs_2),
    .io_outs_3(ces_0_10_io_outs_3)
  );
  Element ces_0_11 ( // @[MockArray.scala 36:52]
    .clock(ces_0_11_clock),
    .io_ins_0(ces_0_11_io_ins_0),
    .io_ins_1(ces_0_11_io_ins_1),
    .io_ins_2(ces_0_11_io_ins_2),
    .io_ins_3(ces_0_11_io_ins_3),
    .io_outs_0(ces_0_11_io_outs_0),
    .io_outs_1(ces_0_11_io_outs_1),
    .io_outs_2(ces_0_11_io_outs_2),
    .io_outs_3(ces_0_11_io_outs_3)
  );
  Element ces_0_12 ( // @[MockArray.scala 36:52]
    .clock(ces_0_12_clock),
    .io_ins_0(ces_0_12_io_ins_0),
    .io_ins_1(ces_0_12_io_ins_1),
    .io_ins_2(ces_0_12_io_ins_2),
    .io_ins_3(ces_0_12_io_ins_3),
    .io_outs_0(ces_0_12_io_outs_0),
    .io_outs_1(ces_0_12_io_outs_1),
    .io_outs_2(ces_0_12_io_outs_2),
    .io_outs_3(ces_0_12_io_outs_3)
  );
  Element ces_0_13 ( // @[MockArray.scala 36:52]
    .clock(ces_0_13_clock),
    .io_ins_0(ces_0_13_io_ins_0),
    .io_ins_1(ces_0_13_io_ins_1),
    .io_ins_2(ces_0_13_io_ins_2),
    .io_ins_3(ces_0_13_io_ins_3),
    .io_outs_0(ces_0_13_io_outs_0),
    .io_outs_1(ces_0_13_io_outs_1),
    .io_outs_2(ces_0_13_io_outs_2),
    .io_outs_3(ces_0_13_io_outs_3)
  );
  Element ces_0_14 ( // @[MockArray.scala 36:52]
    .clock(ces_0_14_clock),
    .io_ins_0(ces_0_14_io_ins_0),
    .io_ins_1(ces_0_14_io_ins_1),
    .io_ins_2(ces_0_14_io_ins_2),
    .io_ins_3(ces_0_14_io_ins_3),
    .io_outs_0(ces_0_14_io_outs_0),
    .io_outs_1(ces_0_14_io_outs_1),
    .io_outs_2(ces_0_14_io_outs_2),
    .io_outs_3(ces_0_14_io_outs_3)
  );
  Element ces_0_15 ( // @[MockArray.scala 36:52]
    .clock(ces_0_15_clock),
    .io_ins_0(ces_0_15_io_ins_0),
    .io_ins_1(ces_0_15_io_ins_1),
    .io_ins_2(ces_0_15_io_ins_2),
    .io_ins_3(ces_0_15_io_ins_3),
    .io_outs_0(ces_0_15_io_outs_0),
    .io_outs_1(ces_0_15_io_outs_1),
    .io_outs_2(ces_0_15_io_outs_2),
    .io_outs_3(ces_0_15_io_outs_3)
  );
  Element ces_0_16 ( // @[MockArray.scala 36:52]
    .clock(ces_0_16_clock),
    .io_ins_0(ces_0_16_io_ins_0),
    .io_ins_1(ces_0_16_io_ins_1),
    .io_ins_2(ces_0_16_io_ins_2),
    .io_ins_3(ces_0_16_io_ins_3),
    .io_outs_0(ces_0_16_io_outs_0),
    .io_outs_1(ces_0_16_io_outs_1),
    .io_outs_2(ces_0_16_io_outs_2),
    .io_outs_3(ces_0_16_io_outs_3)
  );
  Element ces_0_17 ( // @[MockArray.scala 36:52]
    .clock(ces_0_17_clock),
    .io_ins_0(ces_0_17_io_ins_0),
    .io_ins_1(ces_0_17_io_ins_1),
    .io_ins_2(ces_0_17_io_ins_2),
    .io_ins_3(ces_0_17_io_ins_3),
    .io_outs_0(ces_0_17_io_outs_0),
    .io_outs_1(ces_0_17_io_outs_1),
    .io_outs_2(ces_0_17_io_outs_2),
    .io_outs_3(ces_0_17_io_outs_3)
  );
  Element ces_0_18 ( // @[MockArray.scala 36:52]
    .clock(ces_0_18_clock),
    .io_ins_0(ces_0_18_io_ins_0),
    .io_ins_1(ces_0_18_io_ins_1),
    .io_ins_2(ces_0_18_io_ins_2),
    .io_ins_3(ces_0_18_io_ins_3),
    .io_outs_0(ces_0_18_io_outs_0),
    .io_outs_1(ces_0_18_io_outs_1),
    .io_outs_2(ces_0_18_io_outs_2),
    .io_outs_3(ces_0_18_io_outs_3)
  );
  Element ces_0_19 ( // @[MockArray.scala 36:52]
    .clock(ces_0_19_clock),
    .io_ins_0(ces_0_19_io_ins_0),
    .io_ins_1(ces_0_19_io_ins_1),
    .io_ins_2(ces_0_19_io_ins_2),
    .io_ins_3(ces_0_19_io_ins_3),
    .io_outs_0(ces_0_19_io_outs_0),
    .io_outs_1(ces_0_19_io_outs_1),
    .io_outs_2(ces_0_19_io_outs_2),
    .io_outs_3(ces_0_19_io_outs_3)
  );
  Element ces_0_20 ( // @[MockArray.scala 36:52]
    .clock(ces_0_20_clock),
    .io_ins_0(ces_0_20_io_ins_0),
    .io_ins_1(ces_0_20_io_ins_1),
    .io_ins_2(ces_0_20_io_ins_2),
    .io_ins_3(ces_0_20_io_ins_3),
    .io_outs_0(ces_0_20_io_outs_0),
    .io_outs_1(ces_0_20_io_outs_1),
    .io_outs_2(ces_0_20_io_outs_2),
    .io_outs_3(ces_0_20_io_outs_3)
  );
  Element ces_0_21 ( // @[MockArray.scala 36:52]
    .clock(ces_0_21_clock),
    .io_ins_0(ces_0_21_io_ins_0),
    .io_ins_1(ces_0_21_io_ins_1),
    .io_ins_2(ces_0_21_io_ins_2),
    .io_ins_3(ces_0_21_io_ins_3),
    .io_outs_0(ces_0_21_io_outs_0),
    .io_outs_1(ces_0_21_io_outs_1),
    .io_outs_2(ces_0_21_io_outs_2),
    .io_outs_3(ces_0_21_io_outs_3)
  );
  Element ces_0_22 ( // @[MockArray.scala 36:52]
    .clock(ces_0_22_clock),
    .io_ins_0(ces_0_22_io_ins_0),
    .io_ins_1(ces_0_22_io_ins_1),
    .io_ins_2(ces_0_22_io_ins_2),
    .io_ins_3(ces_0_22_io_ins_3),
    .io_outs_0(ces_0_22_io_outs_0),
    .io_outs_1(ces_0_22_io_outs_1),
    .io_outs_2(ces_0_22_io_outs_2),
    .io_outs_3(ces_0_22_io_outs_3)
  );
  Element ces_0_23 ( // @[MockArray.scala 36:52]
    .clock(ces_0_23_clock),
    .io_ins_0(ces_0_23_io_ins_0),
    .io_ins_1(ces_0_23_io_ins_1),
    .io_ins_2(ces_0_23_io_ins_2),
    .io_ins_3(ces_0_23_io_ins_3),
    .io_outs_0(ces_0_23_io_outs_0),
    .io_outs_1(ces_0_23_io_outs_1),
    .io_outs_2(ces_0_23_io_outs_2),
    .io_outs_3(ces_0_23_io_outs_3)
  );
  Element ces_0_24 ( // @[MockArray.scala 36:52]
    .clock(ces_0_24_clock),
    .io_ins_0(ces_0_24_io_ins_0),
    .io_ins_1(ces_0_24_io_ins_1),
    .io_ins_2(ces_0_24_io_ins_2),
    .io_ins_3(ces_0_24_io_ins_3),
    .io_outs_0(ces_0_24_io_outs_0),
    .io_outs_1(ces_0_24_io_outs_1),
    .io_outs_2(ces_0_24_io_outs_2),
    .io_outs_3(ces_0_24_io_outs_3)
  );
  Element ces_0_25 ( // @[MockArray.scala 36:52]
    .clock(ces_0_25_clock),
    .io_ins_0(ces_0_25_io_ins_0),
    .io_ins_1(ces_0_25_io_ins_1),
    .io_ins_2(ces_0_25_io_ins_2),
    .io_ins_3(ces_0_25_io_ins_3),
    .io_outs_0(ces_0_25_io_outs_0),
    .io_outs_1(ces_0_25_io_outs_1),
    .io_outs_2(ces_0_25_io_outs_2),
    .io_outs_3(ces_0_25_io_outs_3)
  );
  Element ces_0_26 ( // @[MockArray.scala 36:52]
    .clock(ces_0_26_clock),
    .io_ins_0(ces_0_26_io_ins_0),
    .io_ins_1(ces_0_26_io_ins_1),
    .io_ins_2(ces_0_26_io_ins_2),
    .io_ins_3(ces_0_26_io_ins_3),
    .io_outs_0(ces_0_26_io_outs_0),
    .io_outs_1(ces_0_26_io_outs_1),
    .io_outs_2(ces_0_26_io_outs_2),
    .io_outs_3(ces_0_26_io_outs_3)
  );
  Element ces_0_27 ( // @[MockArray.scala 36:52]
    .clock(ces_0_27_clock),
    .io_ins_0(ces_0_27_io_ins_0),
    .io_ins_1(ces_0_27_io_ins_1),
    .io_ins_2(ces_0_27_io_ins_2),
    .io_ins_3(ces_0_27_io_ins_3),
    .io_outs_0(ces_0_27_io_outs_0),
    .io_outs_1(ces_0_27_io_outs_1),
    .io_outs_2(ces_0_27_io_outs_2),
    .io_outs_3(ces_0_27_io_outs_3)
  );
  Element ces_0_28 ( // @[MockArray.scala 36:52]
    .clock(ces_0_28_clock),
    .io_ins_0(ces_0_28_io_ins_0),
    .io_ins_1(ces_0_28_io_ins_1),
    .io_ins_2(ces_0_28_io_ins_2),
    .io_ins_3(ces_0_28_io_ins_3),
    .io_outs_0(ces_0_28_io_outs_0),
    .io_outs_1(ces_0_28_io_outs_1),
    .io_outs_2(ces_0_28_io_outs_2),
    .io_outs_3(ces_0_28_io_outs_3)
  );
  Element ces_0_29 ( // @[MockArray.scala 36:52]
    .clock(ces_0_29_clock),
    .io_ins_0(ces_0_29_io_ins_0),
    .io_ins_1(ces_0_29_io_ins_1),
    .io_ins_2(ces_0_29_io_ins_2),
    .io_ins_3(ces_0_29_io_ins_3),
    .io_outs_0(ces_0_29_io_outs_0),
    .io_outs_1(ces_0_29_io_outs_1),
    .io_outs_2(ces_0_29_io_outs_2),
    .io_outs_3(ces_0_29_io_outs_3)
  );
  Element ces_0_30 ( // @[MockArray.scala 36:52]
    .clock(ces_0_30_clock),
    .io_ins_0(ces_0_30_io_ins_0),
    .io_ins_1(ces_0_30_io_ins_1),
    .io_ins_2(ces_0_30_io_ins_2),
    .io_ins_3(ces_0_30_io_ins_3),
    .io_outs_0(ces_0_30_io_outs_0),
    .io_outs_1(ces_0_30_io_outs_1),
    .io_outs_2(ces_0_30_io_outs_2),
    .io_outs_3(ces_0_30_io_outs_3)
  );
  Element ces_0_31 ( // @[MockArray.scala 36:52]
    .clock(ces_0_31_clock),
    .io_ins_0(ces_0_31_io_ins_0),
    .io_ins_1(ces_0_31_io_ins_1),
    .io_ins_2(ces_0_31_io_ins_2),
    .io_ins_3(ces_0_31_io_ins_3),
    .io_outs_0(ces_0_31_io_outs_0),
    .io_outs_1(ces_0_31_io_outs_1),
    .io_outs_2(ces_0_31_io_outs_2),
    .io_outs_3(ces_0_31_io_outs_3)
  );
  Element ces_1_0 ( // @[MockArray.scala 36:52]
    .clock(ces_1_0_clock),
    .io_ins_0(ces_1_0_io_ins_0),
    .io_ins_1(ces_1_0_io_ins_1),
    .io_ins_2(ces_1_0_io_ins_2),
    .io_ins_3(ces_1_0_io_ins_3),
    .io_outs_0(ces_1_0_io_outs_0),
    .io_outs_1(ces_1_0_io_outs_1),
    .io_outs_2(ces_1_0_io_outs_2),
    .io_outs_3(ces_1_0_io_outs_3)
  );
  Element ces_1_1 ( // @[MockArray.scala 36:52]
    .clock(ces_1_1_clock),
    .io_ins_0(ces_1_1_io_ins_0),
    .io_ins_1(ces_1_1_io_ins_1),
    .io_ins_2(ces_1_1_io_ins_2),
    .io_ins_3(ces_1_1_io_ins_3),
    .io_outs_0(ces_1_1_io_outs_0),
    .io_outs_1(ces_1_1_io_outs_1),
    .io_outs_2(ces_1_1_io_outs_2),
    .io_outs_3(ces_1_1_io_outs_3)
  );
  Element ces_1_2 ( // @[MockArray.scala 36:52]
    .clock(ces_1_2_clock),
    .io_ins_0(ces_1_2_io_ins_0),
    .io_ins_1(ces_1_2_io_ins_1),
    .io_ins_2(ces_1_2_io_ins_2),
    .io_ins_3(ces_1_2_io_ins_3),
    .io_outs_0(ces_1_2_io_outs_0),
    .io_outs_1(ces_1_2_io_outs_1),
    .io_outs_2(ces_1_2_io_outs_2),
    .io_outs_3(ces_1_2_io_outs_3)
  );
  Element ces_1_3 ( // @[MockArray.scala 36:52]
    .clock(ces_1_3_clock),
    .io_ins_0(ces_1_3_io_ins_0),
    .io_ins_1(ces_1_3_io_ins_1),
    .io_ins_2(ces_1_3_io_ins_2),
    .io_ins_3(ces_1_3_io_ins_3),
    .io_outs_0(ces_1_3_io_outs_0),
    .io_outs_1(ces_1_3_io_outs_1),
    .io_outs_2(ces_1_3_io_outs_2),
    .io_outs_3(ces_1_3_io_outs_3)
  );
  Element ces_1_4 ( // @[MockArray.scala 36:52]
    .clock(ces_1_4_clock),
    .io_ins_0(ces_1_4_io_ins_0),
    .io_ins_1(ces_1_4_io_ins_1),
    .io_ins_2(ces_1_4_io_ins_2),
    .io_ins_3(ces_1_4_io_ins_3),
    .io_outs_0(ces_1_4_io_outs_0),
    .io_outs_1(ces_1_4_io_outs_1),
    .io_outs_2(ces_1_4_io_outs_2),
    .io_outs_3(ces_1_4_io_outs_3)
  );
  Element ces_1_5 ( // @[MockArray.scala 36:52]
    .clock(ces_1_5_clock),
    .io_ins_0(ces_1_5_io_ins_0),
    .io_ins_1(ces_1_5_io_ins_1),
    .io_ins_2(ces_1_5_io_ins_2),
    .io_ins_3(ces_1_5_io_ins_3),
    .io_outs_0(ces_1_5_io_outs_0),
    .io_outs_1(ces_1_5_io_outs_1),
    .io_outs_2(ces_1_5_io_outs_2),
    .io_outs_3(ces_1_5_io_outs_3)
  );
  Element ces_1_6 ( // @[MockArray.scala 36:52]
    .clock(ces_1_6_clock),
    .io_ins_0(ces_1_6_io_ins_0),
    .io_ins_1(ces_1_6_io_ins_1),
    .io_ins_2(ces_1_6_io_ins_2),
    .io_ins_3(ces_1_6_io_ins_3),
    .io_outs_0(ces_1_6_io_outs_0),
    .io_outs_1(ces_1_6_io_outs_1),
    .io_outs_2(ces_1_6_io_outs_2),
    .io_outs_3(ces_1_6_io_outs_3)
  );
  Element ces_1_7 ( // @[MockArray.scala 36:52]
    .clock(ces_1_7_clock),
    .io_ins_0(ces_1_7_io_ins_0),
    .io_ins_1(ces_1_7_io_ins_1),
    .io_ins_2(ces_1_7_io_ins_2),
    .io_ins_3(ces_1_7_io_ins_3),
    .io_outs_0(ces_1_7_io_outs_0),
    .io_outs_1(ces_1_7_io_outs_1),
    .io_outs_2(ces_1_7_io_outs_2),
    .io_outs_3(ces_1_7_io_outs_3)
  );
  Element ces_1_8 ( // @[MockArray.scala 36:52]
    .clock(ces_1_8_clock),
    .io_ins_0(ces_1_8_io_ins_0),
    .io_ins_1(ces_1_8_io_ins_1),
    .io_ins_2(ces_1_8_io_ins_2),
    .io_ins_3(ces_1_8_io_ins_3),
    .io_outs_0(ces_1_8_io_outs_0),
    .io_outs_1(ces_1_8_io_outs_1),
    .io_outs_2(ces_1_8_io_outs_2),
    .io_outs_3(ces_1_8_io_outs_3)
  );
  Element ces_1_9 ( // @[MockArray.scala 36:52]
    .clock(ces_1_9_clock),
    .io_ins_0(ces_1_9_io_ins_0),
    .io_ins_1(ces_1_9_io_ins_1),
    .io_ins_2(ces_1_9_io_ins_2),
    .io_ins_3(ces_1_9_io_ins_3),
    .io_outs_0(ces_1_9_io_outs_0),
    .io_outs_1(ces_1_9_io_outs_1),
    .io_outs_2(ces_1_9_io_outs_2),
    .io_outs_3(ces_1_9_io_outs_3)
  );
  Element ces_1_10 ( // @[MockArray.scala 36:52]
    .clock(ces_1_10_clock),
    .io_ins_0(ces_1_10_io_ins_0),
    .io_ins_1(ces_1_10_io_ins_1),
    .io_ins_2(ces_1_10_io_ins_2),
    .io_ins_3(ces_1_10_io_ins_3),
    .io_outs_0(ces_1_10_io_outs_0),
    .io_outs_1(ces_1_10_io_outs_1),
    .io_outs_2(ces_1_10_io_outs_2),
    .io_outs_3(ces_1_10_io_outs_3)
  );
  Element ces_1_11 ( // @[MockArray.scala 36:52]
    .clock(ces_1_11_clock),
    .io_ins_0(ces_1_11_io_ins_0),
    .io_ins_1(ces_1_11_io_ins_1),
    .io_ins_2(ces_1_11_io_ins_2),
    .io_ins_3(ces_1_11_io_ins_3),
    .io_outs_0(ces_1_11_io_outs_0),
    .io_outs_1(ces_1_11_io_outs_1),
    .io_outs_2(ces_1_11_io_outs_2),
    .io_outs_3(ces_1_11_io_outs_3)
  );
  Element ces_1_12 ( // @[MockArray.scala 36:52]
    .clock(ces_1_12_clock),
    .io_ins_0(ces_1_12_io_ins_0),
    .io_ins_1(ces_1_12_io_ins_1),
    .io_ins_2(ces_1_12_io_ins_2),
    .io_ins_3(ces_1_12_io_ins_3),
    .io_outs_0(ces_1_12_io_outs_0),
    .io_outs_1(ces_1_12_io_outs_1),
    .io_outs_2(ces_1_12_io_outs_2),
    .io_outs_3(ces_1_12_io_outs_3)
  );
  Element ces_1_13 ( // @[MockArray.scala 36:52]
    .clock(ces_1_13_clock),
    .io_ins_0(ces_1_13_io_ins_0),
    .io_ins_1(ces_1_13_io_ins_1),
    .io_ins_2(ces_1_13_io_ins_2),
    .io_ins_3(ces_1_13_io_ins_3),
    .io_outs_0(ces_1_13_io_outs_0),
    .io_outs_1(ces_1_13_io_outs_1),
    .io_outs_2(ces_1_13_io_outs_2),
    .io_outs_3(ces_1_13_io_outs_3)
  );
  Element ces_1_14 ( // @[MockArray.scala 36:52]
    .clock(ces_1_14_clock),
    .io_ins_0(ces_1_14_io_ins_0),
    .io_ins_1(ces_1_14_io_ins_1),
    .io_ins_2(ces_1_14_io_ins_2),
    .io_ins_3(ces_1_14_io_ins_3),
    .io_outs_0(ces_1_14_io_outs_0),
    .io_outs_1(ces_1_14_io_outs_1),
    .io_outs_2(ces_1_14_io_outs_2),
    .io_outs_3(ces_1_14_io_outs_3)
  );
  Element ces_1_15 ( // @[MockArray.scala 36:52]
    .clock(ces_1_15_clock),
    .io_ins_0(ces_1_15_io_ins_0),
    .io_ins_1(ces_1_15_io_ins_1),
    .io_ins_2(ces_1_15_io_ins_2),
    .io_ins_3(ces_1_15_io_ins_3),
    .io_outs_0(ces_1_15_io_outs_0),
    .io_outs_1(ces_1_15_io_outs_1),
    .io_outs_2(ces_1_15_io_outs_2),
    .io_outs_3(ces_1_15_io_outs_3)
  );
  Element ces_1_16 ( // @[MockArray.scala 36:52]
    .clock(ces_1_16_clock),
    .io_ins_0(ces_1_16_io_ins_0),
    .io_ins_1(ces_1_16_io_ins_1),
    .io_ins_2(ces_1_16_io_ins_2),
    .io_ins_3(ces_1_16_io_ins_3),
    .io_outs_0(ces_1_16_io_outs_0),
    .io_outs_1(ces_1_16_io_outs_1),
    .io_outs_2(ces_1_16_io_outs_2),
    .io_outs_3(ces_1_16_io_outs_3)
  );
  Element ces_1_17 ( // @[MockArray.scala 36:52]
    .clock(ces_1_17_clock),
    .io_ins_0(ces_1_17_io_ins_0),
    .io_ins_1(ces_1_17_io_ins_1),
    .io_ins_2(ces_1_17_io_ins_2),
    .io_ins_3(ces_1_17_io_ins_3),
    .io_outs_0(ces_1_17_io_outs_0),
    .io_outs_1(ces_1_17_io_outs_1),
    .io_outs_2(ces_1_17_io_outs_2),
    .io_outs_3(ces_1_17_io_outs_3)
  );
  Element ces_1_18 ( // @[MockArray.scala 36:52]
    .clock(ces_1_18_clock),
    .io_ins_0(ces_1_18_io_ins_0),
    .io_ins_1(ces_1_18_io_ins_1),
    .io_ins_2(ces_1_18_io_ins_2),
    .io_ins_3(ces_1_18_io_ins_3),
    .io_outs_0(ces_1_18_io_outs_0),
    .io_outs_1(ces_1_18_io_outs_1),
    .io_outs_2(ces_1_18_io_outs_2),
    .io_outs_3(ces_1_18_io_outs_3)
  );
  Element ces_1_19 ( // @[MockArray.scala 36:52]
    .clock(ces_1_19_clock),
    .io_ins_0(ces_1_19_io_ins_0),
    .io_ins_1(ces_1_19_io_ins_1),
    .io_ins_2(ces_1_19_io_ins_2),
    .io_ins_3(ces_1_19_io_ins_3),
    .io_outs_0(ces_1_19_io_outs_0),
    .io_outs_1(ces_1_19_io_outs_1),
    .io_outs_2(ces_1_19_io_outs_2),
    .io_outs_3(ces_1_19_io_outs_3)
  );
  Element ces_1_20 ( // @[MockArray.scala 36:52]
    .clock(ces_1_20_clock),
    .io_ins_0(ces_1_20_io_ins_0),
    .io_ins_1(ces_1_20_io_ins_1),
    .io_ins_2(ces_1_20_io_ins_2),
    .io_ins_3(ces_1_20_io_ins_3),
    .io_outs_0(ces_1_20_io_outs_0),
    .io_outs_1(ces_1_20_io_outs_1),
    .io_outs_2(ces_1_20_io_outs_2),
    .io_outs_3(ces_1_20_io_outs_3)
  );
  Element ces_1_21 ( // @[MockArray.scala 36:52]
    .clock(ces_1_21_clock),
    .io_ins_0(ces_1_21_io_ins_0),
    .io_ins_1(ces_1_21_io_ins_1),
    .io_ins_2(ces_1_21_io_ins_2),
    .io_ins_3(ces_1_21_io_ins_3),
    .io_outs_0(ces_1_21_io_outs_0),
    .io_outs_1(ces_1_21_io_outs_1),
    .io_outs_2(ces_1_21_io_outs_2),
    .io_outs_3(ces_1_21_io_outs_3)
  );
  Element ces_1_22 ( // @[MockArray.scala 36:52]
    .clock(ces_1_22_clock),
    .io_ins_0(ces_1_22_io_ins_0),
    .io_ins_1(ces_1_22_io_ins_1),
    .io_ins_2(ces_1_22_io_ins_2),
    .io_ins_3(ces_1_22_io_ins_3),
    .io_outs_0(ces_1_22_io_outs_0),
    .io_outs_1(ces_1_22_io_outs_1),
    .io_outs_2(ces_1_22_io_outs_2),
    .io_outs_3(ces_1_22_io_outs_3)
  );
  Element ces_1_23 ( // @[MockArray.scala 36:52]
    .clock(ces_1_23_clock),
    .io_ins_0(ces_1_23_io_ins_0),
    .io_ins_1(ces_1_23_io_ins_1),
    .io_ins_2(ces_1_23_io_ins_2),
    .io_ins_3(ces_1_23_io_ins_3),
    .io_outs_0(ces_1_23_io_outs_0),
    .io_outs_1(ces_1_23_io_outs_1),
    .io_outs_2(ces_1_23_io_outs_2),
    .io_outs_3(ces_1_23_io_outs_3)
  );
  Element ces_1_24 ( // @[MockArray.scala 36:52]
    .clock(ces_1_24_clock),
    .io_ins_0(ces_1_24_io_ins_0),
    .io_ins_1(ces_1_24_io_ins_1),
    .io_ins_2(ces_1_24_io_ins_2),
    .io_ins_3(ces_1_24_io_ins_3),
    .io_outs_0(ces_1_24_io_outs_0),
    .io_outs_1(ces_1_24_io_outs_1),
    .io_outs_2(ces_1_24_io_outs_2),
    .io_outs_3(ces_1_24_io_outs_3)
  );
  Element ces_1_25 ( // @[MockArray.scala 36:52]
    .clock(ces_1_25_clock),
    .io_ins_0(ces_1_25_io_ins_0),
    .io_ins_1(ces_1_25_io_ins_1),
    .io_ins_2(ces_1_25_io_ins_2),
    .io_ins_3(ces_1_25_io_ins_3),
    .io_outs_0(ces_1_25_io_outs_0),
    .io_outs_1(ces_1_25_io_outs_1),
    .io_outs_2(ces_1_25_io_outs_2),
    .io_outs_3(ces_1_25_io_outs_3)
  );
  Element ces_1_26 ( // @[MockArray.scala 36:52]
    .clock(ces_1_26_clock),
    .io_ins_0(ces_1_26_io_ins_0),
    .io_ins_1(ces_1_26_io_ins_1),
    .io_ins_2(ces_1_26_io_ins_2),
    .io_ins_3(ces_1_26_io_ins_3),
    .io_outs_0(ces_1_26_io_outs_0),
    .io_outs_1(ces_1_26_io_outs_1),
    .io_outs_2(ces_1_26_io_outs_2),
    .io_outs_3(ces_1_26_io_outs_3)
  );
  Element ces_1_27 ( // @[MockArray.scala 36:52]
    .clock(ces_1_27_clock),
    .io_ins_0(ces_1_27_io_ins_0),
    .io_ins_1(ces_1_27_io_ins_1),
    .io_ins_2(ces_1_27_io_ins_2),
    .io_ins_3(ces_1_27_io_ins_3),
    .io_outs_0(ces_1_27_io_outs_0),
    .io_outs_1(ces_1_27_io_outs_1),
    .io_outs_2(ces_1_27_io_outs_2),
    .io_outs_3(ces_1_27_io_outs_3)
  );
  Element ces_1_28 ( // @[MockArray.scala 36:52]
    .clock(ces_1_28_clock),
    .io_ins_0(ces_1_28_io_ins_0),
    .io_ins_1(ces_1_28_io_ins_1),
    .io_ins_2(ces_1_28_io_ins_2),
    .io_ins_3(ces_1_28_io_ins_3),
    .io_outs_0(ces_1_28_io_outs_0),
    .io_outs_1(ces_1_28_io_outs_1),
    .io_outs_2(ces_1_28_io_outs_2),
    .io_outs_3(ces_1_28_io_outs_3)
  );
  Element ces_1_29 ( // @[MockArray.scala 36:52]
    .clock(ces_1_29_clock),
    .io_ins_0(ces_1_29_io_ins_0),
    .io_ins_1(ces_1_29_io_ins_1),
    .io_ins_2(ces_1_29_io_ins_2),
    .io_ins_3(ces_1_29_io_ins_3),
    .io_outs_0(ces_1_29_io_outs_0),
    .io_outs_1(ces_1_29_io_outs_1),
    .io_outs_2(ces_1_29_io_outs_2),
    .io_outs_3(ces_1_29_io_outs_3)
  );
  Element ces_1_30 ( // @[MockArray.scala 36:52]
    .clock(ces_1_30_clock),
    .io_ins_0(ces_1_30_io_ins_0),
    .io_ins_1(ces_1_30_io_ins_1),
    .io_ins_2(ces_1_30_io_ins_2),
    .io_ins_3(ces_1_30_io_ins_3),
    .io_outs_0(ces_1_30_io_outs_0),
    .io_outs_1(ces_1_30_io_outs_1),
    .io_outs_2(ces_1_30_io_outs_2),
    .io_outs_3(ces_1_30_io_outs_3)
  );
  Element ces_1_31 ( // @[MockArray.scala 36:52]
    .clock(ces_1_31_clock),
    .io_ins_0(ces_1_31_io_ins_0),
    .io_ins_1(ces_1_31_io_ins_1),
    .io_ins_2(ces_1_31_io_ins_2),
    .io_ins_3(ces_1_31_io_ins_3),
    .io_outs_0(ces_1_31_io_outs_0),
    .io_outs_1(ces_1_31_io_outs_1),
    .io_outs_2(ces_1_31_io_outs_2),
    .io_outs_3(ces_1_31_io_outs_3)
  );
  Element ces_2_0 ( // @[MockArray.scala 36:52]
    .clock(ces_2_0_clock),
    .io_ins_0(ces_2_0_io_ins_0),
    .io_ins_1(ces_2_0_io_ins_1),
    .io_ins_2(ces_2_0_io_ins_2),
    .io_ins_3(ces_2_0_io_ins_3),
    .io_outs_0(ces_2_0_io_outs_0),
    .io_outs_1(ces_2_0_io_outs_1),
    .io_outs_2(ces_2_0_io_outs_2),
    .io_outs_3(ces_2_0_io_outs_3)
  );
  Element ces_2_1 ( // @[MockArray.scala 36:52]
    .clock(ces_2_1_clock),
    .io_ins_0(ces_2_1_io_ins_0),
    .io_ins_1(ces_2_1_io_ins_1),
    .io_ins_2(ces_2_1_io_ins_2),
    .io_ins_3(ces_2_1_io_ins_3),
    .io_outs_0(ces_2_1_io_outs_0),
    .io_outs_1(ces_2_1_io_outs_1),
    .io_outs_2(ces_2_1_io_outs_2),
    .io_outs_3(ces_2_1_io_outs_3)
  );
  Element ces_2_2 ( // @[MockArray.scala 36:52]
    .clock(ces_2_2_clock),
    .io_ins_0(ces_2_2_io_ins_0),
    .io_ins_1(ces_2_2_io_ins_1),
    .io_ins_2(ces_2_2_io_ins_2),
    .io_ins_3(ces_2_2_io_ins_3),
    .io_outs_0(ces_2_2_io_outs_0),
    .io_outs_1(ces_2_2_io_outs_1),
    .io_outs_2(ces_2_2_io_outs_2),
    .io_outs_3(ces_2_2_io_outs_3)
  );
  Element ces_2_3 ( // @[MockArray.scala 36:52]
    .clock(ces_2_3_clock),
    .io_ins_0(ces_2_3_io_ins_0),
    .io_ins_1(ces_2_3_io_ins_1),
    .io_ins_2(ces_2_3_io_ins_2),
    .io_ins_3(ces_2_3_io_ins_3),
    .io_outs_0(ces_2_3_io_outs_0),
    .io_outs_1(ces_2_3_io_outs_1),
    .io_outs_2(ces_2_3_io_outs_2),
    .io_outs_3(ces_2_3_io_outs_3)
  );
  Element ces_2_4 ( // @[MockArray.scala 36:52]
    .clock(ces_2_4_clock),
    .io_ins_0(ces_2_4_io_ins_0),
    .io_ins_1(ces_2_4_io_ins_1),
    .io_ins_2(ces_2_4_io_ins_2),
    .io_ins_3(ces_2_4_io_ins_3),
    .io_outs_0(ces_2_4_io_outs_0),
    .io_outs_1(ces_2_4_io_outs_1),
    .io_outs_2(ces_2_4_io_outs_2),
    .io_outs_3(ces_2_4_io_outs_3)
  );
  Element ces_2_5 ( // @[MockArray.scala 36:52]
    .clock(ces_2_5_clock),
    .io_ins_0(ces_2_5_io_ins_0),
    .io_ins_1(ces_2_5_io_ins_1),
    .io_ins_2(ces_2_5_io_ins_2),
    .io_ins_3(ces_2_5_io_ins_3),
    .io_outs_0(ces_2_5_io_outs_0),
    .io_outs_1(ces_2_5_io_outs_1),
    .io_outs_2(ces_2_5_io_outs_2),
    .io_outs_3(ces_2_5_io_outs_3)
  );
  Element ces_2_6 ( // @[MockArray.scala 36:52]
    .clock(ces_2_6_clock),
    .io_ins_0(ces_2_6_io_ins_0),
    .io_ins_1(ces_2_6_io_ins_1),
    .io_ins_2(ces_2_6_io_ins_2),
    .io_ins_3(ces_2_6_io_ins_3),
    .io_outs_0(ces_2_6_io_outs_0),
    .io_outs_1(ces_2_6_io_outs_1),
    .io_outs_2(ces_2_6_io_outs_2),
    .io_outs_3(ces_2_6_io_outs_3)
  );
  Element ces_2_7 ( // @[MockArray.scala 36:52]
    .clock(ces_2_7_clock),
    .io_ins_0(ces_2_7_io_ins_0),
    .io_ins_1(ces_2_7_io_ins_1),
    .io_ins_2(ces_2_7_io_ins_2),
    .io_ins_3(ces_2_7_io_ins_3),
    .io_outs_0(ces_2_7_io_outs_0),
    .io_outs_1(ces_2_7_io_outs_1),
    .io_outs_2(ces_2_7_io_outs_2),
    .io_outs_3(ces_2_7_io_outs_3)
  );
  Element ces_2_8 ( // @[MockArray.scala 36:52]
    .clock(ces_2_8_clock),
    .io_ins_0(ces_2_8_io_ins_0),
    .io_ins_1(ces_2_8_io_ins_1),
    .io_ins_2(ces_2_8_io_ins_2),
    .io_ins_3(ces_2_8_io_ins_3),
    .io_outs_0(ces_2_8_io_outs_0),
    .io_outs_1(ces_2_8_io_outs_1),
    .io_outs_2(ces_2_8_io_outs_2),
    .io_outs_3(ces_2_8_io_outs_3)
  );
  Element ces_2_9 ( // @[MockArray.scala 36:52]
    .clock(ces_2_9_clock),
    .io_ins_0(ces_2_9_io_ins_0),
    .io_ins_1(ces_2_9_io_ins_1),
    .io_ins_2(ces_2_9_io_ins_2),
    .io_ins_3(ces_2_9_io_ins_3),
    .io_outs_0(ces_2_9_io_outs_0),
    .io_outs_1(ces_2_9_io_outs_1),
    .io_outs_2(ces_2_9_io_outs_2),
    .io_outs_3(ces_2_9_io_outs_3)
  );
  Element ces_2_10 ( // @[MockArray.scala 36:52]
    .clock(ces_2_10_clock),
    .io_ins_0(ces_2_10_io_ins_0),
    .io_ins_1(ces_2_10_io_ins_1),
    .io_ins_2(ces_2_10_io_ins_2),
    .io_ins_3(ces_2_10_io_ins_3),
    .io_outs_0(ces_2_10_io_outs_0),
    .io_outs_1(ces_2_10_io_outs_1),
    .io_outs_2(ces_2_10_io_outs_2),
    .io_outs_3(ces_2_10_io_outs_3)
  );
  Element ces_2_11 ( // @[MockArray.scala 36:52]
    .clock(ces_2_11_clock),
    .io_ins_0(ces_2_11_io_ins_0),
    .io_ins_1(ces_2_11_io_ins_1),
    .io_ins_2(ces_2_11_io_ins_2),
    .io_ins_3(ces_2_11_io_ins_3),
    .io_outs_0(ces_2_11_io_outs_0),
    .io_outs_1(ces_2_11_io_outs_1),
    .io_outs_2(ces_2_11_io_outs_2),
    .io_outs_3(ces_2_11_io_outs_3)
  );
  Element ces_2_12 ( // @[MockArray.scala 36:52]
    .clock(ces_2_12_clock),
    .io_ins_0(ces_2_12_io_ins_0),
    .io_ins_1(ces_2_12_io_ins_1),
    .io_ins_2(ces_2_12_io_ins_2),
    .io_ins_3(ces_2_12_io_ins_3),
    .io_outs_0(ces_2_12_io_outs_0),
    .io_outs_1(ces_2_12_io_outs_1),
    .io_outs_2(ces_2_12_io_outs_2),
    .io_outs_3(ces_2_12_io_outs_3)
  );
  Element ces_2_13 ( // @[MockArray.scala 36:52]
    .clock(ces_2_13_clock),
    .io_ins_0(ces_2_13_io_ins_0),
    .io_ins_1(ces_2_13_io_ins_1),
    .io_ins_2(ces_2_13_io_ins_2),
    .io_ins_3(ces_2_13_io_ins_3),
    .io_outs_0(ces_2_13_io_outs_0),
    .io_outs_1(ces_2_13_io_outs_1),
    .io_outs_2(ces_2_13_io_outs_2),
    .io_outs_3(ces_2_13_io_outs_3)
  );
  Element ces_2_14 ( // @[MockArray.scala 36:52]
    .clock(ces_2_14_clock),
    .io_ins_0(ces_2_14_io_ins_0),
    .io_ins_1(ces_2_14_io_ins_1),
    .io_ins_2(ces_2_14_io_ins_2),
    .io_ins_3(ces_2_14_io_ins_3),
    .io_outs_0(ces_2_14_io_outs_0),
    .io_outs_1(ces_2_14_io_outs_1),
    .io_outs_2(ces_2_14_io_outs_2),
    .io_outs_3(ces_2_14_io_outs_3)
  );
  Element ces_2_15 ( // @[MockArray.scala 36:52]
    .clock(ces_2_15_clock),
    .io_ins_0(ces_2_15_io_ins_0),
    .io_ins_1(ces_2_15_io_ins_1),
    .io_ins_2(ces_2_15_io_ins_2),
    .io_ins_3(ces_2_15_io_ins_3),
    .io_outs_0(ces_2_15_io_outs_0),
    .io_outs_1(ces_2_15_io_outs_1),
    .io_outs_2(ces_2_15_io_outs_2),
    .io_outs_3(ces_2_15_io_outs_3)
  );
  Element ces_2_16 ( // @[MockArray.scala 36:52]
    .clock(ces_2_16_clock),
    .io_ins_0(ces_2_16_io_ins_0),
    .io_ins_1(ces_2_16_io_ins_1),
    .io_ins_2(ces_2_16_io_ins_2),
    .io_ins_3(ces_2_16_io_ins_3),
    .io_outs_0(ces_2_16_io_outs_0),
    .io_outs_1(ces_2_16_io_outs_1),
    .io_outs_2(ces_2_16_io_outs_2),
    .io_outs_3(ces_2_16_io_outs_3)
  );
  Element ces_2_17 ( // @[MockArray.scala 36:52]
    .clock(ces_2_17_clock),
    .io_ins_0(ces_2_17_io_ins_0),
    .io_ins_1(ces_2_17_io_ins_1),
    .io_ins_2(ces_2_17_io_ins_2),
    .io_ins_3(ces_2_17_io_ins_3),
    .io_outs_0(ces_2_17_io_outs_0),
    .io_outs_1(ces_2_17_io_outs_1),
    .io_outs_2(ces_2_17_io_outs_2),
    .io_outs_3(ces_2_17_io_outs_3)
  );
  Element ces_2_18 ( // @[MockArray.scala 36:52]
    .clock(ces_2_18_clock),
    .io_ins_0(ces_2_18_io_ins_0),
    .io_ins_1(ces_2_18_io_ins_1),
    .io_ins_2(ces_2_18_io_ins_2),
    .io_ins_3(ces_2_18_io_ins_3),
    .io_outs_0(ces_2_18_io_outs_0),
    .io_outs_1(ces_2_18_io_outs_1),
    .io_outs_2(ces_2_18_io_outs_2),
    .io_outs_3(ces_2_18_io_outs_3)
  );
  Element ces_2_19 ( // @[MockArray.scala 36:52]
    .clock(ces_2_19_clock),
    .io_ins_0(ces_2_19_io_ins_0),
    .io_ins_1(ces_2_19_io_ins_1),
    .io_ins_2(ces_2_19_io_ins_2),
    .io_ins_3(ces_2_19_io_ins_3),
    .io_outs_0(ces_2_19_io_outs_0),
    .io_outs_1(ces_2_19_io_outs_1),
    .io_outs_2(ces_2_19_io_outs_2),
    .io_outs_3(ces_2_19_io_outs_3)
  );
  Element ces_2_20 ( // @[MockArray.scala 36:52]
    .clock(ces_2_20_clock),
    .io_ins_0(ces_2_20_io_ins_0),
    .io_ins_1(ces_2_20_io_ins_1),
    .io_ins_2(ces_2_20_io_ins_2),
    .io_ins_3(ces_2_20_io_ins_3),
    .io_outs_0(ces_2_20_io_outs_0),
    .io_outs_1(ces_2_20_io_outs_1),
    .io_outs_2(ces_2_20_io_outs_2),
    .io_outs_3(ces_2_20_io_outs_3)
  );
  Element ces_2_21 ( // @[MockArray.scala 36:52]
    .clock(ces_2_21_clock),
    .io_ins_0(ces_2_21_io_ins_0),
    .io_ins_1(ces_2_21_io_ins_1),
    .io_ins_2(ces_2_21_io_ins_2),
    .io_ins_3(ces_2_21_io_ins_3),
    .io_outs_0(ces_2_21_io_outs_0),
    .io_outs_1(ces_2_21_io_outs_1),
    .io_outs_2(ces_2_21_io_outs_2),
    .io_outs_3(ces_2_21_io_outs_3)
  );
  Element ces_2_22 ( // @[MockArray.scala 36:52]
    .clock(ces_2_22_clock),
    .io_ins_0(ces_2_22_io_ins_0),
    .io_ins_1(ces_2_22_io_ins_1),
    .io_ins_2(ces_2_22_io_ins_2),
    .io_ins_3(ces_2_22_io_ins_3),
    .io_outs_0(ces_2_22_io_outs_0),
    .io_outs_1(ces_2_22_io_outs_1),
    .io_outs_2(ces_2_22_io_outs_2),
    .io_outs_3(ces_2_22_io_outs_3)
  );
  Element ces_2_23 ( // @[MockArray.scala 36:52]
    .clock(ces_2_23_clock),
    .io_ins_0(ces_2_23_io_ins_0),
    .io_ins_1(ces_2_23_io_ins_1),
    .io_ins_2(ces_2_23_io_ins_2),
    .io_ins_3(ces_2_23_io_ins_3),
    .io_outs_0(ces_2_23_io_outs_0),
    .io_outs_1(ces_2_23_io_outs_1),
    .io_outs_2(ces_2_23_io_outs_2),
    .io_outs_3(ces_2_23_io_outs_3)
  );
  Element ces_2_24 ( // @[MockArray.scala 36:52]
    .clock(ces_2_24_clock),
    .io_ins_0(ces_2_24_io_ins_0),
    .io_ins_1(ces_2_24_io_ins_1),
    .io_ins_2(ces_2_24_io_ins_2),
    .io_ins_3(ces_2_24_io_ins_3),
    .io_outs_0(ces_2_24_io_outs_0),
    .io_outs_1(ces_2_24_io_outs_1),
    .io_outs_2(ces_2_24_io_outs_2),
    .io_outs_3(ces_2_24_io_outs_3)
  );
  Element ces_2_25 ( // @[MockArray.scala 36:52]
    .clock(ces_2_25_clock),
    .io_ins_0(ces_2_25_io_ins_0),
    .io_ins_1(ces_2_25_io_ins_1),
    .io_ins_2(ces_2_25_io_ins_2),
    .io_ins_3(ces_2_25_io_ins_3),
    .io_outs_0(ces_2_25_io_outs_0),
    .io_outs_1(ces_2_25_io_outs_1),
    .io_outs_2(ces_2_25_io_outs_2),
    .io_outs_3(ces_2_25_io_outs_3)
  );
  Element ces_2_26 ( // @[MockArray.scala 36:52]
    .clock(ces_2_26_clock),
    .io_ins_0(ces_2_26_io_ins_0),
    .io_ins_1(ces_2_26_io_ins_1),
    .io_ins_2(ces_2_26_io_ins_2),
    .io_ins_3(ces_2_26_io_ins_3),
    .io_outs_0(ces_2_26_io_outs_0),
    .io_outs_1(ces_2_26_io_outs_1),
    .io_outs_2(ces_2_26_io_outs_2),
    .io_outs_3(ces_2_26_io_outs_3)
  );
  Element ces_2_27 ( // @[MockArray.scala 36:52]
    .clock(ces_2_27_clock),
    .io_ins_0(ces_2_27_io_ins_0),
    .io_ins_1(ces_2_27_io_ins_1),
    .io_ins_2(ces_2_27_io_ins_2),
    .io_ins_3(ces_2_27_io_ins_3),
    .io_outs_0(ces_2_27_io_outs_0),
    .io_outs_1(ces_2_27_io_outs_1),
    .io_outs_2(ces_2_27_io_outs_2),
    .io_outs_3(ces_2_27_io_outs_3)
  );
  Element ces_2_28 ( // @[MockArray.scala 36:52]
    .clock(ces_2_28_clock),
    .io_ins_0(ces_2_28_io_ins_0),
    .io_ins_1(ces_2_28_io_ins_1),
    .io_ins_2(ces_2_28_io_ins_2),
    .io_ins_3(ces_2_28_io_ins_3),
    .io_outs_0(ces_2_28_io_outs_0),
    .io_outs_1(ces_2_28_io_outs_1),
    .io_outs_2(ces_2_28_io_outs_2),
    .io_outs_3(ces_2_28_io_outs_3)
  );
  Element ces_2_29 ( // @[MockArray.scala 36:52]
    .clock(ces_2_29_clock),
    .io_ins_0(ces_2_29_io_ins_0),
    .io_ins_1(ces_2_29_io_ins_1),
    .io_ins_2(ces_2_29_io_ins_2),
    .io_ins_3(ces_2_29_io_ins_3),
    .io_outs_0(ces_2_29_io_outs_0),
    .io_outs_1(ces_2_29_io_outs_1),
    .io_outs_2(ces_2_29_io_outs_2),
    .io_outs_3(ces_2_29_io_outs_3)
  );
  Element ces_2_30 ( // @[MockArray.scala 36:52]
    .clock(ces_2_30_clock),
    .io_ins_0(ces_2_30_io_ins_0),
    .io_ins_1(ces_2_30_io_ins_1),
    .io_ins_2(ces_2_30_io_ins_2),
    .io_ins_3(ces_2_30_io_ins_3),
    .io_outs_0(ces_2_30_io_outs_0),
    .io_outs_1(ces_2_30_io_outs_1),
    .io_outs_2(ces_2_30_io_outs_2),
    .io_outs_3(ces_2_30_io_outs_3)
  );
  Element ces_2_31 ( // @[MockArray.scala 36:52]
    .clock(ces_2_31_clock),
    .io_ins_0(ces_2_31_io_ins_0),
    .io_ins_1(ces_2_31_io_ins_1),
    .io_ins_2(ces_2_31_io_ins_2),
    .io_ins_3(ces_2_31_io_ins_3),
    .io_outs_0(ces_2_31_io_outs_0),
    .io_outs_1(ces_2_31_io_outs_1),
    .io_outs_2(ces_2_31_io_outs_2),
    .io_outs_3(ces_2_31_io_outs_3)
  );
  Element ces_3_0 ( // @[MockArray.scala 36:52]
    .clock(ces_3_0_clock),
    .io_ins_0(ces_3_0_io_ins_0),
    .io_ins_1(ces_3_0_io_ins_1),
    .io_ins_2(ces_3_0_io_ins_2),
    .io_ins_3(ces_3_0_io_ins_3),
    .io_outs_0(ces_3_0_io_outs_0),
    .io_outs_1(ces_3_0_io_outs_1),
    .io_outs_2(ces_3_0_io_outs_2),
    .io_outs_3(ces_3_0_io_outs_3)
  );
  Element ces_3_1 ( // @[MockArray.scala 36:52]
    .clock(ces_3_1_clock),
    .io_ins_0(ces_3_1_io_ins_0),
    .io_ins_1(ces_3_1_io_ins_1),
    .io_ins_2(ces_3_1_io_ins_2),
    .io_ins_3(ces_3_1_io_ins_3),
    .io_outs_0(ces_3_1_io_outs_0),
    .io_outs_1(ces_3_1_io_outs_1),
    .io_outs_2(ces_3_1_io_outs_2),
    .io_outs_3(ces_3_1_io_outs_3)
  );
  Element ces_3_2 ( // @[MockArray.scala 36:52]
    .clock(ces_3_2_clock),
    .io_ins_0(ces_3_2_io_ins_0),
    .io_ins_1(ces_3_2_io_ins_1),
    .io_ins_2(ces_3_2_io_ins_2),
    .io_ins_3(ces_3_2_io_ins_3),
    .io_outs_0(ces_3_2_io_outs_0),
    .io_outs_1(ces_3_2_io_outs_1),
    .io_outs_2(ces_3_2_io_outs_2),
    .io_outs_3(ces_3_2_io_outs_3)
  );
  Element ces_3_3 ( // @[MockArray.scala 36:52]
    .clock(ces_3_3_clock),
    .io_ins_0(ces_3_3_io_ins_0),
    .io_ins_1(ces_3_3_io_ins_1),
    .io_ins_2(ces_3_3_io_ins_2),
    .io_ins_3(ces_3_3_io_ins_3),
    .io_outs_0(ces_3_3_io_outs_0),
    .io_outs_1(ces_3_3_io_outs_1),
    .io_outs_2(ces_3_3_io_outs_2),
    .io_outs_3(ces_3_3_io_outs_3)
  );
  Element ces_3_4 ( // @[MockArray.scala 36:52]
    .clock(ces_3_4_clock),
    .io_ins_0(ces_3_4_io_ins_0),
    .io_ins_1(ces_3_4_io_ins_1),
    .io_ins_2(ces_3_4_io_ins_2),
    .io_ins_3(ces_3_4_io_ins_3),
    .io_outs_0(ces_3_4_io_outs_0),
    .io_outs_1(ces_3_4_io_outs_1),
    .io_outs_2(ces_3_4_io_outs_2),
    .io_outs_3(ces_3_4_io_outs_3)
  );
  Element ces_3_5 ( // @[MockArray.scala 36:52]
    .clock(ces_3_5_clock),
    .io_ins_0(ces_3_5_io_ins_0),
    .io_ins_1(ces_3_5_io_ins_1),
    .io_ins_2(ces_3_5_io_ins_2),
    .io_ins_3(ces_3_5_io_ins_3),
    .io_outs_0(ces_3_5_io_outs_0),
    .io_outs_1(ces_3_5_io_outs_1),
    .io_outs_2(ces_3_5_io_outs_2),
    .io_outs_3(ces_3_5_io_outs_3)
  );
  Element ces_3_6 ( // @[MockArray.scala 36:52]
    .clock(ces_3_6_clock),
    .io_ins_0(ces_3_6_io_ins_0),
    .io_ins_1(ces_3_6_io_ins_1),
    .io_ins_2(ces_3_6_io_ins_2),
    .io_ins_3(ces_3_6_io_ins_3),
    .io_outs_0(ces_3_6_io_outs_0),
    .io_outs_1(ces_3_6_io_outs_1),
    .io_outs_2(ces_3_6_io_outs_2),
    .io_outs_3(ces_3_6_io_outs_3)
  );
  Element ces_3_7 ( // @[MockArray.scala 36:52]
    .clock(ces_3_7_clock),
    .io_ins_0(ces_3_7_io_ins_0),
    .io_ins_1(ces_3_7_io_ins_1),
    .io_ins_2(ces_3_7_io_ins_2),
    .io_ins_3(ces_3_7_io_ins_3),
    .io_outs_0(ces_3_7_io_outs_0),
    .io_outs_1(ces_3_7_io_outs_1),
    .io_outs_2(ces_3_7_io_outs_2),
    .io_outs_3(ces_3_7_io_outs_3)
  );
  Element ces_3_8 ( // @[MockArray.scala 36:52]
    .clock(ces_3_8_clock),
    .io_ins_0(ces_3_8_io_ins_0),
    .io_ins_1(ces_3_8_io_ins_1),
    .io_ins_2(ces_3_8_io_ins_2),
    .io_ins_3(ces_3_8_io_ins_3),
    .io_outs_0(ces_3_8_io_outs_0),
    .io_outs_1(ces_3_8_io_outs_1),
    .io_outs_2(ces_3_8_io_outs_2),
    .io_outs_3(ces_3_8_io_outs_3)
  );
  Element ces_3_9 ( // @[MockArray.scala 36:52]
    .clock(ces_3_9_clock),
    .io_ins_0(ces_3_9_io_ins_0),
    .io_ins_1(ces_3_9_io_ins_1),
    .io_ins_2(ces_3_9_io_ins_2),
    .io_ins_3(ces_3_9_io_ins_3),
    .io_outs_0(ces_3_9_io_outs_0),
    .io_outs_1(ces_3_9_io_outs_1),
    .io_outs_2(ces_3_9_io_outs_2),
    .io_outs_3(ces_3_9_io_outs_3)
  );
  Element ces_3_10 ( // @[MockArray.scala 36:52]
    .clock(ces_3_10_clock),
    .io_ins_0(ces_3_10_io_ins_0),
    .io_ins_1(ces_3_10_io_ins_1),
    .io_ins_2(ces_3_10_io_ins_2),
    .io_ins_3(ces_3_10_io_ins_3),
    .io_outs_0(ces_3_10_io_outs_0),
    .io_outs_1(ces_3_10_io_outs_1),
    .io_outs_2(ces_3_10_io_outs_2),
    .io_outs_3(ces_3_10_io_outs_3)
  );
  Element ces_3_11 ( // @[MockArray.scala 36:52]
    .clock(ces_3_11_clock),
    .io_ins_0(ces_3_11_io_ins_0),
    .io_ins_1(ces_3_11_io_ins_1),
    .io_ins_2(ces_3_11_io_ins_2),
    .io_ins_3(ces_3_11_io_ins_3),
    .io_outs_0(ces_3_11_io_outs_0),
    .io_outs_1(ces_3_11_io_outs_1),
    .io_outs_2(ces_3_11_io_outs_2),
    .io_outs_3(ces_3_11_io_outs_3)
  );
  Element ces_3_12 ( // @[MockArray.scala 36:52]
    .clock(ces_3_12_clock),
    .io_ins_0(ces_3_12_io_ins_0),
    .io_ins_1(ces_3_12_io_ins_1),
    .io_ins_2(ces_3_12_io_ins_2),
    .io_ins_3(ces_3_12_io_ins_3),
    .io_outs_0(ces_3_12_io_outs_0),
    .io_outs_1(ces_3_12_io_outs_1),
    .io_outs_2(ces_3_12_io_outs_2),
    .io_outs_3(ces_3_12_io_outs_3)
  );
  Element ces_3_13 ( // @[MockArray.scala 36:52]
    .clock(ces_3_13_clock),
    .io_ins_0(ces_3_13_io_ins_0),
    .io_ins_1(ces_3_13_io_ins_1),
    .io_ins_2(ces_3_13_io_ins_2),
    .io_ins_3(ces_3_13_io_ins_3),
    .io_outs_0(ces_3_13_io_outs_0),
    .io_outs_1(ces_3_13_io_outs_1),
    .io_outs_2(ces_3_13_io_outs_2),
    .io_outs_3(ces_3_13_io_outs_3)
  );
  Element ces_3_14 ( // @[MockArray.scala 36:52]
    .clock(ces_3_14_clock),
    .io_ins_0(ces_3_14_io_ins_0),
    .io_ins_1(ces_3_14_io_ins_1),
    .io_ins_2(ces_3_14_io_ins_2),
    .io_ins_3(ces_3_14_io_ins_3),
    .io_outs_0(ces_3_14_io_outs_0),
    .io_outs_1(ces_3_14_io_outs_1),
    .io_outs_2(ces_3_14_io_outs_2),
    .io_outs_3(ces_3_14_io_outs_3)
  );
  Element ces_3_15 ( // @[MockArray.scala 36:52]
    .clock(ces_3_15_clock),
    .io_ins_0(ces_3_15_io_ins_0),
    .io_ins_1(ces_3_15_io_ins_1),
    .io_ins_2(ces_3_15_io_ins_2),
    .io_ins_3(ces_3_15_io_ins_3),
    .io_outs_0(ces_3_15_io_outs_0),
    .io_outs_1(ces_3_15_io_outs_1),
    .io_outs_2(ces_3_15_io_outs_2),
    .io_outs_3(ces_3_15_io_outs_3)
  );
  Element ces_3_16 ( // @[MockArray.scala 36:52]
    .clock(ces_3_16_clock),
    .io_ins_0(ces_3_16_io_ins_0),
    .io_ins_1(ces_3_16_io_ins_1),
    .io_ins_2(ces_3_16_io_ins_2),
    .io_ins_3(ces_3_16_io_ins_3),
    .io_outs_0(ces_3_16_io_outs_0),
    .io_outs_1(ces_3_16_io_outs_1),
    .io_outs_2(ces_3_16_io_outs_2),
    .io_outs_3(ces_3_16_io_outs_3)
  );
  Element ces_3_17 ( // @[MockArray.scala 36:52]
    .clock(ces_3_17_clock),
    .io_ins_0(ces_3_17_io_ins_0),
    .io_ins_1(ces_3_17_io_ins_1),
    .io_ins_2(ces_3_17_io_ins_2),
    .io_ins_3(ces_3_17_io_ins_3),
    .io_outs_0(ces_3_17_io_outs_0),
    .io_outs_1(ces_3_17_io_outs_1),
    .io_outs_2(ces_3_17_io_outs_2),
    .io_outs_3(ces_3_17_io_outs_3)
  );
  Element ces_3_18 ( // @[MockArray.scala 36:52]
    .clock(ces_3_18_clock),
    .io_ins_0(ces_3_18_io_ins_0),
    .io_ins_1(ces_3_18_io_ins_1),
    .io_ins_2(ces_3_18_io_ins_2),
    .io_ins_3(ces_3_18_io_ins_3),
    .io_outs_0(ces_3_18_io_outs_0),
    .io_outs_1(ces_3_18_io_outs_1),
    .io_outs_2(ces_3_18_io_outs_2),
    .io_outs_3(ces_3_18_io_outs_3)
  );
  Element ces_3_19 ( // @[MockArray.scala 36:52]
    .clock(ces_3_19_clock),
    .io_ins_0(ces_3_19_io_ins_0),
    .io_ins_1(ces_3_19_io_ins_1),
    .io_ins_2(ces_3_19_io_ins_2),
    .io_ins_3(ces_3_19_io_ins_3),
    .io_outs_0(ces_3_19_io_outs_0),
    .io_outs_1(ces_3_19_io_outs_1),
    .io_outs_2(ces_3_19_io_outs_2),
    .io_outs_3(ces_3_19_io_outs_3)
  );
  Element ces_3_20 ( // @[MockArray.scala 36:52]
    .clock(ces_3_20_clock),
    .io_ins_0(ces_3_20_io_ins_0),
    .io_ins_1(ces_3_20_io_ins_1),
    .io_ins_2(ces_3_20_io_ins_2),
    .io_ins_3(ces_3_20_io_ins_3),
    .io_outs_0(ces_3_20_io_outs_0),
    .io_outs_1(ces_3_20_io_outs_1),
    .io_outs_2(ces_3_20_io_outs_2),
    .io_outs_3(ces_3_20_io_outs_3)
  );
  Element ces_3_21 ( // @[MockArray.scala 36:52]
    .clock(ces_3_21_clock),
    .io_ins_0(ces_3_21_io_ins_0),
    .io_ins_1(ces_3_21_io_ins_1),
    .io_ins_2(ces_3_21_io_ins_2),
    .io_ins_3(ces_3_21_io_ins_3),
    .io_outs_0(ces_3_21_io_outs_0),
    .io_outs_1(ces_3_21_io_outs_1),
    .io_outs_2(ces_3_21_io_outs_2),
    .io_outs_3(ces_3_21_io_outs_3)
  );
  Element ces_3_22 ( // @[MockArray.scala 36:52]
    .clock(ces_3_22_clock),
    .io_ins_0(ces_3_22_io_ins_0),
    .io_ins_1(ces_3_22_io_ins_1),
    .io_ins_2(ces_3_22_io_ins_2),
    .io_ins_3(ces_3_22_io_ins_3),
    .io_outs_0(ces_3_22_io_outs_0),
    .io_outs_1(ces_3_22_io_outs_1),
    .io_outs_2(ces_3_22_io_outs_2),
    .io_outs_3(ces_3_22_io_outs_3)
  );
  Element ces_3_23 ( // @[MockArray.scala 36:52]
    .clock(ces_3_23_clock),
    .io_ins_0(ces_3_23_io_ins_0),
    .io_ins_1(ces_3_23_io_ins_1),
    .io_ins_2(ces_3_23_io_ins_2),
    .io_ins_3(ces_3_23_io_ins_3),
    .io_outs_0(ces_3_23_io_outs_0),
    .io_outs_1(ces_3_23_io_outs_1),
    .io_outs_2(ces_3_23_io_outs_2),
    .io_outs_3(ces_3_23_io_outs_3)
  );
  Element ces_3_24 ( // @[MockArray.scala 36:52]
    .clock(ces_3_24_clock),
    .io_ins_0(ces_3_24_io_ins_0),
    .io_ins_1(ces_3_24_io_ins_1),
    .io_ins_2(ces_3_24_io_ins_2),
    .io_ins_3(ces_3_24_io_ins_3),
    .io_outs_0(ces_3_24_io_outs_0),
    .io_outs_1(ces_3_24_io_outs_1),
    .io_outs_2(ces_3_24_io_outs_2),
    .io_outs_3(ces_3_24_io_outs_3)
  );
  Element ces_3_25 ( // @[MockArray.scala 36:52]
    .clock(ces_3_25_clock),
    .io_ins_0(ces_3_25_io_ins_0),
    .io_ins_1(ces_3_25_io_ins_1),
    .io_ins_2(ces_3_25_io_ins_2),
    .io_ins_3(ces_3_25_io_ins_3),
    .io_outs_0(ces_3_25_io_outs_0),
    .io_outs_1(ces_3_25_io_outs_1),
    .io_outs_2(ces_3_25_io_outs_2),
    .io_outs_3(ces_3_25_io_outs_3)
  );
  Element ces_3_26 ( // @[MockArray.scala 36:52]
    .clock(ces_3_26_clock),
    .io_ins_0(ces_3_26_io_ins_0),
    .io_ins_1(ces_3_26_io_ins_1),
    .io_ins_2(ces_3_26_io_ins_2),
    .io_ins_3(ces_3_26_io_ins_3),
    .io_outs_0(ces_3_26_io_outs_0),
    .io_outs_1(ces_3_26_io_outs_1),
    .io_outs_2(ces_3_26_io_outs_2),
    .io_outs_3(ces_3_26_io_outs_3)
  );
  Element ces_3_27 ( // @[MockArray.scala 36:52]
    .clock(ces_3_27_clock),
    .io_ins_0(ces_3_27_io_ins_0),
    .io_ins_1(ces_3_27_io_ins_1),
    .io_ins_2(ces_3_27_io_ins_2),
    .io_ins_3(ces_3_27_io_ins_3),
    .io_outs_0(ces_3_27_io_outs_0),
    .io_outs_1(ces_3_27_io_outs_1),
    .io_outs_2(ces_3_27_io_outs_2),
    .io_outs_3(ces_3_27_io_outs_3)
  );
  Element ces_3_28 ( // @[MockArray.scala 36:52]
    .clock(ces_3_28_clock),
    .io_ins_0(ces_3_28_io_ins_0),
    .io_ins_1(ces_3_28_io_ins_1),
    .io_ins_2(ces_3_28_io_ins_2),
    .io_ins_3(ces_3_28_io_ins_3),
    .io_outs_0(ces_3_28_io_outs_0),
    .io_outs_1(ces_3_28_io_outs_1),
    .io_outs_2(ces_3_28_io_outs_2),
    .io_outs_3(ces_3_28_io_outs_3)
  );
  Element ces_3_29 ( // @[MockArray.scala 36:52]
    .clock(ces_3_29_clock),
    .io_ins_0(ces_3_29_io_ins_0),
    .io_ins_1(ces_3_29_io_ins_1),
    .io_ins_2(ces_3_29_io_ins_2),
    .io_ins_3(ces_3_29_io_ins_3),
    .io_outs_0(ces_3_29_io_outs_0),
    .io_outs_1(ces_3_29_io_outs_1),
    .io_outs_2(ces_3_29_io_outs_2),
    .io_outs_3(ces_3_29_io_outs_3)
  );
  Element ces_3_30 ( // @[MockArray.scala 36:52]
    .clock(ces_3_30_clock),
    .io_ins_0(ces_3_30_io_ins_0),
    .io_ins_1(ces_3_30_io_ins_1),
    .io_ins_2(ces_3_30_io_ins_2),
    .io_ins_3(ces_3_30_io_ins_3),
    .io_outs_0(ces_3_30_io_outs_0),
    .io_outs_1(ces_3_30_io_outs_1),
    .io_outs_2(ces_3_30_io_outs_2),
    .io_outs_3(ces_3_30_io_outs_3)
  );
  Element ces_3_31 ( // @[MockArray.scala 36:52]
    .clock(ces_3_31_clock),
    .io_ins_0(ces_3_31_io_ins_0),
    .io_ins_1(ces_3_31_io_ins_1),
    .io_ins_2(ces_3_31_io_ins_2),
    .io_ins_3(ces_3_31_io_ins_3),
    .io_outs_0(ces_3_31_io_outs_0),
    .io_outs_1(ces_3_31_io_outs_1),
    .io_outs_2(ces_3_31_io_outs_2),
    .io_outs_3(ces_3_31_io_outs_3)
  );
  Element ces_4_0 ( // @[MockArray.scala 36:52]
    .clock(ces_4_0_clock),
    .io_ins_0(ces_4_0_io_ins_0),
    .io_ins_1(ces_4_0_io_ins_1),
    .io_ins_2(ces_4_0_io_ins_2),
    .io_ins_3(ces_4_0_io_ins_3),
    .io_outs_0(ces_4_0_io_outs_0),
    .io_outs_1(ces_4_0_io_outs_1),
    .io_outs_2(ces_4_0_io_outs_2),
    .io_outs_3(ces_4_0_io_outs_3)
  );
  Element ces_4_1 ( // @[MockArray.scala 36:52]
    .clock(ces_4_1_clock),
    .io_ins_0(ces_4_1_io_ins_0),
    .io_ins_1(ces_4_1_io_ins_1),
    .io_ins_2(ces_4_1_io_ins_2),
    .io_ins_3(ces_4_1_io_ins_3),
    .io_outs_0(ces_4_1_io_outs_0),
    .io_outs_1(ces_4_1_io_outs_1),
    .io_outs_2(ces_4_1_io_outs_2),
    .io_outs_3(ces_4_1_io_outs_3)
  );
  Element ces_4_2 ( // @[MockArray.scala 36:52]
    .clock(ces_4_2_clock),
    .io_ins_0(ces_4_2_io_ins_0),
    .io_ins_1(ces_4_2_io_ins_1),
    .io_ins_2(ces_4_2_io_ins_2),
    .io_ins_3(ces_4_2_io_ins_3),
    .io_outs_0(ces_4_2_io_outs_0),
    .io_outs_1(ces_4_2_io_outs_1),
    .io_outs_2(ces_4_2_io_outs_2),
    .io_outs_3(ces_4_2_io_outs_3)
  );
  Element ces_4_3 ( // @[MockArray.scala 36:52]
    .clock(ces_4_3_clock),
    .io_ins_0(ces_4_3_io_ins_0),
    .io_ins_1(ces_4_3_io_ins_1),
    .io_ins_2(ces_4_3_io_ins_2),
    .io_ins_3(ces_4_3_io_ins_3),
    .io_outs_0(ces_4_3_io_outs_0),
    .io_outs_1(ces_4_3_io_outs_1),
    .io_outs_2(ces_4_3_io_outs_2),
    .io_outs_3(ces_4_3_io_outs_3)
  );
  Element ces_4_4 ( // @[MockArray.scala 36:52]
    .clock(ces_4_4_clock),
    .io_ins_0(ces_4_4_io_ins_0),
    .io_ins_1(ces_4_4_io_ins_1),
    .io_ins_2(ces_4_4_io_ins_2),
    .io_ins_3(ces_4_4_io_ins_3),
    .io_outs_0(ces_4_4_io_outs_0),
    .io_outs_1(ces_4_4_io_outs_1),
    .io_outs_2(ces_4_4_io_outs_2),
    .io_outs_3(ces_4_4_io_outs_3)
  );
  Element ces_4_5 ( // @[MockArray.scala 36:52]
    .clock(ces_4_5_clock),
    .io_ins_0(ces_4_5_io_ins_0),
    .io_ins_1(ces_4_5_io_ins_1),
    .io_ins_2(ces_4_5_io_ins_2),
    .io_ins_3(ces_4_5_io_ins_3),
    .io_outs_0(ces_4_5_io_outs_0),
    .io_outs_1(ces_4_5_io_outs_1),
    .io_outs_2(ces_4_5_io_outs_2),
    .io_outs_3(ces_4_5_io_outs_3)
  );
  Element ces_4_6 ( // @[MockArray.scala 36:52]
    .clock(ces_4_6_clock),
    .io_ins_0(ces_4_6_io_ins_0),
    .io_ins_1(ces_4_6_io_ins_1),
    .io_ins_2(ces_4_6_io_ins_2),
    .io_ins_3(ces_4_6_io_ins_3),
    .io_outs_0(ces_4_6_io_outs_0),
    .io_outs_1(ces_4_6_io_outs_1),
    .io_outs_2(ces_4_6_io_outs_2),
    .io_outs_3(ces_4_6_io_outs_3)
  );
  Element ces_4_7 ( // @[MockArray.scala 36:52]
    .clock(ces_4_7_clock),
    .io_ins_0(ces_4_7_io_ins_0),
    .io_ins_1(ces_4_7_io_ins_1),
    .io_ins_2(ces_4_7_io_ins_2),
    .io_ins_3(ces_4_7_io_ins_3),
    .io_outs_0(ces_4_7_io_outs_0),
    .io_outs_1(ces_4_7_io_outs_1),
    .io_outs_2(ces_4_7_io_outs_2),
    .io_outs_3(ces_4_7_io_outs_3)
  );
  Element ces_4_8 ( // @[MockArray.scala 36:52]
    .clock(ces_4_8_clock),
    .io_ins_0(ces_4_8_io_ins_0),
    .io_ins_1(ces_4_8_io_ins_1),
    .io_ins_2(ces_4_8_io_ins_2),
    .io_ins_3(ces_4_8_io_ins_3),
    .io_outs_0(ces_4_8_io_outs_0),
    .io_outs_1(ces_4_8_io_outs_1),
    .io_outs_2(ces_4_8_io_outs_2),
    .io_outs_3(ces_4_8_io_outs_3)
  );
  Element ces_4_9 ( // @[MockArray.scala 36:52]
    .clock(ces_4_9_clock),
    .io_ins_0(ces_4_9_io_ins_0),
    .io_ins_1(ces_4_9_io_ins_1),
    .io_ins_2(ces_4_9_io_ins_2),
    .io_ins_3(ces_4_9_io_ins_3),
    .io_outs_0(ces_4_9_io_outs_0),
    .io_outs_1(ces_4_9_io_outs_1),
    .io_outs_2(ces_4_9_io_outs_2),
    .io_outs_3(ces_4_9_io_outs_3)
  );
  Element ces_4_10 ( // @[MockArray.scala 36:52]
    .clock(ces_4_10_clock),
    .io_ins_0(ces_4_10_io_ins_0),
    .io_ins_1(ces_4_10_io_ins_1),
    .io_ins_2(ces_4_10_io_ins_2),
    .io_ins_3(ces_4_10_io_ins_3),
    .io_outs_0(ces_4_10_io_outs_0),
    .io_outs_1(ces_4_10_io_outs_1),
    .io_outs_2(ces_4_10_io_outs_2),
    .io_outs_3(ces_4_10_io_outs_3)
  );
  Element ces_4_11 ( // @[MockArray.scala 36:52]
    .clock(ces_4_11_clock),
    .io_ins_0(ces_4_11_io_ins_0),
    .io_ins_1(ces_4_11_io_ins_1),
    .io_ins_2(ces_4_11_io_ins_2),
    .io_ins_3(ces_4_11_io_ins_3),
    .io_outs_0(ces_4_11_io_outs_0),
    .io_outs_1(ces_4_11_io_outs_1),
    .io_outs_2(ces_4_11_io_outs_2),
    .io_outs_3(ces_4_11_io_outs_3)
  );
  Element ces_4_12 ( // @[MockArray.scala 36:52]
    .clock(ces_4_12_clock),
    .io_ins_0(ces_4_12_io_ins_0),
    .io_ins_1(ces_4_12_io_ins_1),
    .io_ins_2(ces_4_12_io_ins_2),
    .io_ins_3(ces_4_12_io_ins_3),
    .io_outs_0(ces_4_12_io_outs_0),
    .io_outs_1(ces_4_12_io_outs_1),
    .io_outs_2(ces_4_12_io_outs_2),
    .io_outs_3(ces_4_12_io_outs_3)
  );
  Element ces_4_13 ( // @[MockArray.scala 36:52]
    .clock(ces_4_13_clock),
    .io_ins_0(ces_4_13_io_ins_0),
    .io_ins_1(ces_4_13_io_ins_1),
    .io_ins_2(ces_4_13_io_ins_2),
    .io_ins_3(ces_4_13_io_ins_3),
    .io_outs_0(ces_4_13_io_outs_0),
    .io_outs_1(ces_4_13_io_outs_1),
    .io_outs_2(ces_4_13_io_outs_2),
    .io_outs_3(ces_4_13_io_outs_3)
  );
  Element ces_4_14 ( // @[MockArray.scala 36:52]
    .clock(ces_4_14_clock),
    .io_ins_0(ces_4_14_io_ins_0),
    .io_ins_1(ces_4_14_io_ins_1),
    .io_ins_2(ces_4_14_io_ins_2),
    .io_ins_3(ces_4_14_io_ins_3),
    .io_outs_0(ces_4_14_io_outs_0),
    .io_outs_1(ces_4_14_io_outs_1),
    .io_outs_2(ces_4_14_io_outs_2),
    .io_outs_3(ces_4_14_io_outs_3)
  );
  Element ces_4_15 ( // @[MockArray.scala 36:52]
    .clock(ces_4_15_clock),
    .io_ins_0(ces_4_15_io_ins_0),
    .io_ins_1(ces_4_15_io_ins_1),
    .io_ins_2(ces_4_15_io_ins_2),
    .io_ins_3(ces_4_15_io_ins_3),
    .io_outs_0(ces_4_15_io_outs_0),
    .io_outs_1(ces_4_15_io_outs_1),
    .io_outs_2(ces_4_15_io_outs_2),
    .io_outs_3(ces_4_15_io_outs_3)
  );
  Element ces_4_16 ( // @[MockArray.scala 36:52]
    .clock(ces_4_16_clock),
    .io_ins_0(ces_4_16_io_ins_0),
    .io_ins_1(ces_4_16_io_ins_1),
    .io_ins_2(ces_4_16_io_ins_2),
    .io_ins_3(ces_4_16_io_ins_3),
    .io_outs_0(ces_4_16_io_outs_0),
    .io_outs_1(ces_4_16_io_outs_1),
    .io_outs_2(ces_4_16_io_outs_2),
    .io_outs_3(ces_4_16_io_outs_3)
  );
  Element ces_4_17 ( // @[MockArray.scala 36:52]
    .clock(ces_4_17_clock),
    .io_ins_0(ces_4_17_io_ins_0),
    .io_ins_1(ces_4_17_io_ins_1),
    .io_ins_2(ces_4_17_io_ins_2),
    .io_ins_3(ces_4_17_io_ins_3),
    .io_outs_0(ces_4_17_io_outs_0),
    .io_outs_1(ces_4_17_io_outs_1),
    .io_outs_2(ces_4_17_io_outs_2),
    .io_outs_3(ces_4_17_io_outs_3)
  );
  Element ces_4_18 ( // @[MockArray.scala 36:52]
    .clock(ces_4_18_clock),
    .io_ins_0(ces_4_18_io_ins_0),
    .io_ins_1(ces_4_18_io_ins_1),
    .io_ins_2(ces_4_18_io_ins_2),
    .io_ins_3(ces_4_18_io_ins_3),
    .io_outs_0(ces_4_18_io_outs_0),
    .io_outs_1(ces_4_18_io_outs_1),
    .io_outs_2(ces_4_18_io_outs_2),
    .io_outs_3(ces_4_18_io_outs_3)
  );
  Element ces_4_19 ( // @[MockArray.scala 36:52]
    .clock(ces_4_19_clock),
    .io_ins_0(ces_4_19_io_ins_0),
    .io_ins_1(ces_4_19_io_ins_1),
    .io_ins_2(ces_4_19_io_ins_2),
    .io_ins_3(ces_4_19_io_ins_3),
    .io_outs_0(ces_4_19_io_outs_0),
    .io_outs_1(ces_4_19_io_outs_1),
    .io_outs_2(ces_4_19_io_outs_2),
    .io_outs_3(ces_4_19_io_outs_3)
  );
  Element ces_4_20 ( // @[MockArray.scala 36:52]
    .clock(ces_4_20_clock),
    .io_ins_0(ces_4_20_io_ins_0),
    .io_ins_1(ces_4_20_io_ins_1),
    .io_ins_2(ces_4_20_io_ins_2),
    .io_ins_3(ces_4_20_io_ins_3),
    .io_outs_0(ces_4_20_io_outs_0),
    .io_outs_1(ces_4_20_io_outs_1),
    .io_outs_2(ces_4_20_io_outs_2),
    .io_outs_3(ces_4_20_io_outs_3)
  );
  Element ces_4_21 ( // @[MockArray.scala 36:52]
    .clock(ces_4_21_clock),
    .io_ins_0(ces_4_21_io_ins_0),
    .io_ins_1(ces_4_21_io_ins_1),
    .io_ins_2(ces_4_21_io_ins_2),
    .io_ins_3(ces_4_21_io_ins_3),
    .io_outs_0(ces_4_21_io_outs_0),
    .io_outs_1(ces_4_21_io_outs_1),
    .io_outs_2(ces_4_21_io_outs_2),
    .io_outs_3(ces_4_21_io_outs_3)
  );
  Element ces_4_22 ( // @[MockArray.scala 36:52]
    .clock(ces_4_22_clock),
    .io_ins_0(ces_4_22_io_ins_0),
    .io_ins_1(ces_4_22_io_ins_1),
    .io_ins_2(ces_4_22_io_ins_2),
    .io_ins_3(ces_4_22_io_ins_3),
    .io_outs_0(ces_4_22_io_outs_0),
    .io_outs_1(ces_4_22_io_outs_1),
    .io_outs_2(ces_4_22_io_outs_2),
    .io_outs_3(ces_4_22_io_outs_3)
  );
  Element ces_4_23 ( // @[MockArray.scala 36:52]
    .clock(ces_4_23_clock),
    .io_ins_0(ces_4_23_io_ins_0),
    .io_ins_1(ces_4_23_io_ins_1),
    .io_ins_2(ces_4_23_io_ins_2),
    .io_ins_3(ces_4_23_io_ins_3),
    .io_outs_0(ces_4_23_io_outs_0),
    .io_outs_1(ces_4_23_io_outs_1),
    .io_outs_2(ces_4_23_io_outs_2),
    .io_outs_3(ces_4_23_io_outs_3)
  );
  Element ces_4_24 ( // @[MockArray.scala 36:52]
    .clock(ces_4_24_clock),
    .io_ins_0(ces_4_24_io_ins_0),
    .io_ins_1(ces_4_24_io_ins_1),
    .io_ins_2(ces_4_24_io_ins_2),
    .io_ins_3(ces_4_24_io_ins_3),
    .io_outs_0(ces_4_24_io_outs_0),
    .io_outs_1(ces_4_24_io_outs_1),
    .io_outs_2(ces_4_24_io_outs_2),
    .io_outs_3(ces_4_24_io_outs_3)
  );
  Element ces_4_25 ( // @[MockArray.scala 36:52]
    .clock(ces_4_25_clock),
    .io_ins_0(ces_4_25_io_ins_0),
    .io_ins_1(ces_4_25_io_ins_1),
    .io_ins_2(ces_4_25_io_ins_2),
    .io_ins_3(ces_4_25_io_ins_3),
    .io_outs_0(ces_4_25_io_outs_0),
    .io_outs_1(ces_4_25_io_outs_1),
    .io_outs_2(ces_4_25_io_outs_2),
    .io_outs_3(ces_4_25_io_outs_3)
  );
  Element ces_4_26 ( // @[MockArray.scala 36:52]
    .clock(ces_4_26_clock),
    .io_ins_0(ces_4_26_io_ins_0),
    .io_ins_1(ces_4_26_io_ins_1),
    .io_ins_2(ces_4_26_io_ins_2),
    .io_ins_3(ces_4_26_io_ins_3),
    .io_outs_0(ces_4_26_io_outs_0),
    .io_outs_1(ces_4_26_io_outs_1),
    .io_outs_2(ces_4_26_io_outs_2),
    .io_outs_3(ces_4_26_io_outs_3)
  );
  Element ces_4_27 ( // @[MockArray.scala 36:52]
    .clock(ces_4_27_clock),
    .io_ins_0(ces_4_27_io_ins_0),
    .io_ins_1(ces_4_27_io_ins_1),
    .io_ins_2(ces_4_27_io_ins_2),
    .io_ins_3(ces_4_27_io_ins_3),
    .io_outs_0(ces_4_27_io_outs_0),
    .io_outs_1(ces_4_27_io_outs_1),
    .io_outs_2(ces_4_27_io_outs_2),
    .io_outs_3(ces_4_27_io_outs_3)
  );
  Element ces_4_28 ( // @[MockArray.scala 36:52]
    .clock(ces_4_28_clock),
    .io_ins_0(ces_4_28_io_ins_0),
    .io_ins_1(ces_4_28_io_ins_1),
    .io_ins_2(ces_4_28_io_ins_2),
    .io_ins_3(ces_4_28_io_ins_3),
    .io_outs_0(ces_4_28_io_outs_0),
    .io_outs_1(ces_4_28_io_outs_1),
    .io_outs_2(ces_4_28_io_outs_2),
    .io_outs_3(ces_4_28_io_outs_3)
  );
  Element ces_4_29 ( // @[MockArray.scala 36:52]
    .clock(ces_4_29_clock),
    .io_ins_0(ces_4_29_io_ins_0),
    .io_ins_1(ces_4_29_io_ins_1),
    .io_ins_2(ces_4_29_io_ins_2),
    .io_ins_3(ces_4_29_io_ins_3),
    .io_outs_0(ces_4_29_io_outs_0),
    .io_outs_1(ces_4_29_io_outs_1),
    .io_outs_2(ces_4_29_io_outs_2),
    .io_outs_3(ces_4_29_io_outs_3)
  );
  Element ces_4_30 ( // @[MockArray.scala 36:52]
    .clock(ces_4_30_clock),
    .io_ins_0(ces_4_30_io_ins_0),
    .io_ins_1(ces_4_30_io_ins_1),
    .io_ins_2(ces_4_30_io_ins_2),
    .io_ins_3(ces_4_30_io_ins_3),
    .io_outs_0(ces_4_30_io_outs_0),
    .io_outs_1(ces_4_30_io_outs_1),
    .io_outs_2(ces_4_30_io_outs_2),
    .io_outs_3(ces_4_30_io_outs_3)
  );
  Element ces_4_31 ( // @[MockArray.scala 36:52]
    .clock(ces_4_31_clock),
    .io_ins_0(ces_4_31_io_ins_0),
    .io_ins_1(ces_4_31_io_ins_1),
    .io_ins_2(ces_4_31_io_ins_2),
    .io_ins_3(ces_4_31_io_ins_3),
    .io_outs_0(ces_4_31_io_outs_0),
    .io_outs_1(ces_4_31_io_outs_1),
    .io_outs_2(ces_4_31_io_outs_2),
    .io_outs_3(ces_4_31_io_outs_3)
  );
  Element ces_5_0 ( // @[MockArray.scala 36:52]
    .clock(ces_5_0_clock),
    .io_ins_0(ces_5_0_io_ins_0),
    .io_ins_1(ces_5_0_io_ins_1),
    .io_ins_2(ces_5_0_io_ins_2),
    .io_ins_3(ces_5_0_io_ins_3),
    .io_outs_0(ces_5_0_io_outs_0),
    .io_outs_1(ces_5_0_io_outs_1),
    .io_outs_2(ces_5_0_io_outs_2),
    .io_outs_3(ces_5_0_io_outs_3)
  );
  Element ces_5_1 ( // @[MockArray.scala 36:52]
    .clock(ces_5_1_clock),
    .io_ins_0(ces_5_1_io_ins_0),
    .io_ins_1(ces_5_1_io_ins_1),
    .io_ins_2(ces_5_1_io_ins_2),
    .io_ins_3(ces_5_1_io_ins_3),
    .io_outs_0(ces_5_1_io_outs_0),
    .io_outs_1(ces_5_1_io_outs_1),
    .io_outs_2(ces_5_1_io_outs_2),
    .io_outs_3(ces_5_1_io_outs_3)
  );
  Element ces_5_2 ( // @[MockArray.scala 36:52]
    .clock(ces_5_2_clock),
    .io_ins_0(ces_5_2_io_ins_0),
    .io_ins_1(ces_5_2_io_ins_1),
    .io_ins_2(ces_5_2_io_ins_2),
    .io_ins_3(ces_5_2_io_ins_3),
    .io_outs_0(ces_5_2_io_outs_0),
    .io_outs_1(ces_5_2_io_outs_1),
    .io_outs_2(ces_5_2_io_outs_2),
    .io_outs_3(ces_5_2_io_outs_3)
  );
  Element ces_5_3 ( // @[MockArray.scala 36:52]
    .clock(ces_5_3_clock),
    .io_ins_0(ces_5_3_io_ins_0),
    .io_ins_1(ces_5_3_io_ins_1),
    .io_ins_2(ces_5_3_io_ins_2),
    .io_ins_3(ces_5_3_io_ins_3),
    .io_outs_0(ces_5_3_io_outs_0),
    .io_outs_1(ces_5_3_io_outs_1),
    .io_outs_2(ces_5_3_io_outs_2),
    .io_outs_3(ces_5_3_io_outs_3)
  );
  Element ces_5_4 ( // @[MockArray.scala 36:52]
    .clock(ces_5_4_clock),
    .io_ins_0(ces_5_4_io_ins_0),
    .io_ins_1(ces_5_4_io_ins_1),
    .io_ins_2(ces_5_4_io_ins_2),
    .io_ins_3(ces_5_4_io_ins_3),
    .io_outs_0(ces_5_4_io_outs_0),
    .io_outs_1(ces_5_4_io_outs_1),
    .io_outs_2(ces_5_4_io_outs_2),
    .io_outs_3(ces_5_4_io_outs_3)
  );
  Element ces_5_5 ( // @[MockArray.scala 36:52]
    .clock(ces_5_5_clock),
    .io_ins_0(ces_5_5_io_ins_0),
    .io_ins_1(ces_5_5_io_ins_1),
    .io_ins_2(ces_5_5_io_ins_2),
    .io_ins_3(ces_5_5_io_ins_3),
    .io_outs_0(ces_5_5_io_outs_0),
    .io_outs_1(ces_5_5_io_outs_1),
    .io_outs_2(ces_5_5_io_outs_2),
    .io_outs_3(ces_5_5_io_outs_3)
  );
  Element ces_5_6 ( // @[MockArray.scala 36:52]
    .clock(ces_5_6_clock),
    .io_ins_0(ces_5_6_io_ins_0),
    .io_ins_1(ces_5_6_io_ins_1),
    .io_ins_2(ces_5_6_io_ins_2),
    .io_ins_3(ces_5_6_io_ins_3),
    .io_outs_0(ces_5_6_io_outs_0),
    .io_outs_1(ces_5_6_io_outs_1),
    .io_outs_2(ces_5_6_io_outs_2),
    .io_outs_3(ces_5_6_io_outs_3)
  );
  Element ces_5_7 ( // @[MockArray.scala 36:52]
    .clock(ces_5_7_clock),
    .io_ins_0(ces_5_7_io_ins_0),
    .io_ins_1(ces_5_7_io_ins_1),
    .io_ins_2(ces_5_7_io_ins_2),
    .io_ins_3(ces_5_7_io_ins_3),
    .io_outs_0(ces_5_7_io_outs_0),
    .io_outs_1(ces_5_7_io_outs_1),
    .io_outs_2(ces_5_7_io_outs_2),
    .io_outs_3(ces_5_7_io_outs_3)
  );
  Element ces_5_8 ( // @[MockArray.scala 36:52]
    .clock(ces_5_8_clock),
    .io_ins_0(ces_5_8_io_ins_0),
    .io_ins_1(ces_5_8_io_ins_1),
    .io_ins_2(ces_5_8_io_ins_2),
    .io_ins_3(ces_5_8_io_ins_3),
    .io_outs_0(ces_5_8_io_outs_0),
    .io_outs_1(ces_5_8_io_outs_1),
    .io_outs_2(ces_5_8_io_outs_2),
    .io_outs_3(ces_5_8_io_outs_3)
  );
  Element ces_5_9 ( // @[MockArray.scala 36:52]
    .clock(ces_5_9_clock),
    .io_ins_0(ces_5_9_io_ins_0),
    .io_ins_1(ces_5_9_io_ins_1),
    .io_ins_2(ces_5_9_io_ins_2),
    .io_ins_3(ces_5_9_io_ins_3),
    .io_outs_0(ces_5_9_io_outs_0),
    .io_outs_1(ces_5_9_io_outs_1),
    .io_outs_2(ces_5_9_io_outs_2),
    .io_outs_3(ces_5_9_io_outs_3)
  );
  Element ces_5_10 ( // @[MockArray.scala 36:52]
    .clock(ces_5_10_clock),
    .io_ins_0(ces_5_10_io_ins_0),
    .io_ins_1(ces_5_10_io_ins_1),
    .io_ins_2(ces_5_10_io_ins_2),
    .io_ins_3(ces_5_10_io_ins_3),
    .io_outs_0(ces_5_10_io_outs_0),
    .io_outs_1(ces_5_10_io_outs_1),
    .io_outs_2(ces_5_10_io_outs_2),
    .io_outs_3(ces_5_10_io_outs_3)
  );
  Element ces_5_11 ( // @[MockArray.scala 36:52]
    .clock(ces_5_11_clock),
    .io_ins_0(ces_5_11_io_ins_0),
    .io_ins_1(ces_5_11_io_ins_1),
    .io_ins_2(ces_5_11_io_ins_2),
    .io_ins_3(ces_5_11_io_ins_3),
    .io_outs_0(ces_5_11_io_outs_0),
    .io_outs_1(ces_5_11_io_outs_1),
    .io_outs_2(ces_5_11_io_outs_2),
    .io_outs_3(ces_5_11_io_outs_3)
  );
  Element ces_5_12 ( // @[MockArray.scala 36:52]
    .clock(ces_5_12_clock),
    .io_ins_0(ces_5_12_io_ins_0),
    .io_ins_1(ces_5_12_io_ins_1),
    .io_ins_2(ces_5_12_io_ins_2),
    .io_ins_3(ces_5_12_io_ins_3),
    .io_outs_0(ces_5_12_io_outs_0),
    .io_outs_1(ces_5_12_io_outs_1),
    .io_outs_2(ces_5_12_io_outs_2),
    .io_outs_3(ces_5_12_io_outs_3)
  );
  Element ces_5_13 ( // @[MockArray.scala 36:52]
    .clock(ces_5_13_clock),
    .io_ins_0(ces_5_13_io_ins_0),
    .io_ins_1(ces_5_13_io_ins_1),
    .io_ins_2(ces_5_13_io_ins_2),
    .io_ins_3(ces_5_13_io_ins_3),
    .io_outs_0(ces_5_13_io_outs_0),
    .io_outs_1(ces_5_13_io_outs_1),
    .io_outs_2(ces_5_13_io_outs_2),
    .io_outs_3(ces_5_13_io_outs_3)
  );
  Element ces_5_14 ( // @[MockArray.scala 36:52]
    .clock(ces_5_14_clock),
    .io_ins_0(ces_5_14_io_ins_0),
    .io_ins_1(ces_5_14_io_ins_1),
    .io_ins_2(ces_5_14_io_ins_2),
    .io_ins_3(ces_5_14_io_ins_3),
    .io_outs_0(ces_5_14_io_outs_0),
    .io_outs_1(ces_5_14_io_outs_1),
    .io_outs_2(ces_5_14_io_outs_2),
    .io_outs_3(ces_5_14_io_outs_3)
  );
  Element ces_5_15 ( // @[MockArray.scala 36:52]
    .clock(ces_5_15_clock),
    .io_ins_0(ces_5_15_io_ins_0),
    .io_ins_1(ces_5_15_io_ins_1),
    .io_ins_2(ces_5_15_io_ins_2),
    .io_ins_3(ces_5_15_io_ins_3),
    .io_outs_0(ces_5_15_io_outs_0),
    .io_outs_1(ces_5_15_io_outs_1),
    .io_outs_2(ces_5_15_io_outs_2),
    .io_outs_3(ces_5_15_io_outs_3)
  );
  Element ces_5_16 ( // @[MockArray.scala 36:52]
    .clock(ces_5_16_clock),
    .io_ins_0(ces_5_16_io_ins_0),
    .io_ins_1(ces_5_16_io_ins_1),
    .io_ins_2(ces_5_16_io_ins_2),
    .io_ins_3(ces_5_16_io_ins_3),
    .io_outs_0(ces_5_16_io_outs_0),
    .io_outs_1(ces_5_16_io_outs_1),
    .io_outs_2(ces_5_16_io_outs_2),
    .io_outs_3(ces_5_16_io_outs_3)
  );
  Element ces_5_17 ( // @[MockArray.scala 36:52]
    .clock(ces_5_17_clock),
    .io_ins_0(ces_5_17_io_ins_0),
    .io_ins_1(ces_5_17_io_ins_1),
    .io_ins_2(ces_5_17_io_ins_2),
    .io_ins_3(ces_5_17_io_ins_3),
    .io_outs_0(ces_5_17_io_outs_0),
    .io_outs_1(ces_5_17_io_outs_1),
    .io_outs_2(ces_5_17_io_outs_2),
    .io_outs_3(ces_5_17_io_outs_3)
  );
  Element ces_5_18 ( // @[MockArray.scala 36:52]
    .clock(ces_5_18_clock),
    .io_ins_0(ces_5_18_io_ins_0),
    .io_ins_1(ces_5_18_io_ins_1),
    .io_ins_2(ces_5_18_io_ins_2),
    .io_ins_3(ces_5_18_io_ins_3),
    .io_outs_0(ces_5_18_io_outs_0),
    .io_outs_1(ces_5_18_io_outs_1),
    .io_outs_2(ces_5_18_io_outs_2),
    .io_outs_3(ces_5_18_io_outs_3)
  );
  Element ces_5_19 ( // @[MockArray.scala 36:52]
    .clock(ces_5_19_clock),
    .io_ins_0(ces_5_19_io_ins_0),
    .io_ins_1(ces_5_19_io_ins_1),
    .io_ins_2(ces_5_19_io_ins_2),
    .io_ins_3(ces_5_19_io_ins_3),
    .io_outs_0(ces_5_19_io_outs_0),
    .io_outs_1(ces_5_19_io_outs_1),
    .io_outs_2(ces_5_19_io_outs_2),
    .io_outs_3(ces_5_19_io_outs_3)
  );
  Element ces_5_20 ( // @[MockArray.scala 36:52]
    .clock(ces_5_20_clock),
    .io_ins_0(ces_5_20_io_ins_0),
    .io_ins_1(ces_5_20_io_ins_1),
    .io_ins_2(ces_5_20_io_ins_2),
    .io_ins_3(ces_5_20_io_ins_3),
    .io_outs_0(ces_5_20_io_outs_0),
    .io_outs_1(ces_5_20_io_outs_1),
    .io_outs_2(ces_5_20_io_outs_2),
    .io_outs_3(ces_5_20_io_outs_3)
  );
  Element ces_5_21 ( // @[MockArray.scala 36:52]
    .clock(ces_5_21_clock),
    .io_ins_0(ces_5_21_io_ins_0),
    .io_ins_1(ces_5_21_io_ins_1),
    .io_ins_2(ces_5_21_io_ins_2),
    .io_ins_3(ces_5_21_io_ins_3),
    .io_outs_0(ces_5_21_io_outs_0),
    .io_outs_1(ces_5_21_io_outs_1),
    .io_outs_2(ces_5_21_io_outs_2),
    .io_outs_3(ces_5_21_io_outs_3)
  );
  Element ces_5_22 ( // @[MockArray.scala 36:52]
    .clock(ces_5_22_clock),
    .io_ins_0(ces_5_22_io_ins_0),
    .io_ins_1(ces_5_22_io_ins_1),
    .io_ins_2(ces_5_22_io_ins_2),
    .io_ins_3(ces_5_22_io_ins_3),
    .io_outs_0(ces_5_22_io_outs_0),
    .io_outs_1(ces_5_22_io_outs_1),
    .io_outs_2(ces_5_22_io_outs_2),
    .io_outs_3(ces_5_22_io_outs_3)
  );
  Element ces_5_23 ( // @[MockArray.scala 36:52]
    .clock(ces_5_23_clock),
    .io_ins_0(ces_5_23_io_ins_0),
    .io_ins_1(ces_5_23_io_ins_1),
    .io_ins_2(ces_5_23_io_ins_2),
    .io_ins_3(ces_5_23_io_ins_3),
    .io_outs_0(ces_5_23_io_outs_0),
    .io_outs_1(ces_5_23_io_outs_1),
    .io_outs_2(ces_5_23_io_outs_2),
    .io_outs_3(ces_5_23_io_outs_3)
  );
  Element ces_5_24 ( // @[MockArray.scala 36:52]
    .clock(ces_5_24_clock),
    .io_ins_0(ces_5_24_io_ins_0),
    .io_ins_1(ces_5_24_io_ins_1),
    .io_ins_2(ces_5_24_io_ins_2),
    .io_ins_3(ces_5_24_io_ins_3),
    .io_outs_0(ces_5_24_io_outs_0),
    .io_outs_1(ces_5_24_io_outs_1),
    .io_outs_2(ces_5_24_io_outs_2),
    .io_outs_3(ces_5_24_io_outs_3)
  );
  Element ces_5_25 ( // @[MockArray.scala 36:52]
    .clock(ces_5_25_clock),
    .io_ins_0(ces_5_25_io_ins_0),
    .io_ins_1(ces_5_25_io_ins_1),
    .io_ins_2(ces_5_25_io_ins_2),
    .io_ins_3(ces_5_25_io_ins_3),
    .io_outs_0(ces_5_25_io_outs_0),
    .io_outs_1(ces_5_25_io_outs_1),
    .io_outs_2(ces_5_25_io_outs_2),
    .io_outs_3(ces_5_25_io_outs_3)
  );
  Element ces_5_26 ( // @[MockArray.scala 36:52]
    .clock(ces_5_26_clock),
    .io_ins_0(ces_5_26_io_ins_0),
    .io_ins_1(ces_5_26_io_ins_1),
    .io_ins_2(ces_5_26_io_ins_2),
    .io_ins_3(ces_5_26_io_ins_3),
    .io_outs_0(ces_5_26_io_outs_0),
    .io_outs_1(ces_5_26_io_outs_1),
    .io_outs_2(ces_5_26_io_outs_2),
    .io_outs_3(ces_5_26_io_outs_3)
  );
  Element ces_5_27 ( // @[MockArray.scala 36:52]
    .clock(ces_5_27_clock),
    .io_ins_0(ces_5_27_io_ins_0),
    .io_ins_1(ces_5_27_io_ins_1),
    .io_ins_2(ces_5_27_io_ins_2),
    .io_ins_3(ces_5_27_io_ins_3),
    .io_outs_0(ces_5_27_io_outs_0),
    .io_outs_1(ces_5_27_io_outs_1),
    .io_outs_2(ces_5_27_io_outs_2),
    .io_outs_3(ces_5_27_io_outs_3)
  );
  Element ces_5_28 ( // @[MockArray.scala 36:52]
    .clock(ces_5_28_clock),
    .io_ins_0(ces_5_28_io_ins_0),
    .io_ins_1(ces_5_28_io_ins_1),
    .io_ins_2(ces_5_28_io_ins_2),
    .io_ins_3(ces_5_28_io_ins_3),
    .io_outs_0(ces_5_28_io_outs_0),
    .io_outs_1(ces_5_28_io_outs_1),
    .io_outs_2(ces_5_28_io_outs_2),
    .io_outs_3(ces_5_28_io_outs_3)
  );
  Element ces_5_29 ( // @[MockArray.scala 36:52]
    .clock(ces_5_29_clock),
    .io_ins_0(ces_5_29_io_ins_0),
    .io_ins_1(ces_5_29_io_ins_1),
    .io_ins_2(ces_5_29_io_ins_2),
    .io_ins_3(ces_5_29_io_ins_3),
    .io_outs_0(ces_5_29_io_outs_0),
    .io_outs_1(ces_5_29_io_outs_1),
    .io_outs_2(ces_5_29_io_outs_2),
    .io_outs_3(ces_5_29_io_outs_3)
  );
  Element ces_5_30 ( // @[MockArray.scala 36:52]
    .clock(ces_5_30_clock),
    .io_ins_0(ces_5_30_io_ins_0),
    .io_ins_1(ces_5_30_io_ins_1),
    .io_ins_2(ces_5_30_io_ins_2),
    .io_ins_3(ces_5_30_io_ins_3),
    .io_outs_0(ces_5_30_io_outs_0),
    .io_outs_1(ces_5_30_io_outs_1),
    .io_outs_2(ces_5_30_io_outs_2),
    .io_outs_3(ces_5_30_io_outs_3)
  );
  Element ces_5_31 ( // @[MockArray.scala 36:52]
    .clock(ces_5_31_clock),
    .io_ins_0(ces_5_31_io_ins_0),
    .io_ins_1(ces_5_31_io_ins_1),
    .io_ins_2(ces_5_31_io_ins_2),
    .io_ins_3(ces_5_31_io_ins_3),
    .io_outs_0(ces_5_31_io_outs_0),
    .io_outs_1(ces_5_31_io_outs_1),
    .io_outs_2(ces_5_31_io_outs_2),
    .io_outs_3(ces_5_31_io_outs_3)
  );
  Element ces_6_0 ( // @[MockArray.scala 36:52]
    .clock(ces_6_0_clock),
    .io_ins_0(ces_6_0_io_ins_0),
    .io_ins_1(ces_6_0_io_ins_1),
    .io_ins_2(ces_6_0_io_ins_2),
    .io_ins_3(ces_6_0_io_ins_3),
    .io_outs_0(ces_6_0_io_outs_0),
    .io_outs_1(ces_6_0_io_outs_1),
    .io_outs_2(ces_6_0_io_outs_2),
    .io_outs_3(ces_6_0_io_outs_3)
  );
  Element ces_6_1 ( // @[MockArray.scala 36:52]
    .clock(ces_6_1_clock),
    .io_ins_0(ces_6_1_io_ins_0),
    .io_ins_1(ces_6_1_io_ins_1),
    .io_ins_2(ces_6_1_io_ins_2),
    .io_ins_3(ces_6_1_io_ins_3),
    .io_outs_0(ces_6_1_io_outs_0),
    .io_outs_1(ces_6_1_io_outs_1),
    .io_outs_2(ces_6_1_io_outs_2),
    .io_outs_3(ces_6_1_io_outs_3)
  );
  Element ces_6_2 ( // @[MockArray.scala 36:52]
    .clock(ces_6_2_clock),
    .io_ins_0(ces_6_2_io_ins_0),
    .io_ins_1(ces_6_2_io_ins_1),
    .io_ins_2(ces_6_2_io_ins_2),
    .io_ins_3(ces_6_2_io_ins_3),
    .io_outs_0(ces_6_2_io_outs_0),
    .io_outs_1(ces_6_2_io_outs_1),
    .io_outs_2(ces_6_2_io_outs_2),
    .io_outs_3(ces_6_2_io_outs_3)
  );
  Element ces_6_3 ( // @[MockArray.scala 36:52]
    .clock(ces_6_3_clock),
    .io_ins_0(ces_6_3_io_ins_0),
    .io_ins_1(ces_6_3_io_ins_1),
    .io_ins_2(ces_6_3_io_ins_2),
    .io_ins_3(ces_6_3_io_ins_3),
    .io_outs_0(ces_6_3_io_outs_0),
    .io_outs_1(ces_6_3_io_outs_1),
    .io_outs_2(ces_6_3_io_outs_2),
    .io_outs_3(ces_6_3_io_outs_3)
  );
  Element ces_6_4 ( // @[MockArray.scala 36:52]
    .clock(ces_6_4_clock),
    .io_ins_0(ces_6_4_io_ins_0),
    .io_ins_1(ces_6_4_io_ins_1),
    .io_ins_2(ces_6_4_io_ins_2),
    .io_ins_3(ces_6_4_io_ins_3),
    .io_outs_0(ces_6_4_io_outs_0),
    .io_outs_1(ces_6_4_io_outs_1),
    .io_outs_2(ces_6_4_io_outs_2),
    .io_outs_3(ces_6_4_io_outs_3)
  );
  Element ces_6_5 ( // @[MockArray.scala 36:52]
    .clock(ces_6_5_clock),
    .io_ins_0(ces_6_5_io_ins_0),
    .io_ins_1(ces_6_5_io_ins_1),
    .io_ins_2(ces_6_5_io_ins_2),
    .io_ins_3(ces_6_5_io_ins_3),
    .io_outs_0(ces_6_5_io_outs_0),
    .io_outs_1(ces_6_5_io_outs_1),
    .io_outs_2(ces_6_5_io_outs_2),
    .io_outs_3(ces_6_5_io_outs_3)
  );
  Element ces_6_6 ( // @[MockArray.scala 36:52]
    .clock(ces_6_6_clock),
    .io_ins_0(ces_6_6_io_ins_0),
    .io_ins_1(ces_6_6_io_ins_1),
    .io_ins_2(ces_6_6_io_ins_2),
    .io_ins_3(ces_6_6_io_ins_3),
    .io_outs_0(ces_6_6_io_outs_0),
    .io_outs_1(ces_6_6_io_outs_1),
    .io_outs_2(ces_6_6_io_outs_2),
    .io_outs_3(ces_6_6_io_outs_3)
  );
  Element ces_6_7 ( // @[MockArray.scala 36:52]
    .clock(ces_6_7_clock),
    .io_ins_0(ces_6_7_io_ins_0),
    .io_ins_1(ces_6_7_io_ins_1),
    .io_ins_2(ces_6_7_io_ins_2),
    .io_ins_3(ces_6_7_io_ins_3),
    .io_outs_0(ces_6_7_io_outs_0),
    .io_outs_1(ces_6_7_io_outs_1),
    .io_outs_2(ces_6_7_io_outs_2),
    .io_outs_3(ces_6_7_io_outs_3)
  );
  Element ces_6_8 ( // @[MockArray.scala 36:52]
    .clock(ces_6_8_clock),
    .io_ins_0(ces_6_8_io_ins_0),
    .io_ins_1(ces_6_8_io_ins_1),
    .io_ins_2(ces_6_8_io_ins_2),
    .io_ins_3(ces_6_8_io_ins_3),
    .io_outs_0(ces_6_8_io_outs_0),
    .io_outs_1(ces_6_8_io_outs_1),
    .io_outs_2(ces_6_8_io_outs_2),
    .io_outs_3(ces_6_8_io_outs_3)
  );
  Element ces_6_9 ( // @[MockArray.scala 36:52]
    .clock(ces_6_9_clock),
    .io_ins_0(ces_6_9_io_ins_0),
    .io_ins_1(ces_6_9_io_ins_1),
    .io_ins_2(ces_6_9_io_ins_2),
    .io_ins_3(ces_6_9_io_ins_3),
    .io_outs_0(ces_6_9_io_outs_0),
    .io_outs_1(ces_6_9_io_outs_1),
    .io_outs_2(ces_6_9_io_outs_2),
    .io_outs_3(ces_6_9_io_outs_3)
  );
  Element ces_6_10 ( // @[MockArray.scala 36:52]
    .clock(ces_6_10_clock),
    .io_ins_0(ces_6_10_io_ins_0),
    .io_ins_1(ces_6_10_io_ins_1),
    .io_ins_2(ces_6_10_io_ins_2),
    .io_ins_3(ces_6_10_io_ins_3),
    .io_outs_0(ces_6_10_io_outs_0),
    .io_outs_1(ces_6_10_io_outs_1),
    .io_outs_2(ces_6_10_io_outs_2),
    .io_outs_3(ces_6_10_io_outs_3)
  );
  Element ces_6_11 ( // @[MockArray.scala 36:52]
    .clock(ces_6_11_clock),
    .io_ins_0(ces_6_11_io_ins_0),
    .io_ins_1(ces_6_11_io_ins_1),
    .io_ins_2(ces_6_11_io_ins_2),
    .io_ins_3(ces_6_11_io_ins_3),
    .io_outs_0(ces_6_11_io_outs_0),
    .io_outs_1(ces_6_11_io_outs_1),
    .io_outs_2(ces_6_11_io_outs_2),
    .io_outs_3(ces_6_11_io_outs_3)
  );
  Element ces_6_12 ( // @[MockArray.scala 36:52]
    .clock(ces_6_12_clock),
    .io_ins_0(ces_6_12_io_ins_0),
    .io_ins_1(ces_6_12_io_ins_1),
    .io_ins_2(ces_6_12_io_ins_2),
    .io_ins_3(ces_6_12_io_ins_3),
    .io_outs_0(ces_6_12_io_outs_0),
    .io_outs_1(ces_6_12_io_outs_1),
    .io_outs_2(ces_6_12_io_outs_2),
    .io_outs_3(ces_6_12_io_outs_3)
  );
  Element ces_6_13 ( // @[MockArray.scala 36:52]
    .clock(ces_6_13_clock),
    .io_ins_0(ces_6_13_io_ins_0),
    .io_ins_1(ces_6_13_io_ins_1),
    .io_ins_2(ces_6_13_io_ins_2),
    .io_ins_3(ces_6_13_io_ins_3),
    .io_outs_0(ces_6_13_io_outs_0),
    .io_outs_1(ces_6_13_io_outs_1),
    .io_outs_2(ces_6_13_io_outs_2),
    .io_outs_3(ces_6_13_io_outs_3)
  );
  Element ces_6_14 ( // @[MockArray.scala 36:52]
    .clock(ces_6_14_clock),
    .io_ins_0(ces_6_14_io_ins_0),
    .io_ins_1(ces_6_14_io_ins_1),
    .io_ins_2(ces_6_14_io_ins_2),
    .io_ins_3(ces_6_14_io_ins_3),
    .io_outs_0(ces_6_14_io_outs_0),
    .io_outs_1(ces_6_14_io_outs_1),
    .io_outs_2(ces_6_14_io_outs_2),
    .io_outs_3(ces_6_14_io_outs_3)
  );
  Element ces_6_15 ( // @[MockArray.scala 36:52]
    .clock(ces_6_15_clock),
    .io_ins_0(ces_6_15_io_ins_0),
    .io_ins_1(ces_6_15_io_ins_1),
    .io_ins_2(ces_6_15_io_ins_2),
    .io_ins_3(ces_6_15_io_ins_3),
    .io_outs_0(ces_6_15_io_outs_0),
    .io_outs_1(ces_6_15_io_outs_1),
    .io_outs_2(ces_6_15_io_outs_2),
    .io_outs_3(ces_6_15_io_outs_3)
  );
  Element ces_6_16 ( // @[MockArray.scala 36:52]
    .clock(ces_6_16_clock),
    .io_ins_0(ces_6_16_io_ins_0),
    .io_ins_1(ces_6_16_io_ins_1),
    .io_ins_2(ces_6_16_io_ins_2),
    .io_ins_3(ces_6_16_io_ins_3),
    .io_outs_0(ces_6_16_io_outs_0),
    .io_outs_1(ces_6_16_io_outs_1),
    .io_outs_2(ces_6_16_io_outs_2),
    .io_outs_3(ces_6_16_io_outs_3)
  );
  Element ces_6_17 ( // @[MockArray.scala 36:52]
    .clock(ces_6_17_clock),
    .io_ins_0(ces_6_17_io_ins_0),
    .io_ins_1(ces_6_17_io_ins_1),
    .io_ins_2(ces_6_17_io_ins_2),
    .io_ins_3(ces_6_17_io_ins_3),
    .io_outs_0(ces_6_17_io_outs_0),
    .io_outs_1(ces_6_17_io_outs_1),
    .io_outs_2(ces_6_17_io_outs_2),
    .io_outs_3(ces_6_17_io_outs_3)
  );
  Element ces_6_18 ( // @[MockArray.scala 36:52]
    .clock(ces_6_18_clock),
    .io_ins_0(ces_6_18_io_ins_0),
    .io_ins_1(ces_6_18_io_ins_1),
    .io_ins_2(ces_6_18_io_ins_2),
    .io_ins_3(ces_6_18_io_ins_3),
    .io_outs_0(ces_6_18_io_outs_0),
    .io_outs_1(ces_6_18_io_outs_1),
    .io_outs_2(ces_6_18_io_outs_2),
    .io_outs_3(ces_6_18_io_outs_3)
  );
  Element ces_6_19 ( // @[MockArray.scala 36:52]
    .clock(ces_6_19_clock),
    .io_ins_0(ces_6_19_io_ins_0),
    .io_ins_1(ces_6_19_io_ins_1),
    .io_ins_2(ces_6_19_io_ins_2),
    .io_ins_3(ces_6_19_io_ins_3),
    .io_outs_0(ces_6_19_io_outs_0),
    .io_outs_1(ces_6_19_io_outs_1),
    .io_outs_2(ces_6_19_io_outs_2),
    .io_outs_3(ces_6_19_io_outs_3)
  );
  Element ces_6_20 ( // @[MockArray.scala 36:52]
    .clock(ces_6_20_clock),
    .io_ins_0(ces_6_20_io_ins_0),
    .io_ins_1(ces_6_20_io_ins_1),
    .io_ins_2(ces_6_20_io_ins_2),
    .io_ins_3(ces_6_20_io_ins_3),
    .io_outs_0(ces_6_20_io_outs_0),
    .io_outs_1(ces_6_20_io_outs_1),
    .io_outs_2(ces_6_20_io_outs_2),
    .io_outs_3(ces_6_20_io_outs_3)
  );
  Element ces_6_21 ( // @[MockArray.scala 36:52]
    .clock(ces_6_21_clock),
    .io_ins_0(ces_6_21_io_ins_0),
    .io_ins_1(ces_6_21_io_ins_1),
    .io_ins_2(ces_6_21_io_ins_2),
    .io_ins_3(ces_6_21_io_ins_3),
    .io_outs_0(ces_6_21_io_outs_0),
    .io_outs_1(ces_6_21_io_outs_1),
    .io_outs_2(ces_6_21_io_outs_2),
    .io_outs_3(ces_6_21_io_outs_3)
  );
  Element ces_6_22 ( // @[MockArray.scala 36:52]
    .clock(ces_6_22_clock),
    .io_ins_0(ces_6_22_io_ins_0),
    .io_ins_1(ces_6_22_io_ins_1),
    .io_ins_2(ces_6_22_io_ins_2),
    .io_ins_3(ces_6_22_io_ins_3),
    .io_outs_0(ces_6_22_io_outs_0),
    .io_outs_1(ces_6_22_io_outs_1),
    .io_outs_2(ces_6_22_io_outs_2),
    .io_outs_3(ces_6_22_io_outs_3)
  );
  Element ces_6_23 ( // @[MockArray.scala 36:52]
    .clock(ces_6_23_clock),
    .io_ins_0(ces_6_23_io_ins_0),
    .io_ins_1(ces_6_23_io_ins_1),
    .io_ins_2(ces_6_23_io_ins_2),
    .io_ins_3(ces_6_23_io_ins_3),
    .io_outs_0(ces_6_23_io_outs_0),
    .io_outs_1(ces_6_23_io_outs_1),
    .io_outs_2(ces_6_23_io_outs_2),
    .io_outs_3(ces_6_23_io_outs_3)
  );
  Element ces_6_24 ( // @[MockArray.scala 36:52]
    .clock(ces_6_24_clock),
    .io_ins_0(ces_6_24_io_ins_0),
    .io_ins_1(ces_6_24_io_ins_1),
    .io_ins_2(ces_6_24_io_ins_2),
    .io_ins_3(ces_6_24_io_ins_3),
    .io_outs_0(ces_6_24_io_outs_0),
    .io_outs_1(ces_6_24_io_outs_1),
    .io_outs_2(ces_6_24_io_outs_2),
    .io_outs_3(ces_6_24_io_outs_3)
  );
  Element ces_6_25 ( // @[MockArray.scala 36:52]
    .clock(ces_6_25_clock),
    .io_ins_0(ces_6_25_io_ins_0),
    .io_ins_1(ces_6_25_io_ins_1),
    .io_ins_2(ces_6_25_io_ins_2),
    .io_ins_3(ces_6_25_io_ins_3),
    .io_outs_0(ces_6_25_io_outs_0),
    .io_outs_1(ces_6_25_io_outs_1),
    .io_outs_2(ces_6_25_io_outs_2),
    .io_outs_3(ces_6_25_io_outs_3)
  );
  Element ces_6_26 ( // @[MockArray.scala 36:52]
    .clock(ces_6_26_clock),
    .io_ins_0(ces_6_26_io_ins_0),
    .io_ins_1(ces_6_26_io_ins_1),
    .io_ins_2(ces_6_26_io_ins_2),
    .io_ins_3(ces_6_26_io_ins_3),
    .io_outs_0(ces_6_26_io_outs_0),
    .io_outs_1(ces_6_26_io_outs_1),
    .io_outs_2(ces_6_26_io_outs_2),
    .io_outs_3(ces_6_26_io_outs_3)
  );
  Element ces_6_27 ( // @[MockArray.scala 36:52]
    .clock(ces_6_27_clock),
    .io_ins_0(ces_6_27_io_ins_0),
    .io_ins_1(ces_6_27_io_ins_1),
    .io_ins_2(ces_6_27_io_ins_2),
    .io_ins_3(ces_6_27_io_ins_3),
    .io_outs_0(ces_6_27_io_outs_0),
    .io_outs_1(ces_6_27_io_outs_1),
    .io_outs_2(ces_6_27_io_outs_2),
    .io_outs_3(ces_6_27_io_outs_3)
  );
  Element ces_6_28 ( // @[MockArray.scala 36:52]
    .clock(ces_6_28_clock),
    .io_ins_0(ces_6_28_io_ins_0),
    .io_ins_1(ces_6_28_io_ins_1),
    .io_ins_2(ces_6_28_io_ins_2),
    .io_ins_3(ces_6_28_io_ins_3),
    .io_outs_0(ces_6_28_io_outs_0),
    .io_outs_1(ces_6_28_io_outs_1),
    .io_outs_2(ces_6_28_io_outs_2),
    .io_outs_3(ces_6_28_io_outs_3)
  );
  Element ces_6_29 ( // @[MockArray.scala 36:52]
    .clock(ces_6_29_clock),
    .io_ins_0(ces_6_29_io_ins_0),
    .io_ins_1(ces_6_29_io_ins_1),
    .io_ins_2(ces_6_29_io_ins_2),
    .io_ins_3(ces_6_29_io_ins_3),
    .io_outs_0(ces_6_29_io_outs_0),
    .io_outs_1(ces_6_29_io_outs_1),
    .io_outs_2(ces_6_29_io_outs_2),
    .io_outs_3(ces_6_29_io_outs_3)
  );
  Element ces_6_30 ( // @[MockArray.scala 36:52]
    .clock(ces_6_30_clock),
    .io_ins_0(ces_6_30_io_ins_0),
    .io_ins_1(ces_6_30_io_ins_1),
    .io_ins_2(ces_6_30_io_ins_2),
    .io_ins_3(ces_6_30_io_ins_3),
    .io_outs_0(ces_6_30_io_outs_0),
    .io_outs_1(ces_6_30_io_outs_1),
    .io_outs_2(ces_6_30_io_outs_2),
    .io_outs_3(ces_6_30_io_outs_3)
  );
  Element ces_6_31 ( // @[MockArray.scala 36:52]
    .clock(ces_6_31_clock),
    .io_ins_0(ces_6_31_io_ins_0),
    .io_ins_1(ces_6_31_io_ins_1),
    .io_ins_2(ces_6_31_io_ins_2),
    .io_ins_3(ces_6_31_io_ins_3),
    .io_outs_0(ces_6_31_io_outs_0),
    .io_outs_1(ces_6_31_io_outs_1),
    .io_outs_2(ces_6_31_io_outs_2),
    .io_outs_3(ces_6_31_io_outs_3)
  );
  Element ces_7_0 ( // @[MockArray.scala 36:52]
    .clock(ces_7_0_clock),
    .io_ins_0(ces_7_0_io_ins_0),
    .io_ins_1(ces_7_0_io_ins_1),
    .io_ins_2(ces_7_0_io_ins_2),
    .io_ins_3(ces_7_0_io_ins_3),
    .io_outs_0(ces_7_0_io_outs_0),
    .io_outs_1(ces_7_0_io_outs_1),
    .io_outs_2(ces_7_0_io_outs_2),
    .io_outs_3(ces_7_0_io_outs_3)
  );
  Element ces_7_1 ( // @[MockArray.scala 36:52]
    .clock(ces_7_1_clock),
    .io_ins_0(ces_7_1_io_ins_0),
    .io_ins_1(ces_7_1_io_ins_1),
    .io_ins_2(ces_7_1_io_ins_2),
    .io_ins_3(ces_7_1_io_ins_3),
    .io_outs_0(ces_7_1_io_outs_0),
    .io_outs_1(ces_7_1_io_outs_1),
    .io_outs_2(ces_7_1_io_outs_2),
    .io_outs_3(ces_7_1_io_outs_3)
  );
  Element ces_7_2 ( // @[MockArray.scala 36:52]
    .clock(ces_7_2_clock),
    .io_ins_0(ces_7_2_io_ins_0),
    .io_ins_1(ces_7_2_io_ins_1),
    .io_ins_2(ces_7_2_io_ins_2),
    .io_ins_3(ces_7_2_io_ins_3),
    .io_outs_0(ces_7_2_io_outs_0),
    .io_outs_1(ces_7_2_io_outs_1),
    .io_outs_2(ces_7_2_io_outs_2),
    .io_outs_3(ces_7_2_io_outs_3)
  );
  Element ces_7_3 ( // @[MockArray.scala 36:52]
    .clock(ces_7_3_clock),
    .io_ins_0(ces_7_3_io_ins_0),
    .io_ins_1(ces_7_3_io_ins_1),
    .io_ins_2(ces_7_3_io_ins_2),
    .io_ins_3(ces_7_3_io_ins_3),
    .io_outs_0(ces_7_3_io_outs_0),
    .io_outs_1(ces_7_3_io_outs_1),
    .io_outs_2(ces_7_3_io_outs_2),
    .io_outs_3(ces_7_3_io_outs_3)
  );
  Element ces_7_4 ( // @[MockArray.scala 36:52]
    .clock(ces_7_4_clock),
    .io_ins_0(ces_7_4_io_ins_0),
    .io_ins_1(ces_7_4_io_ins_1),
    .io_ins_2(ces_7_4_io_ins_2),
    .io_ins_3(ces_7_4_io_ins_3),
    .io_outs_0(ces_7_4_io_outs_0),
    .io_outs_1(ces_7_4_io_outs_1),
    .io_outs_2(ces_7_4_io_outs_2),
    .io_outs_3(ces_7_4_io_outs_3)
  );
  Element ces_7_5 ( // @[MockArray.scala 36:52]
    .clock(ces_7_5_clock),
    .io_ins_0(ces_7_5_io_ins_0),
    .io_ins_1(ces_7_5_io_ins_1),
    .io_ins_2(ces_7_5_io_ins_2),
    .io_ins_3(ces_7_5_io_ins_3),
    .io_outs_0(ces_7_5_io_outs_0),
    .io_outs_1(ces_7_5_io_outs_1),
    .io_outs_2(ces_7_5_io_outs_2),
    .io_outs_3(ces_7_5_io_outs_3)
  );
  Element ces_7_6 ( // @[MockArray.scala 36:52]
    .clock(ces_7_6_clock),
    .io_ins_0(ces_7_6_io_ins_0),
    .io_ins_1(ces_7_6_io_ins_1),
    .io_ins_2(ces_7_6_io_ins_2),
    .io_ins_3(ces_7_6_io_ins_3),
    .io_outs_0(ces_7_6_io_outs_0),
    .io_outs_1(ces_7_6_io_outs_1),
    .io_outs_2(ces_7_6_io_outs_2),
    .io_outs_3(ces_7_6_io_outs_3)
  );
  Element ces_7_7 ( // @[MockArray.scala 36:52]
    .clock(ces_7_7_clock),
    .io_ins_0(ces_7_7_io_ins_0),
    .io_ins_1(ces_7_7_io_ins_1),
    .io_ins_2(ces_7_7_io_ins_2),
    .io_ins_3(ces_7_7_io_ins_3),
    .io_outs_0(ces_7_7_io_outs_0),
    .io_outs_1(ces_7_7_io_outs_1),
    .io_outs_2(ces_7_7_io_outs_2),
    .io_outs_3(ces_7_7_io_outs_3)
  );
  Element ces_7_8 ( // @[MockArray.scala 36:52]
    .clock(ces_7_8_clock),
    .io_ins_0(ces_7_8_io_ins_0),
    .io_ins_1(ces_7_8_io_ins_1),
    .io_ins_2(ces_7_8_io_ins_2),
    .io_ins_3(ces_7_8_io_ins_3),
    .io_outs_0(ces_7_8_io_outs_0),
    .io_outs_1(ces_7_8_io_outs_1),
    .io_outs_2(ces_7_8_io_outs_2),
    .io_outs_3(ces_7_8_io_outs_3)
  );
  Element ces_7_9 ( // @[MockArray.scala 36:52]
    .clock(ces_7_9_clock),
    .io_ins_0(ces_7_9_io_ins_0),
    .io_ins_1(ces_7_9_io_ins_1),
    .io_ins_2(ces_7_9_io_ins_2),
    .io_ins_3(ces_7_9_io_ins_3),
    .io_outs_0(ces_7_9_io_outs_0),
    .io_outs_1(ces_7_9_io_outs_1),
    .io_outs_2(ces_7_9_io_outs_2),
    .io_outs_3(ces_7_9_io_outs_3)
  );
  Element ces_7_10 ( // @[MockArray.scala 36:52]
    .clock(ces_7_10_clock),
    .io_ins_0(ces_7_10_io_ins_0),
    .io_ins_1(ces_7_10_io_ins_1),
    .io_ins_2(ces_7_10_io_ins_2),
    .io_ins_3(ces_7_10_io_ins_3),
    .io_outs_0(ces_7_10_io_outs_0),
    .io_outs_1(ces_7_10_io_outs_1),
    .io_outs_2(ces_7_10_io_outs_2),
    .io_outs_3(ces_7_10_io_outs_3)
  );
  Element ces_7_11 ( // @[MockArray.scala 36:52]
    .clock(ces_7_11_clock),
    .io_ins_0(ces_7_11_io_ins_0),
    .io_ins_1(ces_7_11_io_ins_1),
    .io_ins_2(ces_7_11_io_ins_2),
    .io_ins_3(ces_7_11_io_ins_3),
    .io_outs_0(ces_7_11_io_outs_0),
    .io_outs_1(ces_7_11_io_outs_1),
    .io_outs_2(ces_7_11_io_outs_2),
    .io_outs_3(ces_7_11_io_outs_3)
  );
  Element ces_7_12 ( // @[MockArray.scala 36:52]
    .clock(ces_7_12_clock),
    .io_ins_0(ces_7_12_io_ins_0),
    .io_ins_1(ces_7_12_io_ins_1),
    .io_ins_2(ces_7_12_io_ins_2),
    .io_ins_3(ces_7_12_io_ins_3),
    .io_outs_0(ces_7_12_io_outs_0),
    .io_outs_1(ces_7_12_io_outs_1),
    .io_outs_2(ces_7_12_io_outs_2),
    .io_outs_3(ces_7_12_io_outs_3)
  );
  Element ces_7_13 ( // @[MockArray.scala 36:52]
    .clock(ces_7_13_clock),
    .io_ins_0(ces_7_13_io_ins_0),
    .io_ins_1(ces_7_13_io_ins_1),
    .io_ins_2(ces_7_13_io_ins_2),
    .io_ins_3(ces_7_13_io_ins_3),
    .io_outs_0(ces_7_13_io_outs_0),
    .io_outs_1(ces_7_13_io_outs_1),
    .io_outs_2(ces_7_13_io_outs_2),
    .io_outs_3(ces_7_13_io_outs_3)
  );
  Element ces_7_14 ( // @[MockArray.scala 36:52]
    .clock(ces_7_14_clock),
    .io_ins_0(ces_7_14_io_ins_0),
    .io_ins_1(ces_7_14_io_ins_1),
    .io_ins_2(ces_7_14_io_ins_2),
    .io_ins_3(ces_7_14_io_ins_3),
    .io_outs_0(ces_7_14_io_outs_0),
    .io_outs_1(ces_7_14_io_outs_1),
    .io_outs_2(ces_7_14_io_outs_2),
    .io_outs_3(ces_7_14_io_outs_3)
  );
  Element ces_7_15 ( // @[MockArray.scala 36:52]
    .clock(ces_7_15_clock),
    .io_ins_0(ces_7_15_io_ins_0),
    .io_ins_1(ces_7_15_io_ins_1),
    .io_ins_2(ces_7_15_io_ins_2),
    .io_ins_3(ces_7_15_io_ins_3),
    .io_outs_0(ces_7_15_io_outs_0),
    .io_outs_1(ces_7_15_io_outs_1),
    .io_outs_2(ces_7_15_io_outs_2),
    .io_outs_3(ces_7_15_io_outs_3)
  );
  Element ces_7_16 ( // @[MockArray.scala 36:52]
    .clock(ces_7_16_clock),
    .io_ins_0(ces_7_16_io_ins_0),
    .io_ins_1(ces_7_16_io_ins_1),
    .io_ins_2(ces_7_16_io_ins_2),
    .io_ins_3(ces_7_16_io_ins_3),
    .io_outs_0(ces_7_16_io_outs_0),
    .io_outs_1(ces_7_16_io_outs_1),
    .io_outs_2(ces_7_16_io_outs_2),
    .io_outs_3(ces_7_16_io_outs_3)
  );
  Element ces_7_17 ( // @[MockArray.scala 36:52]
    .clock(ces_7_17_clock),
    .io_ins_0(ces_7_17_io_ins_0),
    .io_ins_1(ces_7_17_io_ins_1),
    .io_ins_2(ces_7_17_io_ins_2),
    .io_ins_3(ces_7_17_io_ins_3),
    .io_outs_0(ces_7_17_io_outs_0),
    .io_outs_1(ces_7_17_io_outs_1),
    .io_outs_2(ces_7_17_io_outs_2),
    .io_outs_3(ces_7_17_io_outs_3)
  );
  Element ces_7_18 ( // @[MockArray.scala 36:52]
    .clock(ces_7_18_clock),
    .io_ins_0(ces_7_18_io_ins_0),
    .io_ins_1(ces_7_18_io_ins_1),
    .io_ins_2(ces_7_18_io_ins_2),
    .io_ins_3(ces_7_18_io_ins_3),
    .io_outs_0(ces_7_18_io_outs_0),
    .io_outs_1(ces_7_18_io_outs_1),
    .io_outs_2(ces_7_18_io_outs_2),
    .io_outs_3(ces_7_18_io_outs_3)
  );
  Element ces_7_19 ( // @[MockArray.scala 36:52]
    .clock(ces_7_19_clock),
    .io_ins_0(ces_7_19_io_ins_0),
    .io_ins_1(ces_7_19_io_ins_1),
    .io_ins_2(ces_7_19_io_ins_2),
    .io_ins_3(ces_7_19_io_ins_3),
    .io_outs_0(ces_7_19_io_outs_0),
    .io_outs_1(ces_7_19_io_outs_1),
    .io_outs_2(ces_7_19_io_outs_2),
    .io_outs_3(ces_7_19_io_outs_3)
  );
  Element ces_7_20 ( // @[MockArray.scala 36:52]
    .clock(ces_7_20_clock),
    .io_ins_0(ces_7_20_io_ins_0),
    .io_ins_1(ces_7_20_io_ins_1),
    .io_ins_2(ces_7_20_io_ins_2),
    .io_ins_3(ces_7_20_io_ins_3),
    .io_outs_0(ces_7_20_io_outs_0),
    .io_outs_1(ces_7_20_io_outs_1),
    .io_outs_2(ces_7_20_io_outs_2),
    .io_outs_3(ces_7_20_io_outs_3)
  );
  Element ces_7_21 ( // @[MockArray.scala 36:52]
    .clock(ces_7_21_clock),
    .io_ins_0(ces_7_21_io_ins_0),
    .io_ins_1(ces_7_21_io_ins_1),
    .io_ins_2(ces_7_21_io_ins_2),
    .io_ins_3(ces_7_21_io_ins_3),
    .io_outs_0(ces_7_21_io_outs_0),
    .io_outs_1(ces_7_21_io_outs_1),
    .io_outs_2(ces_7_21_io_outs_2),
    .io_outs_3(ces_7_21_io_outs_3)
  );
  Element ces_7_22 ( // @[MockArray.scala 36:52]
    .clock(ces_7_22_clock),
    .io_ins_0(ces_7_22_io_ins_0),
    .io_ins_1(ces_7_22_io_ins_1),
    .io_ins_2(ces_7_22_io_ins_2),
    .io_ins_3(ces_7_22_io_ins_3),
    .io_outs_0(ces_7_22_io_outs_0),
    .io_outs_1(ces_7_22_io_outs_1),
    .io_outs_2(ces_7_22_io_outs_2),
    .io_outs_3(ces_7_22_io_outs_3)
  );
  Element ces_7_23 ( // @[MockArray.scala 36:52]
    .clock(ces_7_23_clock),
    .io_ins_0(ces_7_23_io_ins_0),
    .io_ins_1(ces_7_23_io_ins_1),
    .io_ins_2(ces_7_23_io_ins_2),
    .io_ins_3(ces_7_23_io_ins_3),
    .io_outs_0(ces_7_23_io_outs_0),
    .io_outs_1(ces_7_23_io_outs_1),
    .io_outs_2(ces_7_23_io_outs_2),
    .io_outs_3(ces_7_23_io_outs_3)
  );
  Element ces_7_24 ( // @[MockArray.scala 36:52]
    .clock(ces_7_24_clock),
    .io_ins_0(ces_7_24_io_ins_0),
    .io_ins_1(ces_7_24_io_ins_1),
    .io_ins_2(ces_7_24_io_ins_2),
    .io_ins_3(ces_7_24_io_ins_3),
    .io_outs_0(ces_7_24_io_outs_0),
    .io_outs_1(ces_7_24_io_outs_1),
    .io_outs_2(ces_7_24_io_outs_2),
    .io_outs_3(ces_7_24_io_outs_3)
  );
  Element ces_7_25 ( // @[MockArray.scala 36:52]
    .clock(ces_7_25_clock),
    .io_ins_0(ces_7_25_io_ins_0),
    .io_ins_1(ces_7_25_io_ins_1),
    .io_ins_2(ces_7_25_io_ins_2),
    .io_ins_3(ces_7_25_io_ins_3),
    .io_outs_0(ces_7_25_io_outs_0),
    .io_outs_1(ces_7_25_io_outs_1),
    .io_outs_2(ces_7_25_io_outs_2),
    .io_outs_3(ces_7_25_io_outs_3)
  );
  Element ces_7_26 ( // @[MockArray.scala 36:52]
    .clock(ces_7_26_clock),
    .io_ins_0(ces_7_26_io_ins_0),
    .io_ins_1(ces_7_26_io_ins_1),
    .io_ins_2(ces_7_26_io_ins_2),
    .io_ins_3(ces_7_26_io_ins_3),
    .io_outs_0(ces_7_26_io_outs_0),
    .io_outs_1(ces_7_26_io_outs_1),
    .io_outs_2(ces_7_26_io_outs_2),
    .io_outs_3(ces_7_26_io_outs_3)
  );
  Element ces_7_27 ( // @[MockArray.scala 36:52]
    .clock(ces_7_27_clock),
    .io_ins_0(ces_7_27_io_ins_0),
    .io_ins_1(ces_7_27_io_ins_1),
    .io_ins_2(ces_7_27_io_ins_2),
    .io_ins_3(ces_7_27_io_ins_3),
    .io_outs_0(ces_7_27_io_outs_0),
    .io_outs_1(ces_7_27_io_outs_1),
    .io_outs_2(ces_7_27_io_outs_2),
    .io_outs_3(ces_7_27_io_outs_3)
  );
  Element ces_7_28 ( // @[MockArray.scala 36:52]
    .clock(ces_7_28_clock),
    .io_ins_0(ces_7_28_io_ins_0),
    .io_ins_1(ces_7_28_io_ins_1),
    .io_ins_2(ces_7_28_io_ins_2),
    .io_ins_3(ces_7_28_io_ins_3),
    .io_outs_0(ces_7_28_io_outs_0),
    .io_outs_1(ces_7_28_io_outs_1),
    .io_outs_2(ces_7_28_io_outs_2),
    .io_outs_3(ces_7_28_io_outs_3)
  );
  Element ces_7_29 ( // @[MockArray.scala 36:52]
    .clock(ces_7_29_clock),
    .io_ins_0(ces_7_29_io_ins_0),
    .io_ins_1(ces_7_29_io_ins_1),
    .io_ins_2(ces_7_29_io_ins_2),
    .io_ins_3(ces_7_29_io_ins_3),
    .io_outs_0(ces_7_29_io_outs_0),
    .io_outs_1(ces_7_29_io_outs_1),
    .io_outs_2(ces_7_29_io_outs_2),
    .io_outs_3(ces_7_29_io_outs_3)
  );
  Element ces_7_30 ( // @[MockArray.scala 36:52]
    .clock(ces_7_30_clock),
    .io_ins_0(ces_7_30_io_ins_0),
    .io_ins_1(ces_7_30_io_ins_1),
    .io_ins_2(ces_7_30_io_ins_2),
    .io_ins_3(ces_7_30_io_ins_3),
    .io_outs_0(ces_7_30_io_outs_0),
    .io_outs_1(ces_7_30_io_outs_1),
    .io_outs_2(ces_7_30_io_outs_2),
    .io_outs_3(ces_7_30_io_outs_3)
  );
  Element ces_7_31 ( // @[MockArray.scala 36:52]
    .clock(ces_7_31_clock),
    .io_ins_0(ces_7_31_io_ins_0),
    .io_ins_1(ces_7_31_io_ins_1),
    .io_ins_2(ces_7_31_io_ins_2),
    .io_ins_3(ces_7_31_io_ins_3),
    .io_outs_0(ces_7_31_io_outs_0),
    .io_outs_1(ces_7_31_io_outs_1),
    .io_outs_2(ces_7_31_io_outs_2),
    .io_outs_3(ces_7_31_io_outs_3)
  );
  Element ces_8_0 ( // @[MockArray.scala 36:52]
    .clock(ces_8_0_clock),
    .io_ins_0(ces_8_0_io_ins_0),
    .io_ins_1(ces_8_0_io_ins_1),
    .io_ins_2(ces_8_0_io_ins_2),
    .io_ins_3(ces_8_0_io_ins_3),
    .io_outs_0(ces_8_0_io_outs_0),
    .io_outs_1(ces_8_0_io_outs_1),
    .io_outs_2(ces_8_0_io_outs_2),
    .io_outs_3(ces_8_0_io_outs_3)
  );
  Element ces_8_1 ( // @[MockArray.scala 36:52]
    .clock(ces_8_1_clock),
    .io_ins_0(ces_8_1_io_ins_0),
    .io_ins_1(ces_8_1_io_ins_1),
    .io_ins_2(ces_8_1_io_ins_2),
    .io_ins_3(ces_8_1_io_ins_3),
    .io_outs_0(ces_8_1_io_outs_0),
    .io_outs_1(ces_8_1_io_outs_1),
    .io_outs_2(ces_8_1_io_outs_2),
    .io_outs_3(ces_8_1_io_outs_3)
  );
  Element ces_8_2 ( // @[MockArray.scala 36:52]
    .clock(ces_8_2_clock),
    .io_ins_0(ces_8_2_io_ins_0),
    .io_ins_1(ces_8_2_io_ins_1),
    .io_ins_2(ces_8_2_io_ins_2),
    .io_ins_3(ces_8_2_io_ins_3),
    .io_outs_0(ces_8_2_io_outs_0),
    .io_outs_1(ces_8_2_io_outs_1),
    .io_outs_2(ces_8_2_io_outs_2),
    .io_outs_3(ces_8_2_io_outs_3)
  );
  Element ces_8_3 ( // @[MockArray.scala 36:52]
    .clock(ces_8_3_clock),
    .io_ins_0(ces_8_3_io_ins_0),
    .io_ins_1(ces_8_3_io_ins_1),
    .io_ins_2(ces_8_3_io_ins_2),
    .io_ins_3(ces_8_3_io_ins_3),
    .io_outs_0(ces_8_3_io_outs_0),
    .io_outs_1(ces_8_3_io_outs_1),
    .io_outs_2(ces_8_3_io_outs_2),
    .io_outs_3(ces_8_3_io_outs_3)
  );
  Element ces_8_4 ( // @[MockArray.scala 36:52]
    .clock(ces_8_4_clock),
    .io_ins_0(ces_8_4_io_ins_0),
    .io_ins_1(ces_8_4_io_ins_1),
    .io_ins_2(ces_8_4_io_ins_2),
    .io_ins_3(ces_8_4_io_ins_3),
    .io_outs_0(ces_8_4_io_outs_0),
    .io_outs_1(ces_8_4_io_outs_1),
    .io_outs_2(ces_8_4_io_outs_2),
    .io_outs_3(ces_8_4_io_outs_3)
  );
  Element ces_8_5 ( // @[MockArray.scala 36:52]
    .clock(ces_8_5_clock),
    .io_ins_0(ces_8_5_io_ins_0),
    .io_ins_1(ces_8_5_io_ins_1),
    .io_ins_2(ces_8_5_io_ins_2),
    .io_ins_3(ces_8_5_io_ins_3),
    .io_outs_0(ces_8_5_io_outs_0),
    .io_outs_1(ces_8_5_io_outs_1),
    .io_outs_2(ces_8_5_io_outs_2),
    .io_outs_3(ces_8_5_io_outs_3)
  );
  Element ces_8_6 ( // @[MockArray.scala 36:52]
    .clock(ces_8_6_clock),
    .io_ins_0(ces_8_6_io_ins_0),
    .io_ins_1(ces_8_6_io_ins_1),
    .io_ins_2(ces_8_6_io_ins_2),
    .io_ins_3(ces_8_6_io_ins_3),
    .io_outs_0(ces_8_6_io_outs_0),
    .io_outs_1(ces_8_6_io_outs_1),
    .io_outs_2(ces_8_6_io_outs_2),
    .io_outs_3(ces_8_6_io_outs_3)
  );
  Element ces_8_7 ( // @[MockArray.scala 36:52]
    .clock(ces_8_7_clock),
    .io_ins_0(ces_8_7_io_ins_0),
    .io_ins_1(ces_8_7_io_ins_1),
    .io_ins_2(ces_8_7_io_ins_2),
    .io_ins_3(ces_8_7_io_ins_3),
    .io_outs_0(ces_8_7_io_outs_0),
    .io_outs_1(ces_8_7_io_outs_1),
    .io_outs_2(ces_8_7_io_outs_2),
    .io_outs_3(ces_8_7_io_outs_3)
  );
  Element ces_8_8 ( // @[MockArray.scala 36:52]
    .clock(ces_8_8_clock),
    .io_ins_0(ces_8_8_io_ins_0),
    .io_ins_1(ces_8_8_io_ins_1),
    .io_ins_2(ces_8_8_io_ins_2),
    .io_ins_3(ces_8_8_io_ins_3),
    .io_outs_0(ces_8_8_io_outs_0),
    .io_outs_1(ces_8_8_io_outs_1),
    .io_outs_2(ces_8_8_io_outs_2),
    .io_outs_3(ces_8_8_io_outs_3)
  );
  Element ces_8_9 ( // @[MockArray.scala 36:52]
    .clock(ces_8_9_clock),
    .io_ins_0(ces_8_9_io_ins_0),
    .io_ins_1(ces_8_9_io_ins_1),
    .io_ins_2(ces_8_9_io_ins_2),
    .io_ins_3(ces_8_9_io_ins_3),
    .io_outs_0(ces_8_9_io_outs_0),
    .io_outs_1(ces_8_9_io_outs_1),
    .io_outs_2(ces_8_9_io_outs_2),
    .io_outs_3(ces_8_9_io_outs_3)
  );
  Element ces_8_10 ( // @[MockArray.scala 36:52]
    .clock(ces_8_10_clock),
    .io_ins_0(ces_8_10_io_ins_0),
    .io_ins_1(ces_8_10_io_ins_1),
    .io_ins_2(ces_8_10_io_ins_2),
    .io_ins_3(ces_8_10_io_ins_3),
    .io_outs_0(ces_8_10_io_outs_0),
    .io_outs_1(ces_8_10_io_outs_1),
    .io_outs_2(ces_8_10_io_outs_2),
    .io_outs_3(ces_8_10_io_outs_3)
  );
  Element ces_8_11 ( // @[MockArray.scala 36:52]
    .clock(ces_8_11_clock),
    .io_ins_0(ces_8_11_io_ins_0),
    .io_ins_1(ces_8_11_io_ins_1),
    .io_ins_2(ces_8_11_io_ins_2),
    .io_ins_3(ces_8_11_io_ins_3),
    .io_outs_0(ces_8_11_io_outs_0),
    .io_outs_1(ces_8_11_io_outs_1),
    .io_outs_2(ces_8_11_io_outs_2),
    .io_outs_3(ces_8_11_io_outs_3)
  );
  Element ces_8_12 ( // @[MockArray.scala 36:52]
    .clock(ces_8_12_clock),
    .io_ins_0(ces_8_12_io_ins_0),
    .io_ins_1(ces_8_12_io_ins_1),
    .io_ins_2(ces_8_12_io_ins_2),
    .io_ins_3(ces_8_12_io_ins_3),
    .io_outs_0(ces_8_12_io_outs_0),
    .io_outs_1(ces_8_12_io_outs_1),
    .io_outs_2(ces_8_12_io_outs_2),
    .io_outs_3(ces_8_12_io_outs_3)
  );
  Element ces_8_13 ( // @[MockArray.scala 36:52]
    .clock(ces_8_13_clock),
    .io_ins_0(ces_8_13_io_ins_0),
    .io_ins_1(ces_8_13_io_ins_1),
    .io_ins_2(ces_8_13_io_ins_2),
    .io_ins_3(ces_8_13_io_ins_3),
    .io_outs_0(ces_8_13_io_outs_0),
    .io_outs_1(ces_8_13_io_outs_1),
    .io_outs_2(ces_8_13_io_outs_2),
    .io_outs_3(ces_8_13_io_outs_3)
  );
  Element ces_8_14 ( // @[MockArray.scala 36:52]
    .clock(ces_8_14_clock),
    .io_ins_0(ces_8_14_io_ins_0),
    .io_ins_1(ces_8_14_io_ins_1),
    .io_ins_2(ces_8_14_io_ins_2),
    .io_ins_3(ces_8_14_io_ins_3),
    .io_outs_0(ces_8_14_io_outs_0),
    .io_outs_1(ces_8_14_io_outs_1),
    .io_outs_2(ces_8_14_io_outs_2),
    .io_outs_3(ces_8_14_io_outs_3)
  );
  Element ces_8_15 ( // @[MockArray.scala 36:52]
    .clock(ces_8_15_clock),
    .io_ins_0(ces_8_15_io_ins_0),
    .io_ins_1(ces_8_15_io_ins_1),
    .io_ins_2(ces_8_15_io_ins_2),
    .io_ins_3(ces_8_15_io_ins_3),
    .io_outs_0(ces_8_15_io_outs_0),
    .io_outs_1(ces_8_15_io_outs_1),
    .io_outs_2(ces_8_15_io_outs_2),
    .io_outs_3(ces_8_15_io_outs_3)
  );
  Element ces_8_16 ( // @[MockArray.scala 36:52]
    .clock(ces_8_16_clock),
    .io_ins_0(ces_8_16_io_ins_0),
    .io_ins_1(ces_8_16_io_ins_1),
    .io_ins_2(ces_8_16_io_ins_2),
    .io_ins_3(ces_8_16_io_ins_3),
    .io_outs_0(ces_8_16_io_outs_0),
    .io_outs_1(ces_8_16_io_outs_1),
    .io_outs_2(ces_8_16_io_outs_2),
    .io_outs_3(ces_8_16_io_outs_3)
  );
  Element ces_8_17 ( // @[MockArray.scala 36:52]
    .clock(ces_8_17_clock),
    .io_ins_0(ces_8_17_io_ins_0),
    .io_ins_1(ces_8_17_io_ins_1),
    .io_ins_2(ces_8_17_io_ins_2),
    .io_ins_3(ces_8_17_io_ins_3),
    .io_outs_0(ces_8_17_io_outs_0),
    .io_outs_1(ces_8_17_io_outs_1),
    .io_outs_2(ces_8_17_io_outs_2),
    .io_outs_3(ces_8_17_io_outs_3)
  );
  Element ces_8_18 ( // @[MockArray.scala 36:52]
    .clock(ces_8_18_clock),
    .io_ins_0(ces_8_18_io_ins_0),
    .io_ins_1(ces_8_18_io_ins_1),
    .io_ins_2(ces_8_18_io_ins_2),
    .io_ins_3(ces_8_18_io_ins_3),
    .io_outs_0(ces_8_18_io_outs_0),
    .io_outs_1(ces_8_18_io_outs_1),
    .io_outs_2(ces_8_18_io_outs_2),
    .io_outs_3(ces_8_18_io_outs_3)
  );
  Element ces_8_19 ( // @[MockArray.scala 36:52]
    .clock(ces_8_19_clock),
    .io_ins_0(ces_8_19_io_ins_0),
    .io_ins_1(ces_8_19_io_ins_1),
    .io_ins_2(ces_8_19_io_ins_2),
    .io_ins_3(ces_8_19_io_ins_3),
    .io_outs_0(ces_8_19_io_outs_0),
    .io_outs_1(ces_8_19_io_outs_1),
    .io_outs_2(ces_8_19_io_outs_2),
    .io_outs_3(ces_8_19_io_outs_3)
  );
  Element ces_8_20 ( // @[MockArray.scala 36:52]
    .clock(ces_8_20_clock),
    .io_ins_0(ces_8_20_io_ins_0),
    .io_ins_1(ces_8_20_io_ins_1),
    .io_ins_2(ces_8_20_io_ins_2),
    .io_ins_3(ces_8_20_io_ins_3),
    .io_outs_0(ces_8_20_io_outs_0),
    .io_outs_1(ces_8_20_io_outs_1),
    .io_outs_2(ces_8_20_io_outs_2),
    .io_outs_3(ces_8_20_io_outs_3)
  );
  Element ces_8_21 ( // @[MockArray.scala 36:52]
    .clock(ces_8_21_clock),
    .io_ins_0(ces_8_21_io_ins_0),
    .io_ins_1(ces_8_21_io_ins_1),
    .io_ins_2(ces_8_21_io_ins_2),
    .io_ins_3(ces_8_21_io_ins_3),
    .io_outs_0(ces_8_21_io_outs_0),
    .io_outs_1(ces_8_21_io_outs_1),
    .io_outs_2(ces_8_21_io_outs_2),
    .io_outs_3(ces_8_21_io_outs_3)
  );
  Element ces_8_22 ( // @[MockArray.scala 36:52]
    .clock(ces_8_22_clock),
    .io_ins_0(ces_8_22_io_ins_0),
    .io_ins_1(ces_8_22_io_ins_1),
    .io_ins_2(ces_8_22_io_ins_2),
    .io_ins_3(ces_8_22_io_ins_3),
    .io_outs_0(ces_8_22_io_outs_0),
    .io_outs_1(ces_8_22_io_outs_1),
    .io_outs_2(ces_8_22_io_outs_2),
    .io_outs_3(ces_8_22_io_outs_3)
  );
  Element ces_8_23 ( // @[MockArray.scala 36:52]
    .clock(ces_8_23_clock),
    .io_ins_0(ces_8_23_io_ins_0),
    .io_ins_1(ces_8_23_io_ins_1),
    .io_ins_2(ces_8_23_io_ins_2),
    .io_ins_3(ces_8_23_io_ins_3),
    .io_outs_0(ces_8_23_io_outs_0),
    .io_outs_1(ces_8_23_io_outs_1),
    .io_outs_2(ces_8_23_io_outs_2),
    .io_outs_3(ces_8_23_io_outs_3)
  );
  Element ces_8_24 ( // @[MockArray.scala 36:52]
    .clock(ces_8_24_clock),
    .io_ins_0(ces_8_24_io_ins_0),
    .io_ins_1(ces_8_24_io_ins_1),
    .io_ins_2(ces_8_24_io_ins_2),
    .io_ins_3(ces_8_24_io_ins_3),
    .io_outs_0(ces_8_24_io_outs_0),
    .io_outs_1(ces_8_24_io_outs_1),
    .io_outs_2(ces_8_24_io_outs_2),
    .io_outs_3(ces_8_24_io_outs_3)
  );
  Element ces_8_25 ( // @[MockArray.scala 36:52]
    .clock(ces_8_25_clock),
    .io_ins_0(ces_8_25_io_ins_0),
    .io_ins_1(ces_8_25_io_ins_1),
    .io_ins_2(ces_8_25_io_ins_2),
    .io_ins_3(ces_8_25_io_ins_3),
    .io_outs_0(ces_8_25_io_outs_0),
    .io_outs_1(ces_8_25_io_outs_1),
    .io_outs_2(ces_8_25_io_outs_2),
    .io_outs_3(ces_8_25_io_outs_3)
  );
  Element ces_8_26 ( // @[MockArray.scala 36:52]
    .clock(ces_8_26_clock),
    .io_ins_0(ces_8_26_io_ins_0),
    .io_ins_1(ces_8_26_io_ins_1),
    .io_ins_2(ces_8_26_io_ins_2),
    .io_ins_3(ces_8_26_io_ins_3),
    .io_outs_0(ces_8_26_io_outs_0),
    .io_outs_1(ces_8_26_io_outs_1),
    .io_outs_2(ces_8_26_io_outs_2),
    .io_outs_3(ces_8_26_io_outs_3)
  );
  Element ces_8_27 ( // @[MockArray.scala 36:52]
    .clock(ces_8_27_clock),
    .io_ins_0(ces_8_27_io_ins_0),
    .io_ins_1(ces_8_27_io_ins_1),
    .io_ins_2(ces_8_27_io_ins_2),
    .io_ins_3(ces_8_27_io_ins_3),
    .io_outs_0(ces_8_27_io_outs_0),
    .io_outs_1(ces_8_27_io_outs_1),
    .io_outs_2(ces_8_27_io_outs_2),
    .io_outs_3(ces_8_27_io_outs_3)
  );
  Element ces_8_28 ( // @[MockArray.scala 36:52]
    .clock(ces_8_28_clock),
    .io_ins_0(ces_8_28_io_ins_0),
    .io_ins_1(ces_8_28_io_ins_1),
    .io_ins_2(ces_8_28_io_ins_2),
    .io_ins_3(ces_8_28_io_ins_3),
    .io_outs_0(ces_8_28_io_outs_0),
    .io_outs_1(ces_8_28_io_outs_1),
    .io_outs_2(ces_8_28_io_outs_2),
    .io_outs_3(ces_8_28_io_outs_3)
  );
  Element ces_8_29 ( // @[MockArray.scala 36:52]
    .clock(ces_8_29_clock),
    .io_ins_0(ces_8_29_io_ins_0),
    .io_ins_1(ces_8_29_io_ins_1),
    .io_ins_2(ces_8_29_io_ins_2),
    .io_ins_3(ces_8_29_io_ins_3),
    .io_outs_0(ces_8_29_io_outs_0),
    .io_outs_1(ces_8_29_io_outs_1),
    .io_outs_2(ces_8_29_io_outs_2),
    .io_outs_3(ces_8_29_io_outs_3)
  );
  Element ces_8_30 ( // @[MockArray.scala 36:52]
    .clock(ces_8_30_clock),
    .io_ins_0(ces_8_30_io_ins_0),
    .io_ins_1(ces_8_30_io_ins_1),
    .io_ins_2(ces_8_30_io_ins_2),
    .io_ins_3(ces_8_30_io_ins_3),
    .io_outs_0(ces_8_30_io_outs_0),
    .io_outs_1(ces_8_30_io_outs_1),
    .io_outs_2(ces_8_30_io_outs_2),
    .io_outs_3(ces_8_30_io_outs_3)
  );
  Element ces_8_31 ( // @[MockArray.scala 36:52]
    .clock(ces_8_31_clock),
    .io_ins_0(ces_8_31_io_ins_0),
    .io_ins_1(ces_8_31_io_ins_1),
    .io_ins_2(ces_8_31_io_ins_2),
    .io_ins_3(ces_8_31_io_ins_3),
    .io_outs_0(ces_8_31_io_outs_0),
    .io_outs_1(ces_8_31_io_outs_1),
    .io_outs_2(ces_8_31_io_outs_2),
    .io_outs_3(ces_8_31_io_outs_3)
  );
  Element ces_9_0 ( // @[MockArray.scala 36:52]
    .clock(ces_9_0_clock),
    .io_ins_0(ces_9_0_io_ins_0),
    .io_ins_1(ces_9_0_io_ins_1),
    .io_ins_2(ces_9_0_io_ins_2),
    .io_ins_3(ces_9_0_io_ins_3),
    .io_outs_0(ces_9_0_io_outs_0),
    .io_outs_1(ces_9_0_io_outs_1),
    .io_outs_2(ces_9_0_io_outs_2),
    .io_outs_3(ces_9_0_io_outs_3)
  );
  Element ces_9_1 ( // @[MockArray.scala 36:52]
    .clock(ces_9_1_clock),
    .io_ins_0(ces_9_1_io_ins_0),
    .io_ins_1(ces_9_1_io_ins_1),
    .io_ins_2(ces_9_1_io_ins_2),
    .io_ins_3(ces_9_1_io_ins_3),
    .io_outs_0(ces_9_1_io_outs_0),
    .io_outs_1(ces_9_1_io_outs_1),
    .io_outs_2(ces_9_1_io_outs_2),
    .io_outs_3(ces_9_1_io_outs_3)
  );
  Element ces_9_2 ( // @[MockArray.scala 36:52]
    .clock(ces_9_2_clock),
    .io_ins_0(ces_9_2_io_ins_0),
    .io_ins_1(ces_9_2_io_ins_1),
    .io_ins_2(ces_9_2_io_ins_2),
    .io_ins_3(ces_9_2_io_ins_3),
    .io_outs_0(ces_9_2_io_outs_0),
    .io_outs_1(ces_9_2_io_outs_1),
    .io_outs_2(ces_9_2_io_outs_2),
    .io_outs_3(ces_9_2_io_outs_3)
  );
  Element ces_9_3 ( // @[MockArray.scala 36:52]
    .clock(ces_9_3_clock),
    .io_ins_0(ces_9_3_io_ins_0),
    .io_ins_1(ces_9_3_io_ins_1),
    .io_ins_2(ces_9_3_io_ins_2),
    .io_ins_3(ces_9_3_io_ins_3),
    .io_outs_0(ces_9_3_io_outs_0),
    .io_outs_1(ces_9_3_io_outs_1),
    .io_outs_2(ces_9_3_io_outs_2),
    .io_outs_3(ces_9_3_io_outs_3)
  );
  Element ces_9_4 ( // @[MockArray.scala 36:52]
    .clock(ces_9_4_clock),
    .io_ins_0(ces_9_4_io_ins_0),
    .io_ins_1(ces_9_4_io_ins_1),
    .io_ins_2(ces_9_4_io_ins_2),
    .io_ins_3(ces_9_4_io_ins_3),
    .io_outs_0(ces_9_4_io_outs_0),
    .io_outs_1(ces_9_4_io_outs_1),
    .io_outs_2(ces_9_4_io_outs_2),
    .io_outs_3(ces_9_4_io_outs_3)
  );
  Element ces_9_5 ( // @[MockArray.scala 36:52]
    .clock(ces_9_5_clock),
    .io_ins_0(ces_9_5_io_ins_0),
    .io_ins_1(ces_9_5_io_ins_1),
    .io_ins_2(ces_9_5_io_ins_2),
    .io_ins_3(ces_9_5_io_ins_3),
    .io_outs_0(ces_9_5_io_outs_0),
    .io_outs_1(ces_9_5_io_outs_1),
    .io_outs_2(ces_9_5_io_outs_2),
    .io_outs_3(ces_9_5_io_outs_3)
  );
  Element ces_9_6 ( // @[MockArray.scala 36:52]
    .clock(ces_9_6_clock),
    .io_ins_0(ces_9_6_io_ins_0),
    .io_ins_1(ces_9_6_io_ins_1),
    .io_ins_2(ces_9_6_io_ins_2),
    .io_ins_3(ces_9_6_io_ins_3),
    .io_outs_0(ces_9_6_io_outs_0),
    .io_outs_1(ces_9_6_io_outs_1),
    .io_outs_2(ces_9_6_io_outs_2),
    .io_outs_3(ces_9_6_io_outs_3)
  );
  Element ces_9_7 ( // @[MockArray.scala 36:52]
    .clock(ces_9_7_clock),
    .io_ins_0(ces_9_7_io_ins_0),
    .io_ins_1(ces_9_7_io_ins_1),
    .io_ins_2(ces_9_7_io_ins_2),
    .io_ins_3(ces_9_7_io_ins_3),
    .io_outs_0(ces_9_7_io_outs_0),
    .io_outs_1(ces_9_7_io_outs_1),
    .io_outs_2(ces_9_7_io_outs_2),
    .io_outs_3(ces_9_7_io_outs_3)
  );
  Element ces_9_8 ( // @[MockArray.scala 36:52]
    .clock(ces_9_8_clock),
    .io_ins_0(ces_9_8_io_ins_0),
    .io_ins_1(ces_9_8_io_ins_1),
    .io_ins_2(ces_9_8_io_ins_2),
    .io_ins_3(ces_9_8_io_ins_3),
    .io_outs_0(ces_9_8_io_outs_0),
    .io_outs_1(ces_9_8_io_outs_1),
    .io_outs_2(ces_9_8_io_outs_2),
    .io_outs_3(ces_9_8_io_outs_3)
  );
  Element ces_9_9 ( // @[MockArray.scala 36:52]
    .clock(ces_9_9_clock),
    .io_ins_0(ces_9_9_io_ins_0),
    .io_ins_1(ces_9_9_io_ins_1),
    .io_ins_2(ces_9_9_io_ins_2),
    .io_ins_3(ces_9_9_io_ins_3),
    .io_outs_0(ces_9_9_io_outs_0),
    .io_outs_1(ces_9_9_io_outs_1),
    .io_outs_2(ces_9_9_io_outs_2),
    .io_outs_3(ces_9_9_io_outs_3)
  );
  Element ces_9_10 ( // @[MockArray.scala 36:52]
    .clock(ces_9_10_clock),
    .io_ins_0(ces_9_10_io_ins_0),
    .io_ins_1(ces_9_10_io_ins_1),
    .io_ins_2(ces_9_10_io_ins_2),
    .io_ins_3(ces_9_10_io_ins_3),
    .io_outs_0(ces_9_10_io_outs_0),
    .io_outs_1(ces_9_10_io_outs_1),
    .io_outs_2(ces_9_10_io_outs_2),
    .io_outs_3(ces_9_10_io_outs_3)
  );
  Element ces_9_11 ( // @[MockArray.scala 36:52]
    .clock(ces_9_11_clock),
    .io_ins_0(ces_9_11_io_ins_0),
    .io_ins_1(ces_9_11_io_ins_1),
    .io_ins_2(ces_9_11_io_ins_2),
    .io_ins_3(ces_9_11_io_ins_3),
    .io_outs_0(ces_9_11_io_outs_0),
    .io_outs_1(ces_9_11_io_outs_1),
    .io_outs_2(ces_9_11_io_outs_2),
    .io_outs_3(ces_9_11_io_outs_3)
  );
  Element ces_9_12 ( // @[MockArray.scala 36:52]
    .clock(ces_9_12_clock),
    .io_ins_0(ces_9_12_io_ins_0),
    .io_ins_1(ces_9_12_io_ins_1),
    .io_ins_2(ces_9_12_io_ins_2),
    .io_ins_3(ces_9_12_io_ins_3),
    .io_outs_0(ces_9_12_io_outs_0),
    .io_outs_1(ces_9_12_io_outs_1),
    .io_outs_2(ces_9_12_io_outs_2),
    .io_outs_3(ces_9_12_io_outs_3)
  );
  Element ces_9_13 ( // @[MockArray.scala 36:52]
    .clock(ces_9_13_clock),
    .io_ins_0(ces_9_13_io_ins_0),
    .io_ins_1(ces_9_13_io_ins_1),
    .io_ins_2(ces_9_13_io_ins_2),
    .io_ins_3(ces_9_13_io_ins_3),
    .io_outs_0(ces_9_13_io_outs_0),
    .io_outs_1(ces_9_13_io_outs_1),
    .io_outs_2(ces_9_13_io_outs_2),
    .io_outs_3(ces_9_13_io_outs_3)
  );
  Element ces_9_14 ( // @[MockArray.scala 36:52]
    .clock(ces_9_14_clock),
    .io_ins_0(ces_9_14_io_ins_0),
    .io_ins_1(ces_9_14_io_ins_1),
    .io_ins_2(ces_9_14_io_ins_2),
    .io_ins_3(ces_9_14_io_ins_3),
    .io_outs_0(ces_9_14_io_outs_0),
    .io_outs_1(ces_9_14_io_outs_1),
    .io_outs_2(ces_9_14_io_outs_2),
    .io_outs_3(ces_9_14_io_outs_3)
  );
  Element ces_9_15 ( // @[MockArray.scala 36:52]
    .clock(ces_9_15_clock),
    .io_ins_0(ces_9_15_io_ins_0),
    .io_ins_1(ces_9_15_io_ins_1),
    .io_ins_2(ces_9_15_io_ins_2),
    .io_ins_3(ces_9_15_io_ins_3),
    .io_outs_0(ces_9_15_io_outs_0),
    .io_outs_1(ces_9_15_io_outs_1),
    .io_outs_2(ces_9_15_io_outs_2),
    .io_outs_3(ces_9_15_io_outs_3)
  );
  Element ces_9_16 ( // @[MockArray.scala 36:52]
    .clock(ces_9_16_clock),
    .io_ins_0(ces_9_16_io_ins_0),
    .io_ins_1(ces_9_16_io_ins_1),
    .io_ins_2(ces_9_16_io_ins_2),
    .io_ins_3(ces_9_16_io_ins_3),
    .io_outs_0(ces_9_16_io_outs_0),
    .io_outs_1(ces_9_16_io_outs_1),
    .io_outs_2(ces_9_16_io_outs_2),
    .io_outs_3(ces_9_16_io_outs_3)
  );
  Element ces_9_17 ( // @[MockArray.scala 36:52]
    .clock(ces_9_17_clock),
    .io_ins_0(ces_9_17_io_ins_0),
    .io_ins_1(ces_9_17_io_ins_1),
    .io_ins_2(ces_9_17_io_ins_2),
    .io_ins_3(ces_9_17_io_ins_3),
    .io_outs_0(ces_9_17_io_outs_0),
    .io_outs_1(ces_9_17_io_outs_1),
    .io_outs_2(ces_9_17_io_outs_2),
    .io_outs_3(ces_9_17_io_outs_3)
  );
  Element ces_9_18 ( // @[MockArray.scala 36:52]
    .clock(ces_9_18_clock),
    .io_ins_0(ces_9_18_io_ins_0),
    .io_ins_1(ces_9_18_io_ins_1),
    .io_ins_2(ces_9_18_io_ins_2),
    .io_ins_3(ces_9_18_io_ins_3),
    .io_outs_0(ces_9_18_io_outs_0),
    .io_outs_1(ces_9_18_io_outs_1),
    .io_outs_2(ces_9_18_io_outs_2),
    .io_outs_3(ces_9_18_io_outs_3)
  );
  Element ces_9_19 ( // @[MockArray.scala 36:52]
    .clock(ces_9_19_clock),
    .io_ins_0(ces_9_19_io_ins_0),
    .io_ins_1(ces_9_19_io_ins_1),
    .io_ins_2(ces_9_19_io_ins_2),
    .io_ins_3(ces_9_19_io_ins_3),
    .io_outs_0(ces_9_19_io_outs_0),
    .io_outs_1(ces_9_19_io_outs_1),
    .io_outs_2(ces_9_19_io_outs_2),
    .io_outs_3(ces_9_19_io_outs_3)
  );
  Element ces_9_20 ( // @[MockArray.scala 36:52]
    .clock(ces_9_20_clock),
    .io_ins_0(ces_9_20_io_ins_0),
    .io_ins_1(ces_9_20_io_ins_1),
    .io_ins_2(ces_9_20_io_ins_2),
    .io_ins_3(ces_9_20_io_ins_3),
    .io_outs_0(ces_9_20_io_outs_0),
    .io_outs_1(ces_9_20_io_outs_1),
    .io_outs_2(ces_9_20_io_outs_2),
    .io_outs_3(ces_9_20_io_outs_3)
  );
  Element ces_9_21 ( // @[MockArray.scala 36:52]
    .clock(ces_9_21_clock),
    .io_ins_0(ces_9_21_io_ins_0),
    .io_ins_1(ces_9_21_io_ins_1),
    .io_ins_2(ces_9_21_io_ins_2),
    .io_ins_3(ces_9_21_io_ins_3),
    .io_outs_0(ces_9_21_io_outs_0),
    .io_outs_1(ces_9_21_io_outs_1),
    .io_outs_2(ces_9_21_io_outs_2),
    .io_outs_3(ces_9_21_io_outs_3)
  );
  Element ces_9_22 ( // @[MockArray.scala 36:52]
    .clock(ces_9_22_clock),
    .io_ins_0(ces_9_22_io_ins_0),
    .io_ins_1(ces_9_22_io_ins_1),
    .io_ins_2(ces_9_22_io_ins_2),
    .io_ins_3(ces_9_22_io_ins_3),
    .io_outs_0(ces_9_22_io_outs_0),
    .io_outs_1(ces_9_22_io_outs_1),
    .io_outs_2(ces_9_22_io_outs_2),
    .io_outs_3(ces_9_22_io_outs_3)
  );
  Element ces_9_23 ( // @[MockArray.scala 36:52]
    .clock(ces_9_23_clock),
    .io_ins_0(ces_9_23_io_ins_0),
    .io_ins_1(ces_9_23_io_ins_1),
    .io_ins_2(ces_9_23_io_ins_2),
    .io_ins_3(ces_9_23_io_ins_3),
    .io_outs_0(ces_9_23_io_outs_0),
    .io_outs_1(ces_9_23_io_outs_1),
    .io_outs_2(ces_9_23_io_outs_2),
    .io_outs_3(ces_9_23_io_outs_3)
  );
  Element ces_9_24 ( // @[MockArray.scala 36:52]
    .clock(ces_9_24_clock),
    .io_ins_0(ces_9_24_io_ins_0),
    .io_ins_1(ces_9_24_io_ins_1),
    .io_ins_2(ces_9_24_io_ins_2),
    .io_ins_3(ces_9_24_io_ins_3),
    .io_outs_0(ces_9_24_io_outs_0),
    .io_outs_1(ces_9_24_io_outs_1),
    .io_outs_2(ces_9_24_io_outs_2),
    .io_outs_3(ces_9_24_io_outs_3)
  );
  Element ces_9_25 ( // @[MockArray.scala 36:52]
    .clock(ces_9_25_clock),
    .io_ins_0(ces_9_25_io_ins_0),
    .io_ins_1(ces_9_25_io_ins_1),
    .io_ins_2(ces_9_25_io_ins_2),
    .io_ins_3(ces_9_25_io_ins_3),
    .io_outs_0(ces_9_25_io_outs_0),
    .io_outs_1(ces_9_25_io_outs_1),
    .io_outs_2(ces_9_25_io_outs_2),
    .io_outs_3(ces_9_25_io_outs_3)
  );
  Element ces_9_26 ( // @[MockArray.scala 36:52]
    .clock(ces_9_26_clock),
    .io_ins_0(ces_9_26_io_ins_0),
    .io_ins_1(ces_9_26_io_ins_1),
    .io_ins_2(ces_9_26_io_ins_2),
    .io_ins_3(ces_9_26_io_ins_3),
    .io_outs_0(ces_9_26_io_outs_0),
    .io_outs_1(ces_9_26_io_outs_1),
    .io_outs_2(ces_9_26_io_outs_2),
    .io_outs_3(ces_9_26_io_outs_3)
  );
  Element ces_9_27 ( // @[MockArray.scala 36:52]
    .clock(ces_9_27_clock),
    .io_ins_0(ces_9_27_io_ins_0),
    .io_ins_1(ces_9_27_io_ins_1),
    .io_ins_2(ces_9_27_io_ins_2),
    .io_ins_3(ces_9_27_io_ins_3),
    .io_outs_0(ces_9_27_io_outs_0),
    .io_outs_1(ces_9_27_io_outs_1),
    .io_outs_2(ces_9_27_io_outs_2),
    .io_outs_3(ces_9_27_io_outs_3)
  );
  Element ces_9_28 ( // @[MockArray.scala 36:52]
    .clock(ces_9_28_clock),
    .io_ins_0(ces_9_28_io_ins_0),
    .io_ins_1(ces_9_28_io_ins_1),
    .io_ins_2(ces_9_28_io_ins_2),
    .io_ins_3(ces_9_28_io_ins_3),
    .io_outs_0(ces_9_28_io_outs_0),
    .io_outs_1(ces_9_28_io_outs_1),
    .io_outs_2(ces_9_28_io_outs_2),
    .io_outs_3(ces_9_28_io_outs_3)
  );
  Element ces_9_29 ( // @[MockArray.scala 36:52]
    .clock(ces_9_29_clock),
    .io_ins_0(ces_9_29_io_ins_0),
    .io_ins_1(ces_9_29_io_ins_1),
    .io_ins_2(ces_9_29_io_ins_2),
    .io_ins_3(ces_9_29_io_ins_3),
    .io_outs_0(ces_9_29_io_outs_0),
    .io_outs_1(ces_9_29_io_outs_1),
    .io_outs_2(ces_9_29_io_outs_2),
    .io_outs_3(ces_9_29_io_outs_3)
  );
  Element ces_9_30 ( // @[MockArray.scala 36:52]
    .clock(ces_9_30_clock),
    .io_ins_0(ces_9_30_io_ins_0),
    .io_ins_1(ces_9_30_io_ins_1),
    .io_ins_2(ces_9_30_io_ins_2),
    .io_ins_3(ces_9_30_io_ins_3),
    .io_outs_0(ces_9_30_io_outs_0),
    .io_outs_1(ces_9_30_io_outs_1),
    .io_outs_2(ces_9_30_io_outs_2),
    .io_outs_3(ces_9_30_io_outs_3)
  );
  Element ces_9_31 ( // @[MockArray.scala 36:52]
    .clock(ces_9_31_clock),
    .io_ins_0(ces_9_31_io_ins_0),
    .io_ins_1(ces_9_31_io_ins_1),
    .io_ins_2(ces_9_31_io_ins_2),
    .io_ins_3(ces_9_31_io_ins_3),
    .io_outs_0(ces_9_31_io_outs_0),
    .io_outs_1(ces_9_31_io_outs_1),
    .io_outs_2(ces_9_31_io_outs_2),
    .io_outs_3(ces_9_31_io_outs_3)
  );
  Element ces_10_0 ( // @[MockArray.scala 36:52]
    .clock(ces_10_0_clock),
    .io_ins_0(ces_10_0_io_ins_0),
    .io_ins_1(ces_10_0_io_ins_1),
    .io_ins_2(ces_10_0_io_ins_2),
    .io_ins_3(ces_10_0_io_ins_3),
    .io_outs_0(ces_10_0_io_outs_0),
    .io_outs_1(ces_10_0_io_outs_1),
    .io_outs_2(ces_10_0_io_outs_2),
    .io_outs_3(ces_10_0_io_outs_3)
  );
  Element ces_10_1 ( // @[MockArray.scala 36:52]
    .clock(ces_10_1_clock),
    .io_ins_0(ces_10_1_io_ins_0),
    .io_ins_1(ces_10_1_io_ins_1),
    .io_ins_2(ces_10_1_io_ins_2),
    .io_ins_3(ces_10_1_io_ins_3),
    .io_outs_0(ces_10_1_io_outs_0),
    .io_outs_1(ces_10_1_io_outs_1),
    .io_outs_2(ces_10_1_io_outs_2),
    .io_outs_3(ces_10_1_io_outs_3)
  );
  Element ces_10_2 ( // @[MockArray.scala 36:52]
    .clock(ces_10_2_clock),
    .io_ins_0(ces_10_2_io_ins_0),
    .io_ins_1(ces_10_2_io_ins_1),
    .io_ins_2(ces_10_2_io_ins_2),
    .io_ins_3(ces_10_2_io_ins_3),
    .io_outs_0(ces_10_2_io_outs_0),
    .io_outs_1(ces_10_2_io_outs_1),
    .io_outs_2(ces_10_2_io_outs_2),
    .io_outs_3(ces_10_2_io_outs_3)
  );
  Element ces_10_3 ( // @[MockArray.scala 36:52]
    .clock(ces_10_3_clock),
    .io_ins_0(ces_10_3_io_ins_0),
    .io_ins_1(ces_10_3_io_ins_1),
    .io_ins_2(ces_10_3_io_ins_2),
    .io_ins_3(ces_10_3_io_ins_3),
    .io_outs_0(ces_10_3_io_outs_0),
    .io_outs_1(ces_10_3_io_outs_1),
    .io_outs_2(ces_10_3_io_outs_2),
    .io_outs_3(ces_10_3_io_outs_3)
  );
  Element ces_10_4 ( // @[MockArray.scala 36:52]
    .clock(ces_10_4_clock),
    .io_ins_0(ces_10_4_io_ins_0),
    .io_ins_1(ces_10_4_io_ins_1),
    .io_ins_2(ces_10_4_io_ins_2),
    .io_ins_3(ces_10_4_io_ins_3),
    .io_outs_0(ces_10_4_io_outs_0),
    .io_outs_1(ces_10_4_io_outs_1),
    .io_outs_2(ces_10_4_io_outs_2),
    .io_outs_3(ces_10_4_io_outs_3)
  );
  Element ces_10_5 ( // @[MockArray.scala 36:52]
    .clock(ces_10_5_clock),
    .io_ins_0(ces_10_5_io_ins_0),
    .io_ins_1(ces_10_5_io_ins_1),
    .io_ins_2(ces_10_5_io_ins_2),
    .io_ins_3(ces_10_5_io_ins_3),
    .io_outs_0(ces_10_5_io_outs_0),
    .io_outs_1(ces_10_5_io_outs_1),
    .io_outs_2(ces_10_5_io_outs_2),
    .io_outs_3(ces_10_5_io_outs_3)
  );
  Element ces_10_6 ( // @[MockArray.scala 36:52]
    .clock(ces_10_6_clock),
    .io_ins_0(ces_10_6_io_ins_0),
    .io_ins_1(ces_10_6_io_ins_1),
    .io_ins_2(ces_10_6_io_ins_2),
    .io_ins_3(ces_10_6_io_ins_3),
    .io_outs_0(ces_10_6_io_outs_0),
    .io_outs_1(ces_10_6_io_outs_1),
    .io_outs_2(ces_10_6_io_outs_2),
    .io_outs_3(ces_10_6_io_outs_3)
  );
  Element ces_10_7 ( // @[MockArray.scala 36:52]
    .clock(ces_10_7_clock),
    .io_ins_0(ces_10_7_io_ins_0),
    .io_ins_1(ces_10_7_io_ins_1),
    .io_ins_2(ces_10_7_io_ins_2),
    .io_ins_3(ces_10_7_io_ins_3),
    .io_outs_0(ces_10_7_io_outs_0),
    .io_outs_1(ces_10_7_io_outs_1),
    .io_outs_2(ces_10_7_io_outs_2),
    .io_outs_3(ces_10_7_io_outs_3)
  );
  Element ces_10_8 ( // @[MockArray.scala 36:52]
    .clock(ces_10_8_clock),
    .io_ins_0(ces_10_8_io_ins_0),
    .io_ins_1(ces_10_8_io_ins_1),
    .io_ins_2(ces_10_8_io_ins_2),
    .io_ins_3(ces_10_8_io_ins_3),
    .io_outs_0(ces_10_8_io_outs_0),
    .io_outs_1(ces_10_8_io_outs_1),
    .io_outs_2(ces_10_8_io_outs_2),
    .io_outs_3(ces_10_8_io_outs_3)
  );
  Element ces_10_9 ( // @[MockArray.scala 36:52]
    .clock(ces_10_9_clock),
    .io_ins_0(ces_10_9_io_ins_0),
    .io_ins_1(ces_10_9_io_ins_1),
    .io_ins_2(ces_10_9_io_ins_2),
    .io_ins_3(ces_10_9_io_ins_3),
    .io_outs_0(ces_10_9_io_outs_0),
    .io_outs_1(ces_10_9_io_outs_1),
    .io_outs_2(ces_10_9_io_outs_2),
    .io_outs_3(ces_10_9_io_outs_3)
  );
  Element ces_10_10 ( // @[MockArray.scala 36:52]
    .clock(ces_10_10_clock),
    .io_ins_0(ces_10_10_io_ins_0),
    .io_ins_1(ces_10_10_io_ins_1),
    .io_ins_2(ces_10_10_io_ins_2),
    .io_ins_3(ces_10_10_io_ins_3),
    .io_outs_0(ces_10_10_io_outs_0),
    .io_outs_1(ces_10_10_io_outs_1),
    .io_outs_2(ces_10_10_io_outs_2),
    .io_outs_3(ces_10_10_io_outs_3)
  );
  Element ces_10_11 ( // @[MockArray.scala 36:52]
    .clock(ces_10_11_clock),
    .io_ins_0(ces_10_11_io_ins_0),
    .io_ins_1(ces_10_11_io_ins_1),
    .io_ins_2(ces_10_11_io_ins_2),
    .io_ins_3(ces_10_11_io_ins_3),
    .io_outs_0(ces_10_11_io_outs_0),
    .io_outs_1(ces_10_11_io_outs_1),
    .io_outs_2(ces_10_11_io_outs_2),
    .io_outs_3(ces_10_11_io_outs_3)
  );
  Element ces_10_12 ( // @[MockArray.scala 36:52]
    .clock(ces_10_12_clock),
    .io_ins_0(ces_10_12_io_ins_0),
    .io_ins_1(ces_10_12_io_ins_1),
    .io_ins_2(ces_10_12_io_ins_2),
    .io_ins_3(ces_10_12_io_ins_3),
    .io_outs_0(ces_10_12_io_outs_0),
    .io_outs_1(ces_10_12_io_outs_1),
    .io_outs_2(ces_10_12_io_outs_2),
    .io_outs_3(ces_10_12_io_outs_3)
  );
  Element ces_10_13 ( // @[MockArray.scala 36:52]
    .clock(ces_10_13_clock),
    .io_ins_0(ces_10_13_io_ins_0),
    .io_ins_1(ces_10_13_io_ins_1),
    .io_ins_2(ces_10_13_io_ins_2),
    .io_ins_3(ces_10_13_io_ins_3),
    .io_outs_0(ces_10_13_io_outs_0),
    .io_outs_1(ces_10_13_io_outs_1),
    .io_outs_2(ces_10_13_io_outs_2),
    .io_outs_3(ces_10_13_io_outs_3)
  );
  Element ces_10_14 ( // @[MockArray.scala 36:52]
    .clock(ces_10_14_clock),
    .io_ins_0(ces_10_14_io_ins_0),
    .io_ins_1(ces_10_14_io_ins_1),
    .io_ins_2(ces_10_14_io_ins_2),
    .io_ins_3(ces_10_14_io_ins_3),
    .io_outs_0(ces_10_14_io_outs_0),
    .io_outs_1(ces_10_14_io_outs_1),
    .io_outs_2(ces_10_14_io_outs_2),
    .io_outs_3(ces_10_14_io_outs_3)
  );
  Element ces_10_15 ( // @[MockArray.scala 36:52]
    .clock(ces_10_15_clock),
    .io_ins_0(ces_10_15_io_ins_0),
    .io_ins_1(ces_10_15_io_ins_1),
    .io_ins_2(ces_10_15_io_ins_2),
    .io_ins_3(ces_10_15_io_ins_3),
    .io_outs_0(ces_10_15_io_outs_0),
    .io_outs_1(ces_10_15_io_outs_1),
    .io_outs_2(ces_10_15_io_outs_2),
    .io_outs_3(ces_10_15_io_outs_3)
  );
  Element ces_10_16 ( // @[MockArray.scala 36:52]
    .clock(ces_10_16_clock),
    .io_ins_0(ces_10_16_io_ins_0),
    .io_ins_1(ces_10_16_io_ins_1),
    .io_ins_2(ces_10_16_io_ins_2),
    .io_ins_3(ces_10_16_io_ins_3),
    .io_outs_0(ces_10_16_io_outs_0),
    .io_outs_1(ces_10_16_io_outs_1),
    .io_outs_2(ces_10_16_io_outs_2),
    .io_outs_3(ces_10_16_io_outs_3)
  );
  Element ces_10_17 ( // @[MockArray.scala 36:52]
    .clock(ces_10_17_clock),
    .io_ins_0(ces_10_17_io_ins_0),
    .io_ins_1(ces_10_17_io_ins_1),
    .io_ins_2(ces_10_17_io_ins_2),
    .io_ins_3(ces_10_17_io_ins_3),
    .io_outs_0(ces_10_17_io_outs_0),
    .io_outs_1(ces_10_17_io_outs_1),
    .io_outs_2(ces_10_17_io_outs_2),
    .io_outs_3(ces_10_17_io_outs_3)
  );
  Element ces_10_18 ( // @[MockArray.scala 36:52]
    .clock(ces_10_18_clock),
    .io_ins_0(ces_10_18_io_ins_0),
    .io_ins_1(ces_10_18_io_ins_1),
    .io_ins_2(ces_10_18_io_ins_2),
    .io_ins_3(ces_10_18_io_ins_3),
    .io_outs_0(ces_10_18_io_outs_0),
    .io_outs_1(ces_10_18_io_outs_1),
    .io_outs_2(ces_10_18_io_outs_2),
    .io_outs_3(ces_10_18_io_outs_3)
  );
  Element ces_10_19 ( // @[MockArray.scala 36:52]
    .clock(ces_10_19_clock),
    .io_ins_0(ces_10_19_io_ins_0),
    .io_ins_1(ces_10_19_io_ins_1),
    .io_ins_2(ces_10_19_io_ins_2),
    .io_ins_3(ces_10_19_io_ins_3),
    .io_outs_0(ces_10_19_io_outs_0),
    .io_outs_1(ces_10_19_io_outs_1),
    .io_outs_2(ces_10_19_io_outs_2),
    .io_outs_3(ces_10_19_io_outs_3)
  );
  Element ces_10_20 ( // @[MockArray.scala 36:52]
    .clock(ces_10_20_clock),
    .io_ins_0(ces_10_20_io_ins_0),
    .io_ins_1(ces_10_20_io_ins_1),
    .io_ins_2(ces_10_20_io_ins_2),
    .io_ins_3(ces_10_20_io_ins_3),
    .io_outs_0(ces_10_20_io_outs_0),
    .io_outs_1(ces_10_20_io_outs_1),
    .io_outs_2(ces_10_20_io_outs_2),
    .io_outs_3(ces_10_20_io_outs_3)
  );
  Element ces_10_21 ( // @[MockArray.scala 36:52]
    .clock(ces_10_21_clock),
    .io_ins_0(ces_10_21_io_ins_0),
    .io_ins_1(ces_10_21_io_ins_1),
    .io_ins_2(ces_10_21_io_ins_2),
    .io_ins_3(ces_10_21_io_ins_3),
    .io_outs_0(ces_10_21_io_outs_0),
    .io_outs_1(ces_10_21_io_outs_1),
    .io_outs_2(ces_10_21_io_outs_2),
    .io_outs_3(ces_10_21_io_outs_3)
  );
  Element ces_10_22 ( // @[MockArray.scala 36:52]
    .clock(ces_10_22_clock),
    .io_ins_0(ces_10_22_io_ins_0),
    .io_ins_1(ces_10_22_io_ins_1),
    .io_ins_2(ces_10_22_io_ins_2),
    .io_ins_3(ces_10_22_io_ins_3),
    .io_outs_0(ces_10_22_io_outs_0),
    .io_outs_1(ces_10_22_io_outs_1),
    .io_outs_2(ces_10_22_io_outs_2),
    .io_outs_3(ces_10_22_io_outs_3)
  );
  Element ces_10_23 ( // @[MockArray.scala 36:52]
    .clock(ces_10_23_clock),
    .io_ins_0(ces_10_23_io_ins_0),
    .io_ins_1(ces_10_23_io_ins_1),
    .io_ins_2(ces_10_23_io_ins_2),
    .io_ins_3(ces_10_23_io_ins_3),
    .io_outs_0(ces_10_23_io_outs_0),
    .io_outs_1(ces_10_23_io_outs_1),
    .io_outs_2(ces_10_23_io_outs_2),
    .io_outs_3(ces_10_23_io_outs_3)
  );
  Element ces_10_24 ( // @[MockArray.scala 36:52]
    .clock(ces_10_24_clock),
    .io_ins_0(ces_10_24_io_ins_0),
    .io_ins_1(ces_10_24_io_ins_1),
    .io_ins_2(ces_10_24_io_ins_2),
    .io_ins_3(ces_10_24_io_ins_3),
    .io_outs_0(ces_10_24_io_outs_0),
    .io_outs_1(ces_10_24_io_outs_1),
    .io_outs_2(ces_10_24_io_outs_2),
    .io_outs_3(ces_10_24_io_outs_3)
  );
  Element ces_10_25 ( // @[MockArray.scala 36:52]
    .clock(ces_10_25_clock),
    .io_ins_0(ces_10_25_io_ins_0),
    .io_ins_1(ces_10_25_io_ins_1),
    .io_ins_2(ces_10_25_io_ins_2),
    .io_ins_3(ces_10_25_io_ins_3),
    .io_outs_0(ces_10_25_io_outs_0),
    .io_outs_1(ces_10_25_io_outs_1),
    .io_outs_2(ces_10_25_io_outs_2),
    .io_outs_3(ces_10_25_io_outs_3)
  );
  Element ces_10_26 ( // @[MockArray.scala 36:52]
    .clock(ces_10_26_clock),
    .io_ins_0(ces_10_26_io_ins_0),
    .io_ins_1(ces_10_26_io_ins_1),
    .io_ins_2(ces_10_26_io_ins_2),
    .io_ins_3(ces_10_26_io_ins_3),
    .io_outs_0(ces_10_26_io_outs_0),
    .io_outs_1(ces_10_26_io_outs_1),
    .io_outs_2(ces_10_26_io_outs_2),
    .io_outs_3(ces_10_26_io_outs_3)
  );
  Element ces_10_27 ( // @[MockArray.scala 36:52]
    .clock(ces_10_27_clock),
    .io_ins_0(ces_10_27_io_ins_0),
    .io_ins_1(ces_10_27_io_ins_1),
    .io_ins_2(ces_10_27_io_ins_2),
    .io_ins_3(ces_10_27_io_ins_3),
    .io_outs_0(ces_10_27_io_outs_0),
    .io_outs_1(ces_10_27_io_outs_1),
    .io_outs_2(ces_10_27_io_outs_2),
    .io_outs_3(ces_10_27_io_outs_3)
  );
  Element ces_10_28 ( // @[MockArray.scala 36:52]
    .clock(ces_10_28_clock),
    .io_ins_0(ces_10_28_io_ins_0),
    .io_ins_1(ces_10_28_io_ins_1),
    .io_ins_2(ces_10_28_io_ins_2),
    .io_ins_3(ces_10_28_io_ins_3),
    .io_outs_0(ces_10_28_io_outs_0),
    .io_outs_1(ces_10_28_io_outs_1),
    .io_outs_2(ces_10_28_io_outs_2),
    .io_outs_3(ces_10_28_io_outs_3)
  );
  Element ces_10_29 ( // @[MockArray.scala 36:52]
    .clock(ces_10_29_clock),
    .io_ins_0(ces_10_29_io_ins_0),
    .io_ins_1(ces_10_29_io_ins_1),
    .io_ins_2(ces_10_29_io_ins_2),
    .io_ins_3(ces_10_29_io_ins_3),
    .io_outs_0(ces_10_29_io_outs_0),
    .io_outs_1(ces_10_29_io_outs_1),
    .io_outs_2(ces_10_29_io_outs_2),
    .io_outs_3(ces_10_29_io_outs_3)
  );
  Element ces_10_30 ( // @[MockArray.scala 36:52]
    .clock(ces_10_30_clock),
    .io_ins_0(ces_10_30_io_ins_0),
    .io_ins_1(ces_10_30_io_ins_1),
    .io_ins_2(ces_10_30_io_ins_2),
    .io_ins_3(ces_10_30_io_ins_3),
    .io_outs_0(ces_10_30_io_outs_0),
    .io_outs_1(ces_10_30_io_outs_1),
    .io_outs_2(ces_10_30_io_outs_2),
    .io_outs_3(ces_10_30_io_outs_3)
  );
  Element ces_10_31 ( // @[MockArray.scala 36:52]
    .clock(ces_10_31_clock),
    .io_ins_0(ces_10_31_io_ins_0),
    .io_ins_1(ces_10_31_io_ins_1),
    .io_ins_2(ces_10_31_io_ins_2),
    .io_ins_3(ces_10_31_io_ins_3),
    .io_outs_0(ces_10_31_io_outs_0),
    .io_outs_1(ces_10_31_io_outs_1),
    .io_outs_2(ces_10_31_io_outs_2),
    .io_outs_3(ces_10_31_io_outs_3)
  );
  Element ces_11_0 ( // @[MockArray.scala 36:52]
    .clock(ces_11_0_clock),
    .io_ins_0(ces_11_0_io_ins_0),
    .io_ins_1(ces_11_0_io_ins_1),
    .io_ins_2(ces_11_0_io_ins_2),
    .io_ins_3(ces_11_0_io_ins_3),
    .io_outs_0(ces_11_0_io_outs_0),
    .io_outs_1(ces_11_0_io_outs_1),
    .io_outs_2(ces_11_0_io_outs_2),
    .io_outs_3(ces_11_0_io_outs_3)
  );
  Element ces_11_1 ( // @[MockArray.scala 36:52]
    .clock(ces_11_1_clock),
    .io_ins_0(ces_11_1_io_ins_0),
    .io_ins_1(ces_11_1_io_ins_1),
    .io_ins_2(ces_11_1_io_ins_2),
    .io_ins_3(ces_11_1_io_ins_3),
    .io_outs_0(ces_11_1_io_outs_0),
    .io_outs_1(ces_11_1_io_outs_1),
    .io_outs_2(ces_11_1_io_outs_2),
    .io_outs_3(ces_11_1_io_outs_3)
  );
  Element ces_11_2 ( // @[MockArray.scala 36:52]
    .clock(ces_11_2_clock),
    .io_ins_0(ces_11_2_io_ins_0),
    .io_ins_1(ces_11_2_io_ins_1),
    .io_ins_2(ces_11_2_io_ins_2),
    .io_ins_3(ces_11_2_io_ins_3),
    .io_outs_0(ces_11_2_io_outs_0),
    .io_outs_1(ces_11_2_io_outs_1),
    .io_outs_2(ces_11_2_io_outs_2),
    .io_outs_3(ces_11_2_io_outs_3)
  );
  Element ces_11_3 ( // @[MockArray.scala 36:52]
    .clock(ces_11_3_clock),
    .io_ins_0(ces_11_3_io_ins_0),
    .io_ins_1(ces_11_3_io_ins_1),
    .io_ins_2(ces_11_3_io_ins_2),
    .io_ins_3(ces_11_3_io_ins_3),
    .io_outs_0(ces_11_3_io_outs_0),
    .io_outs_1(ces_11_3_io_outs_1),
    .io_outs_2(ces_11_3_io_outs_2),
    .io_outs_3(ces_11_3_io_outs_3)
  );
  Element ces_11_4 ( // @[MockArray.scala 36:52]
    .clock(ces_11_4_clock),
    .io_ins_0(ces_11_4_io_ins_0),
    .io_ins_1(ces_11_4_io_ins_1),
    .io_ins_2(ces_11_4_io_ins_2),
    .io_ins_3(ces_11_4_io_ins_3),
    .io_outs_0(ces_11_4_io_outs_0),
    .io_outs_1(ces_11_4_io_outs_1),
    .io_outs_2(ces_11_4_io_outs_2),
    .io_outs_3(ces_11_4_io_outs_3)
  );
  Element ces_11_5 ( // @[MockArray.scala 36:52]
    .clock(ces_11_5_clock),
    .io_ins_0(ces_11_5_io_ins_0),
    .io_ins_1(ces_11_5_io_ins_1),
    .io_ins_2(ces_11_5_io_ins_2),
    .io_ins_3(ces_11_5_io_ins_3),
    .io_outs_0(ces_11_5_io_outs_0),
    .io_outs_1(ces_11_5_io_outs_1),
    .io_outs_2(ces_11_5_io_outs_2),
    .io_outs_3(ces_11_5_io_outs_3)
  );
  Element ces_11_6 ( // @[MockArray.scala 36:52]
    .clock(ces_11_6_clock),
    .io_ins_0(ces_11_6_io_ins_0),
    .io_ins_1(ces_11_6_io_ins_1),
    .io_ins_2(ces_11_6_io_ins_2),
    .io_ins_3(ces_11_6_io_ins_3),
    .io_outs_0(ces_11_6_io_outs_0),
    .io_outs_1(ces_11_6_io_outs_1),
    .io_outs_2(ces_11_6_io_outs_2),
    .io_outs_3(ces_11_6_io_outs_3)
  );
  Element ces_11_7 ( // @[MockArray.scala 36:52]
    .clock(ces_11_7_clock),
    .io_ins_0(ces_11_7_io_ins_0),
    .io_ins_1(ces_11_7_io_ins_1),
    .io_ins_2(ces_11_7_io_ins_2),
    .io_ins_3(ces_11_7_io_ins_3),
    .io_outs_0(ces_11_7_io_outs_0),
    .io_outs_1(ces_11_7_io_outs_1),
    .io_outs_2(ces_11_7_io_outs_2),
    .io_outs_3(ces_11_7_io_outs_3)
  );
  Element ces_11_8 ( // @[MockArray.scala 36:52]
    .clock(ces_11_8_clock),
    .io_ins_0(ces_11_8_io_ins_0),
    .io_ins_1(ces_11_8_io_ins_1),
    .io_ins_2(ces_11_8_io_ins_2),
    .io_ins_3(ces_11_8_io_ins_3),
    .io_outs_0(ces_11_8_io_outs_0),
    .io_outs_1(ces_11_8_io_outs_1),
    .io_outs_2(ces_11_8_io_outs_2),
    .io_outs_3(ces_11_8_io_outs_3)
  );
  Element ces_11_9 ( // @[MockArray.scala 36:52]
    .clock(ces_11_9_clock),
    .io_ins_0(ces_11_9_io_ins_0),
    .io_ins_1(ces_11_9_io_ins_1),
    .io_ins_2(ces_11_9_io_ins_2),
    .io_ins_3(ces_11_9_io_ins_3),
    .io_outs_0(ces_11_9_io_outs_0),
    .io_outs_1(ces_11_9_io_outs_1),
    .io_outs_2(ces_11_9_io_outs_2),
    .io_outs_3(ces_11_9_io_outs_3)
  );
  Element ces_11_10 ( // @[MockArray.scala 36:52]
    .clock(ces_11_10_clock),
    .io_ins_0(ces_11_10_io_ins_0),
    .io_ins_1(ces_11_10_io_ins_1),
    .io_ins_2(ces_11_10_io_ins_2),
    .io_ins_3(ces_11_10_io_ins_3),
    .io_outs_0(ces_11_10_io_outs_0),
    .io_outs_1(ces_11_10_io_outs_1),
    .io_outs_2(ces_11_10_io_outs_2),
    .io_outs_3(ces_11_10_io_outs_3)
  );
  Element ces_11_11 ( // @[MockArray.scala 36:52]
    .clock(ces_11_11_clock),
    .io_ins_0(ces_11_11_io_ins_0),
    .io_ins_1(ces_11_11_io_ins_1),
    .io_ins_2(ces_11_11_io_ins_2),
    .io_ins_3(ces_11_11_io_ins_3),
    .io_outs_0(ces_11_11_io_outs_0),
    .io_outs_1(ces_11_11_io_outs_1),
    .io_outs_2(ces_11_11_io_outs_2),
    .io_outs_3(ces_11_11_io_outs_3)
  );
  Element ces_11_12 ( // @[MockArray.scala 36:52]
    .clock(ces_11_12_clock),
    .io_ins_0(ces_11_12_io_ins_0),
    .io_ins_1(ces_11_12_io_ins_1),
    .io_ins_2(ces_11_12_io_ins_2),
    .io_ins_3(ces_11_12_io_ins_3),
    .io_outs_0(ces_11_12_io_outs_0),
    .io_outs_1(ces_11_12_io_outs_1),
    .io_outs_2(ces_11_12_io_outs_2),
    .io_outs_3(ces_11_12_io_outs_3)
  );
  Element ces_11_13 ( // @[MockArray.scala 36:52]
    .clock(ces_11_13_clock),
    .io_ins_0(ces_11_13_io_ins_0),
    .io_ins_1(ces_11_13_io_ins_1),
    .io_ins_2(ces_11_13_io_ins_2),
    .io_ins_3(ces_11_13_io_ins_3),
    .io_outs_0(ces_11_13_io_outs_0),
    .io_outs_1(ces_11_13_io_outs_1),
    .io_outs_2(ces_11_13_io_outs_2),
    .io_outs_3(ces_11_13_io_outs_3)
  );
  Element ces_11_14 ( // @[MockArray.scala 36:52]
    .clock(ces_11_14_clock),
    .io_ins_0(ces_11_14_io_ins_0),
    .io_ins_1(ces_11_14_io_ins_1),
    .io_ins_2(ces_11_14_io_ins_2),
    .io_ins_3(ces_11_14_io_ins_3),
    .io_outs_0(ces_11_14_io_outs_0),
    .io_outs_1(ces_11_14_io_outs_1),
    .io_outs_2(ces_11_14_io_outs_2),
    .io_outs_3(ces_11_14_io_outs_3)
  );
  Element ces_11_15 ( // @[MockArray.scala 36:52]
    .clock(ces_11_15_clock),
    .io_ins_0(ces_11_15_io_ins_0),
    .io_ins_1(ces_11_15_io_ins_1),
    .io_ins_2(ces_11_15_io_ins_2),
    .io_ins_3(ces_11_15_io_ins_3),
    .io_outs_0(ces_11_15_io_outs_0),
    .io_outs_1(ces_11_15_io_outs_1),
    .io_outs_2(ces_11_15_io_outs_2),
    .io_outs_3(ces_11_15_io_outs_3)
  );
  Element ces_11_16 ( // @[MockArray.scala 36:52]
    .clock(ces_11_16_clock),
    .io_ins_0(ces_11_16_io_ins_0),
    .io_ins_1(ces_11_16_io_ins_1),
    .io_ins_2(ces_11_16_io_ins_2),
    .io_ins_3(ces_11_16_io_ins_3),
    .io_outs_0(ces_11_16_io_outs_0),
    .io_outs_1(ces_11_16_io_outs_1),
    .io_outs_2(ces_11_16_io_outs_2),
    .io_outs_3(ces_11_16_io_outs_3)
  );
  Element ces_11_17 ( // @[MockArray.scala 36:52]
    .clock(ces_11_17_clock),
    .io_ins_0(ces_11_17_io_ins_0),
    .io_ins_1(ces_11_17_io_ins_1),
    .io_ins_2(ces_11_17_io_ins_2),
    .io_ins_3(ces_11_17_io_ins_3),
    .io_outs_0(ces_11_17_io_outs_0),
    .io_outs_1(ces_11_17_io_outs_1),
    .io_outs_2(ces_11_17_io_outs_2),
    .io_outs_3(ces_11_17_io_outs_3)
  );
  Element ces_11_18 ( // @[MockArray.scala 36:52]
    .clock(ces_11_18_clock),
    .io_ins_0(ces_11_18_io_ins_0),
    .io_ins_1(ces_11_18_io_ins_1),
    .io_ins_2(ces_11_18_io_ins_2),
    .io_ins_3(ces_11_18_io_ins_3),
    .io_outs_0(ces_11_18_io_outs_0),
    .io_outs_1(ces_11_18_io_outs_1),
    .io_outs_2(ces_11_18_io_outs_2),
    .io_outs_3(ces_11_18_io_outs_3)
  );
  Element ces_11_19 ( // @[MockArray.scala 36:52]
    .clock(ces_11_19_clock),
    .io_ins_0(ces_11_19_io_ins_0),
    .io_ins_1(ces_11_19_io_ins_1),
    .io_ins_2(ces_11_19_io_ins_2),
    .io_ins_3(ces_11_19_io_ins_3),
    .io_outs_0(ces_11_19_io_outs_0),
    .io_outs_1(ces_11_19_io_outs_1),
    .io_outs_2(ces_11_19_io_outs_2),
    .io_outs_3(ces_11_19_io_outs_3)
  );
  Element ces_11_20 ( // @[MockArray.scala 36:52]
    .clock(ces_11_20_clock),
    .io_ins_0(ces_11_20_io_ins_0),
    .io_ins_1(ces_11_20_io_ins_1),
    .io_ins_2(ces_11_20_io_ins_2),
    .io_ins_3(ces_11_20_io_ins_3),
    .io_outs_0(ces_11_20_io_outs_0),
    .io_outs_1(ces_11_20_io_outs_1),
    .io_outs_2(ces_11_20_io_outs_2),
    .io_outs_3(ces_11_20_io_outs_3)
  );
  Element ces_11_21 ( // @[MockArray.scala 36:52]
    .clock(ces_11_21_clock),
    .io_ins_0(ces_11_21_io_ins_0),
    .io_ins_1(ces_11_21_io_ins_1),
    .io_ins_2(ces_11_21_io_ins_2),
    .io_ins_3(ces_11_21_io_ins_3),
    .io_outs_0(ces_11_21_io_outs_0),
    .io_outs_1(ces_11_21_io_outs_1),
    .io_outs_2(ces_11_21_io_outs_2),
    .io_outs_3(ces_11_21_io_outs_3)
  );
  Element ces_11_22 ( // @[MockArray.scala 36:52]
    .clock(ces_11_22_clock),
    .io_ins_0(ces_11_22_io_ins_0),
    .io_ins_1(ces_11_22_io_ins_1),
    .io_ins_2(ces_11_22_io_ins_2),
    .io_ins_3(ces_11_22_io_ins_3),
    .io_outs_0(ces_11_22_io_outs_0),
    .io_outs_1(ces_11_22_io_outs_1),
    .io_outs_2(ces_11_22_io_outs_2),
    .io_outs_3(ces_11_22_io_outs_3)
  );
  Element ces_11_23 ( // @[MockArray.scala 36:52]
    .clock(ces_11_23_clock),
    .io_ins_0(ces_11_23_io_ins_0),
    .io_ins_1(ces_11_23_io_ins_1),
    .io_ins_2(ces_11_23_io_ins_2),
    .io_ins_3(ces_11_23_io_ins_3),
    .io_outs_0(ces_11_23_io_outs_0),
    .io_outs_1(ces_11_23_io_outs_1),
    .io_outs_2(ces_11_23_io_outs_2),
    .io_outs_3(ces_11_23_io_outs_3)
  );
  Element ces_11_24 ( // @[MockArray.scala 36:52]
    .clock(ces_11_24_clock),
    .io_ins_0(ces_11_24_io_ins_0),
    .io_ins_1(ces_11_24_io_ins_1),
    .io_ins_2(ces_11_24_io_ins_2),
    .io_ins_3(ces_11_24_io_ins_3),
    .io_outs_0(ces_11_24_io_outs_0),
    .io_outs_1(ces_11_24_io_outs_1),
    .io_outs_2(ces_11_24_io_outs_2),
    .io_outs_3(ces_11_24_io_outs_3)
  );
  Element ces_11_25 ( // @[MockArray.scala 36:52]
    .clock(ces_11_25_clock),
    .io_ins_0(ces_11_25_io_ins_0),
    .io_ins_1(ces_11_25_io_ins_1),
    .io_ins_2(ces_11_25_io_ins_2),
    .io_ins_3(ces_11_25_io_ins_3),
    .io_outs_0(ces_11_25_io_outs_0),
    .io_outs_1(ces_11_25_io_outs_1),
    .io_outs_2(ces_11_25_io_outs_2),
    .io_outs_3(ces_11_25_io_outs_3)
  );
  Element ces_11_26 ( // @[MockArray.scala 36:52]
    .clock(ces_11_26_clock),
    .io_ins_0(ces_11_26_io_ins_0),
    .io_ins_1(ces_11_26_io_ins_1),
    .io_ins_2(ces_11_26_io_ins_2),
    .io_ins_3(ces_11_26_io_ins_3),
    .io_outs_0(ces_11_26_io_outs_0),
    .io_outs_1(ces_11_26_io_outs_1),
    .io_outs_2(ces_11_26_io_outs_2),
    .io_outs_3(ces_11_26_io_outs_3)
  );
  Element ces_11_27 ( // @[MockArray.scala 36:52]
    .clock(ces_11_27_clock),
    .io_ins_0(ces_11_27_io_ins_0),
    .io_ins_1(ces_11_27_io_ins_1),
    .io_ins_2(ces_11_27_io_ins_2),
    .io_ins_3(ces_11_27_io_ins_3),
    .io_outs_0(ces_11_27_io_outs_0),
    .io_outs_1(ces_11_27_io_outs_1),
    .io_outs_2(ces_11_27_io_outs_2),
    .io_outs_3(ces_11_27_io_outs_3)
  );
  Element ces_11_28 ( // @[MockArray.scala 36:52]
    .clock(ces_11_28_clock),
    .io_ins_0(ces_11_28_io_ins_0),
    .io_ins_1(ces_11_28_io_ins_1),
    .io_ins_2(ces_11_28_io_ins_2),
    .io_ins_3(ces_11_28_io_ins_3),
    .io_outs_0(ces_11_28_io_outs_0),
    .io_outs_1(ces_11_28_io_outs_1),
    .io_outs_2(ces_11_28_io_outs_2),
    .io_outs_3(ces_11_28_io_outs_3)
  );
  Element ces_11_29 ( // @[MockArray.scala 36:52]
    .clock(ces_11_29_clock),
    .io_ins_0(ces_11_29_io_ins_0),
    .io_ins_1(ces_11_29_io_ins_1),
    .io_ins_2(ces_11_29_io_ins_2),
    .io_ins_3(ces_11_29_io_ins_3),
    .io_outs_0(ces_11_29_io_outs_0),
    .io_outs_1(ces_11_29_io_outs_1),
    .io_outs_2(ces_11_29_io_outs_2),
    .io_outs_3(ces_11_29_io_outs_3)
  );
  Element ces_11_30 ( // @[MockArray.scala 36:52]
    .clock(ces_11_30_clock),
    .io_ins_0(ces_11_30_io_ins_0),
    .io_ins_1(ces_11_30_io_ins_1),
    .io_ins_2(ces_11_30_io_ins_2),
    .io_ins_3(ces_11_30_io_ins_3),
    .io_outs_0(ces_11_30_io_outs_0),
    .io_outs_1(ces_11_30_io_outs_1),
    .io_outs_2(ces_11_30_io_outs_2),
    .io_outs_3(ces_11_30_io_outs_3)
  );
  Element ces_11_31 ( // @[MockArray.scala 36:52]
    .clock(ces_11_31_clock),
    .io_ins_0(ces_11_31_io_ins_0),
    .io_ins_1(ces_11_31_io_ins_1),
    .io_ins_2(ces_11_31_io_ins_2),
    .io_ins_3(ces_11_31_io_ins_3),
    .io_outs_0(ces_11_31_io_outs_0),
    .io_outs_1(ces_11_31_io_outs_1),
    .io_outs_2(ces_11_31_io_outs_2),
    .io_outs_3(ces_11_31_io_outs_3)
  );
  Element ces_12_0 ( // @[MockArray.scala 36:52]
    .clock(ces_12_0_clock),
    .io_ins_0(ces_12_0_io_ins_0),
    .io_ins_1(ces_12_0_io_ins_1),
    .io_ins_2(ces_12_0_io_ins_2),
    .io_ins_3(ces_12_0_io_ins_3),
    .io_outs_0(ces_12_0_io_outs_0),
    .io_outs_1(ces_12_0_io_outs_1),
    .io_outs_2(ces_12_0_io_outs_2),
    .io_outs_3(ces_12_0_io_outs_3)
  );
  Element ces_12_1 ( // @[MockArray.scala 36:52]
    .clock(ces_12_1_clock),
    .io_ins_0(ces_12_1_io_ins_0),
    .io_ins_1(ces_12_1_io_ins_1),
    .io_ins_2(ces_12_1_io_ins_2),
    .io_ins_3(ces_12_1_io_ins_3),
    .io_outs_0(ces_12_1_io_outs_0),
    .io_outs_1(ces_12_1_io_outs_1),
    .io_outs_2(ces_12_1_io_outs_2),
    .io_outs_3(ces_12_1_io_outs_3)
  );
  Element ces_12_2 ( // @[MockArray.scala 36:52]
    .clock(ces_12_2_clock),
    .io_ins_0(ces_12_2_io_ins_0),
    .io_ins_1(ces_12_2_io_ins_1),
    .io_ins_2(ces_12_2_io_ins_2),
    .io_ins_3(ces_12_2_io_ins_3),
    .io_outs_0(ces_12_2_io_outs_0),
    .io_outs_1(ces_12_2_io_outs_1),
    .io_outs_2(ces_12_2_io_outs_2),
    .io_outs_3(ces_12_2_io_outs_3)
  );
  Element ces_12_3 ( // @[MockArray.scala 36:52]
    .clock(ces_12_3_clock),
    .io_ins_0(ces_12_3_io_ins_0),
    .io_ins_1(ces_12_3_io_ins_1),
    .io_ins_2(ces_12_3_io_ins_2),
    .io_ins_3(ces_12_3_io_ins_3),
    .io_outs_0(ces_12_3_io_outs_0),
    .io_outs_1(ces_12_3_io_outs_1),
    .io_outs_2(ces_12_3_io_outs_2),
    .io_outs_3(ces_12_3_io_outs_3)
  );
  Element ces_12_4 ( // @[MockArray.scala 36:52]
    .clock(ces_12_4_clock),
    .io_ins_0(ces_12_4_io_ins_0),
    .io_ins_1(ces_12_4_io_ins_1),
    .io_ins_2(ces_12_4_io_ins_2),
    .io_ins_3(ces_12_4_io_ins_3),
    .io_outs_0(ces_12_4_io_outs_0),
    .io_outs_1(ces_12_4_io_outs_1),
    .io_outs_2(ces_12_4_io_outs_2),
    .io_outs_3(ces_12_4_io_outs_3)
  );
  Element ces_12_5 ( // @[MockArray.scala 36:52]
    .clock(ces_12_5_clock),
    .io_ins_0(ces_12_5_io_ins_0),
    .io_ins_1(ces_12_5_io_ins_1),
    .io_ins_2(ces_12_5_io_ins_2),
    .io_ins_3(ces_12_5_io_ins_3),
    .io_outs_0(ces_12_5_io_outs_0),
    .io_outs_1(ces_12_5_io_outs_1),
    .io_outs_2(ces_12_5_io_outs_2),
    .io_outs_3(ces_12_5_io_outs_3)
  );
  Element ces_12_6 ( // @[MockArray.scala 36:52]
    .clock(ces_12_6_clock),
    .io_ins_0(ces_12_6_io_ins_0),
    .io_ins_1(ces_12_6_io_ins_1),
    .io_ins_2(ces_12_6_io_ins_2),
    .io_ins_3(ces_12_6_io_ins_3),
    .io_outs_0(ces_12_6_io_outs_0),
    .io_outs_1(ces_12_6_io_outs_1),
    .io_outs_2(ces_12_6_io_outs_2),
    .io_outs_3(ces_12_6_io_outs_3)
  );
  Element ces_12_7 ( // @[MockArray.scala 36:52]
    .clock(ces_12_7_clock),
    .io_ins_0(ces_12_7_io_ins_0),
    .io_ins_1(ces_12_7_io_ins_1),
    .io_ins_2(ces_12_7_io_ins_2),
    .io_ins_3(ces_12_7_io_ins_3),
    .io_outs_0(ces_12_7_io_outs_0),
    .io_outs_1(ces_12_7_io_outs_1),
    .io_outs_2(ces_12_7_io_outs_2),
    .io_outs_3(ces_12_7_io_outs_3)
  );
  Element ces_12_8 ( // @[MockArray.scala 36:52]
    .clock(ces_12_8_clock),
    .io_ins_0(ces_12_8_io_ins_0),
    .io_ins_1(ces_12_8_io_ins_1),
    .io_ins_2(ces_12_8_io_ins_2),
    .io_ins_3(ces_12_8_io_ins_3),
    .io_outs_0(ces_12_8_io_outs_0),
    .io_outs_1(ces_12_8_io_outs_1),
    .io_outs_2(ces_12_8_io_outs_2),
    .io_outs_3(ces_12_8_io_outs_3)
  );
  Element ces_12_9 ( // @[MockArray.scala 36:52]
    .clock(ces_12_9_clock),
    .io_ins_0(ces_12_9_io_ins_0),
    .io_ins_1(ces_12_9_io_ins_1),
    .io_ins_2(ces_12_9_io_ins_2),
    .io_ins_3(ces_12_9_io_ins_3),
    .io_outs_0(ces_12_9_io_outs_0),
    .io_outs_1(ces_12_9_io_outs_1),
    .io_outs_2(ces_12_9_io_outs_2),
    .io_outs_3(ces_12_9_io_outs_3)
  );
  Element ces_12_10 ( // @[MockArray.scala 36:52]
    .clock(ces_12_10_clock),
    .io_ins_0(ces_12_10_io_ins_0),
    .io_ins_1(ces_12_10_io_ins_1),
    .io_ins_2(ces_12_10_io_ins_2),
    .io_ins_3(ces_12_10_io_ins_3),
    .io_outs_0(ces_12_10_io_outs_0),
    .io_outs_1(ces_12_10_io_outs_1),
    .io_outs_2(ces_12_10_io_outs_2),
    .io_outs_3(ces_12_10_io_outs_3)
  );
  Element ces_12_11 ( // @[MockArray.scala 36:52]
    .clock(ces_12_11_clock),
    .io_ins_0(ces_12_11_io_ins_0),
    .io_ins_1(ces_12_11_io_ins_1),
    .io_ins_2(ces_12_11_io_ins_2),
    .io_ins_3(ces_12_11_io_ins_3),
    .io_outs_0(ces_12_11_io_outs_0),
    .io_outs_1(ces_12_11_io_outs_1),
    .io_outs_2(ces_12_11_io_outs_2),
    .io_outs_3(ces_12_11_io_outs_3)
  );
  Element ces_12_12 ( // @[MockArray.scala 36:52]
    .clock(ces_12_12_clock),
    .io_ins_0(ces_12_12_io_ins_0),
    .io_ins_1(ces_12_12_io_ins_1),
    .io_ins_2(ces_12_12_io_ins_2),
    .io_ins_3(ces_12_12_io_ins_3),
    .io_outs_0(ces_12_12_io_outs_0),
    .io_outs_1(ces_12_12_io_outs_1),
    .io_outs_2(ces_12_12_io_outs_2),
    .io_outs_3(ces_12_12_io_outs_3)
  );
  Element ces_12_13 ( // @[MockArray.scala 36:52]
    .clock(ces_12_13_clock),
    .io_ins_0(ces_12_13_io_ins_0),
    .io_ins_1(ces_12_13_io_ins_1),
    .io_ins_2(ces_12_13_io_ins_2),
    .io_ins_3(ces_12_13_io_ins_3),
    .io_outs_0(ces_12_13_io_outs_0),
    .io_outs_1(ces_12_13_io_outs_1),
    .io_outs_2(ces_12_13_io_outs_2),
    .io_outs_3(ces_12_13_io_outs_3)
  );
  Element ces_12_14 ( // @[MockArray.scala 36:52]
    .clock(ces_12_14_clock),
    .io_ins_0(ces_12_14_io_ins_0),
    .io_ins_1(ces_12_14_io_ins_1),
    .io_ins_2(ces_12_14_io_ins_2),
    .io_ins_3(ces_12_14_io_ins_3),
    .io_outs_0(ces_12_14_io_outs_0),
    .io_outs_1(ces_12_14_io_outs_1),
    .io_outs_2(ces_12_14_io_outs_2),
    .io_outs_3(ces_12_14_io_outs_3)
  );
  Element ces_12_15 ( // @[MockArray.scala 36:52]
    .clock(ces_12_15_clock),
    .io_ins_0(ces_12_15_io_ins_0),
    .io_ins_1(ces_12_15_io_ins_1),
    .io_ins_2(ces_12_15_io_ins_2),
    .io_ins_3(ces_12_15_io_ins_3),
    .io_outs_0(ces_12_15_io_outs_0),
    .io_outs_1(ces_12_15_io_outs_1),
    .io_outs_2(ces_12_15_io_outs_2),
    .io_outs_3(ces_12_15_io_outs_3)
  );
  Element ces_12_16 ( // @[MockArray.scala 36:52]
    .clock(ces_12_16_clock),
    .io_ins_0(ces_12_16_io_ins_0),
    .io_ins_1(ces_12_16_io_ins_1),
    .io_ins_2(ces_12_16_io_ins_2),
    .io_ins_3(ces_12_16_io_ins_3),
    .io_outs_0(ces_12_16_io_outs_0),
    .io_outs_1(ces_12_16_io_outs_1),
    .io_outs_2(ces_12_16_io_outs_2),
    .io_outs_3(ces_12_16_io_outs_3)
  );
  Element ces_12_17 ( // @[MockArray.scala 36:52]
    .clock(ces_12_17_clock),
    .io_ins_0(ces_12_17_io_ins_0),
    .io_ins_1(ces_12_17_io_ins_1),
    .io_ins_2(ces_12_17_io_ins_2),
    .io_ins_3(ces_12_17_io_ins_3),
    .io_outs_0(ces_12_17_io_outs_0),
    .io_outs_1(ces_12_17_io_outs_1),
    .io_outs_2(ces_12_17_io_outs_2),
    .io_outs_3(ces_12_17_io_outs_3)
  );
  Element ces_12_18 ( // @[MockArray.scala 36:52]
    .clock(ces_12_18_clock),
    .io_ins_0(ces_12_18_io_ins_0),
    .io_ins_1(ces_12_18_io_ins_1),
    .io_ins_2(ces_12_18_io_ins_2),
    .io_ins_3(ces_12_18_io_ins_3),
    .io_outs_0(ces_12_18_io_outs_0),
    .io_outs_1(ces_12_18_io_outs_1),
    .io_outs_2(ces_12_18_io_outs_2),
    .io_outs_3(ces_12_18_io_outs_3)
  );
  Element ces_12_19 ( // @[MockArray.scala 36:52]
    .clock(ces_12_19_clock),
    .io_ins_0(ces_12_19_io_ins_0),
    .io_ins_1(ces_12_19_io_ins_1),
    .io_ins_2(ces_12_19_io_ins_2),
    .io_ins_3(ces_12_19_io_ins_3),
    .io_outs_0(ces_12_19_io_outs_0),
    .io_outs_1(ces_12_19_io_outs_1),
    .io_outs_2(ces_12_19_io_outs_2),
    .io_outs_3(ces_12_19_io_outs_3)
  );
  Element ces_12_20 ( // @[MockArray.scala 36:52]
    .clock(ces_12_20_clock),
    .io_ins_0(ces_12_20_io_ins_0),
    .io_ins_1(ces_12_20_io_ins_1),
    .io_ins_2(ces_12_20_io_ins_2),
    .io_ins_3(ces_12_20_io_ins_3),
    .io_outs_0(ces_12_20_io_outs_0),
    .io_outs_1(ces_12_20_io_outs_1),
    .io_outs_2(ces_12_20_io_outs_2),
    .io_outs_3(ces_12_20_io_outs_3)
  );
  Element ces_12_21 ( // @[MockArray.scala 36:52]
    .clock(ces_12_21_clock),
    .io_ins_0(ces_12_21_io_ins_0),
    .io_ins_1(ces_12_21_io_ins_1),
    .io_ins_2(ces_12_21_io_ins_2),
    .io_ins_3(ces_12_21_io_ins_3),
    .io_outs_0(ces_12_21_io_outs_0),
    .io_outs_1(ces_12_21_io_outs_1),
    .io_outs_2(ces_12_21_io_outs_2),
    .io_outs_3(ces_12_21_io_outs_3)
  );
  Element ces_12_22 ( // @[MockArray.scala 36:52]
    .clock(ces_12_22_clock),
    .io_ins_0(ces_12_22_io_ins_0),
    .io_ins_1(ces_12_22_io_ins_1),
    .io_ins_2(ces_12_22_io_ins_2),
    .io_ins_3(ces_12_22_io_ins_3),
    .io_outs_0(ces_12_22_io_outs_0),
    .io_outs_1(ces_12_22_io_outs_1),
    .io_outs_2(ces_12_22_io_outs_2),
    .io_outs_3(ces_12_22_io_outs_3)
  );
  Element ces_12_23 ( // @[MockArray.scala 36:52]
    .clock(ces_12_23_clock),
    .io_ins_0(ces_12_23_io_ins_0),
    .io_ins_1(ces_12_23_io_ins_1),
    .io_ins_2(ces_12_23_io_ins_2),
    .io_ins_3(ces_12_23_io_ins_3),
    .io_outs_0(ces_12_23_io_outs_0),
    .io_outs_1(ces_12_23_io_outs_1),
    .io_outs_2(ces_12_23_io_outs_2),
    .io_outs_3(ces_12_23_io_outs_3)
  );
  Element ces_12_24 ( // @[MockArray.scala 36:52]
    .clock(ces_12_24_clock),
    .io_ins_0(ces_12_24_io_ins_0),
    .io_ins_1(ces_12_24_io_ins_1),
    .io_ins_2(ces_12_24_io_ins_2),
    .io_ins_3(ces_12_24_io_ins_3),
    .io_outs_0(ces_12_24_io_outs_0),
    .io_outs_1(ces_12_24_io_outs_1),
    .io_outs_2(ces_12_24_io_outs_2),
    .io_outs_3(ces_12_24_io_outs_3)
  );
  Element ces_12_25 ( // @[MockArray.scala 36:52]
    .clock(ces_12_25_clock),
    .io_ins_0(ces_12_25_io_ins_0),
    .io_ins_1(ces_12_25_io_ins_1),
    .io_ins_2(ces_12_25_io_ins_2),
    .io_ins_3(ces_12_25_io_ins_3),
    .io_outs_0(ces_12_25_io_outs_0),
    .io_outs_1(ces_12_25_io_outs_1),
    .io_outs_2(ces_12_25_io_outs_2),
    .io_outs_3(ces_12_25_io_outs_3)
  );
  Element ces_12_26 ( // @[MockArray.scala 36:52]
    .clock(ces_12_26_clock),
    .io_ins_0(ces_12_26_io_ins_0),
    .io_ins_1(ces_12_26_io_ins_1),
    .io_ins_2(ces_12_26_io_ins_2),
    .io_ins_3(ces_12_26_io_ins_3),
    .io_outs_0(ces_12_26_io_outs_0),
    .io_outs_1(ces_12_26_io_outs_1),
    .io_outs_2(ces_12_26_io_outs_2),
    .io_outs_3(ces_12_26_io_outs_3)
  );
  Element ces_12_27 ( // @[MockArray.scala 36:52]
    .clock(ces_12_27_clock),
    .io_ins_0(ces_12_27_io_ins_0),
    .io_ins_1(ces_12_27_io_ins_1),
    .io_ins_2(ces_12_27_io_ins_2),
    .io_ins_3(ces_12_27_io_ins_3),
    .io_outs_0(ces_12_27_io_outs_0),
    .io_outs_1(ces_12_27_io_outs_1),
    .io_outs_2(ces_12_27_io_outs_2),
    .io_outs_3(ces_12_27_io_outs_3)
  );
  Element ces_12_28 ( // @[MockArray.scala 36:52]
    .clock(ces_12_28_clock),
    .io_ins_0(ces_12_28_io_ins_0),
    .io_ins_1(ces_12_28_io_ins_1),
    .io_ins_2(ces_12_28_io_ins_2),
    .io_ins_3(ces_12_28_io_ins_3),
    .io_outs_0(ces_12_28_io_outs_0),
    .io_outs_1(ces_12_28_io_outs_1),
    .io_outs_2(ces_12_28_io_outs_2),
    .io_outs_3(ces_12_28_io_outs_3)
  );
  Element ces_12_29 ( // @[MockArray.scala 36:52]
    .clock(ces_12_29_clock),
    .io_ins_0(ces_12_29_io_ins_0),
    .io_ins_1(ces_12_29_io_ins_1),
    .io_ins_2(ces_12_29_io_ins_2),
    .io_ins_3(ces_12_29_io_ins_3),
    .io_outs_0(ces_12_29_io_outs_0),
    .io_outs_1(ces_12_29_io_outs_1),
    .io_outs_2(ces_12_29_io_outs_2),
    .io_outs_3(ces_12_29_io_outs_3)
  );
  Element ces_12_30 ( // @[MockArray.scala 36:52]
    .clock(ces_12_30_clock),
    .io_ins_0(ces_12_30_io_ins_0),
    .io_ins_1(ces_12_30_io_ins_1),
    .io_ins_2(ces_12_30_io_ins_2),
    .io_ins_3(ces_12_30_io_ins_3),
    .io_outs_0(ces_12_30_io_outs_0),
    .io_outs_1(ces_12_30_io_outs_1),
    .io_outs_2(ces_12_30_io_outs_2),
    .io_outs_3(ces_12_30_io_outs_3)
  );
  Element ces_12_31 ( // @[MockArray.scala 36:52]
    .clock(ces_12_31_clock),
    .io_ins_0(ces_12_31_io_ins_0),
    .io_ins_1(ces_12_31_io_ins_1),
    .io_ins_2(ces_12_31_io_ins_2),
    .io_ins_3(ces_12_31_io_ins_3),
    .io_outs_0(ces_12_31_io_outs_0),
    .io_outs_1(ces_12_31_io_outs_1),
    .io_outs_2(ces_12_31_io_outs_2),
    .io_outs_3(ces_12_31_io_outs_3)
  );
  Element ces_13_0 ( // @[MockArray.scala 36:52]
    .clock(ces_13_0_clock),
    .io_ins_0(ces_13_0_io_ins_0),
    .io_ins_1(ces_13_0_io_ins_1),
    .io_ins_2(ces_13_0_io_ins_2),
    .io_ins_3(ces_13_0_io_ins_3),
    .io_outs_0(ces_13_0_io_outs_0),
    .io_outs_1(ces_13_0_io_outs_1),
    .io_outs_2(ces_13_0_io_outs_2),
    .io_outs_3(ces_13_0_io_outs_3)
  );
  Element ces_13_1 ( // @[MockArray.scala 36:52]
    .clock(ces_13_1_clock),
    .io_ins_0(ces_13_1_io_ins_0),
    .io_ins_1(ces_13_1_io_ins_1),
    .io_ins_2(ces_13_1_io_ins_2),
    .io_ins_3(ces_13_1_io_ins_3),
    .io_outs_0(ces_13_1_io_outs_0),
    .io_outs_1(ces_13_1_io_outs_1),
    .io_outs_2(ces_13_1_io_outs_2),
    .io_outs_3(ces_13_1_io_outs_3)
  );
  Element ces_13_2 ( // @[MockArray.scala 36:52]
    .clock(ces_13_2_clock),
    .io_ins_0(ces_13_2_io_ins_0),
    .io_ins_1(ces_13_2_io_ins_1),
    .io_ins_2(ces_13_2_io_ins_2),
    .io_ins_3(ces_13_2_io_ins_3),
    .io_outs_0(ces_13_2_io_outs_0),
    .io_outs_1(ces_13_2_io_outs_1),
    .io_outs_2(ces_13_2_io_outs_2),
    .io_outs_3(ces_13_2_io_outs_3)
  );
  Element ces_13_3 ( // @[MockArray.scala 36:52]
    .clock(ces_13_3_clock),
    .io_ins_0(ces_13_3_io_ins_0),
    .io_ins_1(ces_13_3_io_ins_1),
    .io_ins_2(ces_13_3_io_ins_2),
    .io_ins_3(ces_13_3_io_ins_3),
    .io_outs_0(ces_13_3_io_outs_0),
    .io_outs_1(ces_13_3_io_outs_1),
    .io_outs_2(ces_13_3_io_outs_2),
    .io_outs_3(ces_13_3_io_outs_3)
  );
  Element ces_13_4 ( // @[MockArray.scala 36:52]
    .clock(ces_13_4_clock),
    .io_ins_0(ces_13_4_io_ins_0),
    .io_ins_1(ces_13_4_io_ins_1),
    .io_ins_2(ces_13_4_io_ins_2),
    .io_ins_3(ces_13_4_io_ins_3),
    .io_outs_0(ces_13_4_io_outs_0),
    .io_outs_1(ces_13_4_io_outs_1),
    .io_outs_2(ces_13_4_io_outs_2),
    .io_outs_3(ces_13_4_io_outs_3)
  );
  Element ces_13_5 ( // @[MockArray.scala 36:52]
    .clock(ces_13_5_clock),
    .io_ins_0(ces_13_5_io_ins_0),
    .io_ins_1(ces_13_5_io_ins_1),
    .io_ins_2(ces_13_5_io_ins_2),
    .io_ins_3(ces_13_5_io_ins_3),
    .io_outs_0(ces_13_5_io_outs_0),
    .io_outs_1(ces_13_5_io_outs_1),
    .io_outs_2(ces_13_5_io_outs_2),
    .io_outs_3(ces_13_5_io_outs_3)
  );
  Element ces_13_6 ( // @[MockArray.scala 36:52]
    .clock(ces_13_6_clock),
    .io_ins_0(ces_13_6_io_ins_0),
    .io_ins_1(ces_13_6_io_ins_1),
    .io_ins_2(ces_13_6_io_ins_2),
    .io_ins_3(ces_13_6_io_ins_3),
    .io_outs_0(ces_13_6_io_outs_0),
    .io_outs_1(ces_13_6_io_outs_1),
    .io_outs_2(ces_13_6_io_outs_2),
    .io_outs_3(ces_13_6_io_outs_3)
  );
  Element ces_13_7 ( // @[MockArray.scala 36:52]
    .clock(ces_13_7_clock),
    .io_ins_0(ces_13_7_io_ins_0),
    .io_ins_1(ces_13_7_io_ins_1),
    .io_ins_2(ces_13_7_io_ins_2),
    .io_ins_3(ces_13_7_io_ins_3),
    .io_outs_0(ces_13_7_io_outs_0),
    .io_outs_1(ces_13_7_io_outs_1),
    .io_outs_2(ces_13_7_io_outs_2),
    .io_outs_3(ces_13_7_io_outs_3)
  );
  Element ces_13_8 ( // @[MockArray.scala 36:52]
    .clock(ces_13_8_clock),
    .io_ins_0(ces_13_8_io_ins_0),
    .io_ins_1(ces_13_8_io_ins_1),
    .io_ins_2(ces_13_8_io_ins_2),
    .io_ins_3(ces_13_8_io_ins_3),
    .io_outs_0(ces_13_8_io_outs_0),
    .io_outs_1(ces_13_8_io_outs_1),
    .io_outs_2(ces_13_8_io_outs_2),
    .io_outs_3(ces_13_8_io_outs_3)
  );
  Element ces_13_9 ( // @[MockArray.scala 36:52]
    .clock(ces_13_9_clock),
    .io_ins_0(ces_13_9_io_ins_0),
    .io_ins_1(ces_13_9_io_ins_1),
    .io_ins_2(ces_13_9_io_ins_2),
    .io_ins_3(ces_13_9_io_ins_3),
    .io_outs_0(ces_13_9_io_outs_0),
    .io_outs_1(ces_13_9_io_outs_1),
    .io_outs_2(ces_13_9_io_outs_2),
    .io_outs_3(ces_13_9_io_outs_3)
  );
  Element ces_13_10 ( // @[MockArray.scala 36:52]
    .clock(ces_13_10_clock),
    .io_ins_0(ces_13_10_io_ins_0),
    .io_ins_1(ces_13_10_io_ins_1),
    .io_ins_2(ces_13_10_io_ins_2),
    .io_ins_3(ces_13_10_io_ins_3),
    .io_outs_0(ces_13_10_io_outs_0),
    .io_outs_1(ces_13_10_io_outs_1),
    .io_outs_2(ces_13_10_io_outs_2),
    .io_outs_3(ces_13_10_io_outs_3)
  );
  Element ces_13_11 ( // @[MockArray.scala 36:52]
    .clock(ces_13_11_clock),
    .io_ins_0(ces_13_11_io_ins_0),
    .io_ins_1(ces_13_11_io_ins_1),
    .io_ins_2(ces_13_11_io_ins_2),
    .io_ins_3(ces_13_11_io_ins_3),
    .io_outs_0(ces_13_11_io_outs_0),
    .io_outs_1(ces_13_11_io_outs_1),
    .io_outs_2(ces_13_11_io_outs_2),
    .io_outs_3(ces_13_11_io_outs_3)
  );
  Element ces_13_12 ( // @[MockArray.scala 36:52]
    .clock(ces_13_12_clock),
    .io_ins_0(ces_13_12_io_ins_0),
    .io_ins_1(ces_13_12_io_ins_1),
    .io_ins_2(ces_13_12_io_ins_2),
    .io_ins_3(ces_13_12_io_ins_3),
    .io_outs_0(ces_13_12_io_outs_0),
    .io_outs_1(ces_13_12_io_outs_1),
    .io_outs_2(ces_13_12_io_outs_2),
    .io_outs_3(ces_13_12_io_outs_3)
  );
  Element ces_13_13 ( // @[MockArray.scala 36:52]
    .clock(ces_13_13_clock),
    .io_ins_0(ces_13_13_io_ins_0),
    .io_ins_1(ces_13_13_io_ins_1),
    .io_ins_2(ces_13_13_io_ins_2),
    .io_ins_3(ces_13_13_io_ins_3),
    .io_outs_0(ces_13_13_io_outs_0),
    .io_outs_1(ces_13_13_io_outs_1),
    .io_outs_2(ces_13_13_io_outs_2),
    .io_outs_3(ces_13_13_io_outs_3)
  );
  Element ces_13_14 ( // @[MockArray.scala 36:52]
    .clock(ces_13_14_clock),
    .io_ins_0(ces_13_14_io_ins_0),
    .io_ins_1(ces_13_14_io_ins_1),
    .io_ins_2(ces_13_14_io_ins_2),
    .io_ins_3(ces_13_14_io_ins_3),
    .io_outs_0(ces_13_14_io_outs_0),
    .io_outs_1(ces_13_14_io_outs_1),
    .io_outs_2(ces_13_14_io_outs_2),
    .io_outs_3(ces_13_14_io_outs_3)
  );
  Element ces_13_15 ( // @[MockArray.scala 36:52]
    .clock(ces_13_15_clock),
    .io_ins_0(ces_13_15_io_ins_0),
    .io_ins_1(ces_13_15_io_ins_1),
    .io_ins_2(ces_13_15_io_ins_2),
    .io_ins_3(ces_13_15_io_ins_3),
    .io_outs_0(ces_13_15_io_outs_0),
    .io_outs_1(ces_13_15_io_outs_1),
    .io_outs_2(ces_13_15_io_outs_2),
    .io_outs_3(ces_13_15_io_outs_3)
  );
  Element ces_13_16 ( // @[MockArray.scala 36:52]
    .clock(ces_13_16_clock),
    .io_ins_0(ces_13_16_io_ins_0),
    .io_ins_1(ces_13_16_io_ins_1),
    .io_ins_2(ces_13_16_io_ins_2),
    .io_ins_3(ces_13_16_io_ins_3),
    .io_outs_0(ces_13_16_io_outs_0),
    .io_outs_1(ces_13_16_io_outs_1),
    .io_outs_2(ces_13_16_io_outs_2),
    .io_outs_3(ces_13_16_io_outs_3)
  );
  Element ces_13_17 ( // @[MockArray.scala 36:52]
    .clock(ces_13_17_clock),
    .io_ins_0(ces_13_17_io_ins_0),
    .io_ins_1(ces_13_17_io_ins_1),
    .io_ins_2(ces_13_17_io_ins_2),
    .io_ins_3(ces_13_17_io_ins_3),
    .io_outs_0(ces_13_17_io_outs_0),
    .io_outs_1(ces_13_17_io_outs_1),
    .io_outs_2(ces_13_17_io_outs_2),
    .io_outs_3(ces_13_17_io_outs_3)
  );
  Element ces_13_18 ( // @[MockArray.scala 36:52]
    .clock(ces_13_18_clock),
    .io_ins_0(ces_13_18_io_ins_0),
    .io_ins_1(ces_13_18_io_ins_1),
    .io_ins_2(ces_13_18_io_ins_2),
    .io_ins_3(ces_13_18_io_ins_3),
    .io_outs_0(ces_13_18_io_outs_0),
    .io_outs_1(ces_13_18_io_outs_1),
    .io_outs_2(ces_13_18_io_outs_2),
    .io_outs_3(ces_13_18_io_outs_3)
  );
  Element ces_13_19 ( // @[MockArray.scala 36:52]
    .clock(ces_13_19_clock),
    .io_ins_0(ces_13_19_io_ins_0),
    .io_ins_1(ces_13_19_io_ins_1),
    .io_ins_2(ces_13_19_io_ins_2),
    .io_ins_3(ces_13_19_io_ins_3),
    .io_outs_0(ces_13_19_io_outs_0),
    .io_outs_1(ces_13_19_io_outs_1),
    .io_outs_2(ces_13_19_io_outs_2),
    .io_outs_3(ces_13_19_io_outs_3)
  );
  Element ces_13_20 ( // @[MockArray.scala 36:52]
    .clock(ces_13_20_clock),
    .io_ins_0(ces_13_20_io_ins_0),
    .io_ins_1(ces_13_20_io_ins_1),
    .io_ins_2(ces_13_20_io_ins_2),
    .io_ins_3(ces_13_20_io_ins_3),
    .io_outs_0(ces_13_20_io_outs_0),
    .io_outs_1(ces_13_20_io_outs_1),
    .io_outs_2(ces_13_20_io_outs_2),
    .io_outs_3(ces_13_20_io_outs_3)
  );
  Element ces_13_21 ( // @[MockArray.scala 36:52]
    .clock(ces_13_21_clock),
    .io_ins_0(ces_13_21_io_ins_0),
    .io_ins_1(ces_13_21_io_ins_1),
    .io_ins_2(ces_13_21_io_ins_2),
    .io_ins_3(ces_13_21_io_ins_3),
    .io_outs_0(ces_13_21_io_outs_0),
    .io_outs_1(ces_13_21_io_outs_1),
    .io_outs_2(ces_13_21_io_outs_2),
    .io_outs_3(ces_13_21_io_outs_3)
  );
  Element ces_13_22 ( // @[MockArray.scala 36:52]
    .clock(ces_13_22_clock),
    .io_ins_0(ces_13_22_io_ins_0),
    .io_ins_1(ces_13_22_io_ins_1),
    .io_ins_2(ces_13_22_io_ins_2),
    .io_ins_3(ces_13_22_io_ins_3),
    .io_outs_0(ces_13_22_io_outs_0),
    .io_outs_1(ces_13_22_io_outs_1),
    .io_outs_2(ces_13_22_io_outs_2),
    .io_outs_3(ces_13_22_io_outs_3)
  );
  Element ces_13_23 ( // @[MockArray.scala 36:52]
    .clock(ces_13_23_clock),
    .io_ins_0(ces_13_23_io_ins_0),
    .io_ins_1(ces_13_23_io_ins_1),
    .io_ins_2(ces_13_23_io_ins_2),
    .io_ins_3(ces_13_23_io_ins_3),
    .io_outs_0(ces_13_23_io_outs_0),
    .io_outs_1(ces_13_23_io_outs_1),
    .io_outs_2(ces_13_23_io_outs_2),
    .io_outs_3(ces_13_23_io_outs_3)
  );
  Element ces_13_24 ( // @[MockArray.scala 36:52]
    .clock(ces_13_24_clock),
    .io_ins_0(ces_13_24_io_ins_0),
    .io_ins_1(ces_13_24_io_ins_1),
    .io_ins_2(ces_13_24_io_ins_2),
    .io_ins_3(ces_13_24_io_ins_3),
    .io_outs_0(ces_13_24_io_outs_0),
    .io_outs_1(ces_13_24_io_outs_1),
    .io_outs_2(ces_13_24_io_outs_2),
    .io_outs_3(ces_13_24_io_outs_3)
  );
  Element ces_13_25 ( // @[MockArray.scala 36:52]
    .clock(ces_13_25_clock),
    .io_ins_0(ces_13_25_io_ins_0),
    .io_ins_1(ces_13_25_io_ins_1),
    .io_ins_2(ces_13_25_io_ins_2),
    .io_ins_3(ces_13_25_io_ins_3),
    .io_outs_0(ces_13_25_io_outs_0),
    .io_outs_1(ces_13_25_io_outs_1),
    .io_outs_2(ces_13_25_io_outs_2),
    .io_outs_3(ces_13_25_io_outs_3)
  );
  Element ces_13_26 ( // @[MockArray.scala 36:52]
    .clock(ces_13_26_clock),
    .io_ins_0(ces_13_26_io_ins_0),
    .io_ins_1(ces_13_26_io_ins_1),
    .io_ins_2(ces_13_26_io_ins_2),
    .io_ins_3(ces_13_26_io_ins_3),
    .io_outs_0(ces_13_26_io_outs_0),
    .io_outs_1(ces_13_26_io_outs_1),
    .io_outs_2(ces_13_26_io_outs_2),
    .io_outs_3(ces_13_26_io_outs_3)
  );
  Element ces_13_27 ( // @[MockArray.scala 36:52]
    .clock(ces_13_27_clock),
    .io_ins_0(ces_13_27_io_ins_0),
    .io_ins_1(ces_13_27_io_ins_1),
    .io_ins_2(ces_13_27_io_ins_2),
    .io_ins_3(ces_13_27_io_ins_3),
    .io_outs_0(ces_13_27_io_outs_0),
    .io_outs_1(ces_13_27_io_outs_1),
    .io_outs_2(ces_13_27_io_outs_2),
    .io_outs_3(ces_13_27_io_outs_3)
  );
  Element ces_13_28 ( // @[MockArray.scala 36:52]
    .clock(ces_13_28_clock),
    .io_ins_0(ces_13_28_io_ins_0),
    .io_ins_1(ces_13_28_io_ins_1),
    .io_ins_2(ces_13_28_io_ins_2),
    .io_ins_3(ces_13_28_io_ins_3),
    .io_outs_0(ces_13_28_io_outs_0),
    .io_outs_1(ces_13_28_io_outs_1),
    .io_outs_2(ces_13_28_io_outs_2),
    .io_outs_3(ces_13_28_io_outs_3)
  );
  Element ces_13_29 ( // @[MockArray.scala 36:52]
    .clock(ces_13_29_clock),
    .io_ins_0(ces_13_29_io_ins_0),
    .io_ins_1(ces_13_29_io_ins_1),
    .io_ins_2(ces_13_29_io_ins_2),
    .io_ins_3(ces_13_29_io_ins_3),
    .io_outs_0(ces_13_29_io_outs_0),
    .io_outs_1(ces_13_29_io_outs_1),
    .io_outs_2(ces_13_29_io_outs_2),
    .io_outs_3(ces_13_29_io_outs_3)
  );
  Element ces_13_30 ( // @[MockArray.scala 36:52]
    .clock(ces_13_30_clock),
    .io_ins_0(ces_13_30_io_ins_0),
    .io_ins_1(ces_13_30_io_ins_1),
    .io_ins_2(ces_13_30_io_ins_2),
    .io_ins_3(ces_13_30_io_ins_3),
    .io_outs_0(ces_13_30_io_outs_0),
    .io_outs_1(ces_13_30_io_outs_1),
    .io_outs_2(ces_13_30_io_outs_2),
    .io_outs_3(ces_13_30_io_outs_3)
  );
  Element ces_13_31 ( // @[MockArray.scala 36:52]
    .clock(ces_13_31_clock),
    .io_ins_0(ces_13_31_io_ins_0),
    .io_ins_1(ces_13_31_io_ins_1),
    .io_ins_2(ces_13_31_io_ins_2),
    .io_ins_3(ces_13_31_io_ins_3),
    .io_outs_0(ces_13_31_io_outs_0),
    .io_outs_1(ces_13_31_io_outs_1),
    .io_outs_2(ces_13_31_io_outs_2),
    .io_outs_3(ces_13_31_io_outs_3)
  );
  Element ces_14_0 ( // @[MockArray.scala 36:52]
    .clock(ces_14_0_clock),
    .io_ins_0(ces_14_0_io_ins_0),
    .io_ins_1(ces_14_0_io_ins_1),
    .io_ins_2(ces_14_0_io_ins_2),
    .io_ins_3(ces_14_0_io_ins_3),
    .io_outs_0(ces_14_0_io_outs_0),
    .io_outs_1(ces_14_0_io_outs_1),
    .io_outs_2(ces_14_0_io_outs_2),
    .io_outs_3(ces_14_0_io_outs_3)
  );
  Element ces_14_1 ( // @[MockArray.scala 36:52]
    .clock(ces_14_1_clock),
    .io_ins_0(ces_14_1_io_ins_0),
    .io_ins_1(ces_14_1_io_ins_1),
    .io_ins_2(ces_14_1_io_ins_2),
    .io_ins_3(ces_14_1_io_ins_3),
    .io_outs_0(ces_14_1_io_outs_0),
    .io_outs_1(ces_14_1_io_outs_1),
    .io_outs_2(ces_14_1_io_outs_2),
    .io_outs_3(ces_14_1_io_outs_3)
  );
  Element ces_14_2 ( // @[MockArray.scala 36:52]
    .clock(ces_14_2_clock),
    .io_ins_0(ces_14_2_io_ins_0),
    .io_ins_1(ces_14_2_io_ins_1),
    .io_ins_2(ces_14_2_io_ins_2),
    .io_ins_3(ces_14_2_io_ins_3),
    .io_outs_0(ces_14_2_io_outs_0),
    .io_outs_1(ces_14_2_io_outs_1),
    .io_outs_2(ces_14_2_io_outs_2),
    .io_outs_3(ces_14_2_io_outs_3)
  );
  Element ces_14_3 ( // @[MockArray.scala 36:52]
    .clock(ces_14_3_clock),
    .io_ins_0(ces_14_3_io_ins_0),
    .io_ins_1(ces_14_3_io_ins_1),
    .io_ins_2(ces_14_3_io_ins_2),
    .io_ins_3(ces_14_3_io_ins_3),
    .io_outs_0(ces_14_3_io_outs_0),
    .io_outs_1(ces_14_3_io_outs_1),
    .io_outs_2(ces_14_3_io_outs_2),
    .io_outs_3(ces_14_3_io_outs_3)
  );
  Element ces_14_4 ( // @[MockArray.scala 36:52]
    .clock(ces_14_4_clock),
    .io_ins_0(ces_14_4_io_ins_0),
    .io_ins_1(ces_14_4_io_ins_1),
    .io_ins_2(ces_14_4_io_ins_2),
    .io_ins_3(ces_14_4_io_ins_3),
    .io_outs_0(ces_14_4_io_outs_0),
    .io_outs_1(ces_14_4_io_outs_1),
    .io_outs_2(ces_14_4_io_outs_2),
    .io_outs_3(ces_14_4_io_outs_3)
  );
  Element ces_14_5 ( // @[MockArray.scala 36:52]
    .clock(ces_14_5_clock),
    .io_ins_0(ces_14_5_io_ins_0),
    .io_ins_1(ces_14_5_io_ins_1),
    .io_ins_2(ces_14_5_io_ins_2),
    .io_ins_3(ces_14_5_io_ins_3),
    .io_outs_0(ces_14_5_io_outs_0),
    .io_outs_1(ces_14_5_io_outs_1),
    .io_outs_2(ces_14_5_io_outs_2),
    .io_outs_3(ces_14_5_io_outs_3)
  );
  Element ces_14_6 ( // @[MockArray.scala 36:52]
    .clock(ces_14_6_clock),
    .io_ins_0(ces_14_6_io_ins_0),
    .io_ins_1(ces_14_6_io_ins_1),
    .io_ins_2(ces_14_6_io_ins_2),
    .io_ins_3(ces_14_6_io_ins_3),
    .io_outs_0(ces_14_6_io_outs_0),
    .io_outs_1(ces_14_6_io_outs_1),
    .io_outs_2(ces_14_6_io_outs_2),
    .io_outs_3(ces_14_6_io_outs_3)
  );
  Element ces_14_7 ( // @[MockArray.scala 36:52]
    .clock(ces_14_7_clock),
    .io_ins_0(ces_14_7_io_ins_0),
    .io_ins_1(ces_14_7_io_ins_1),
    .io_ins_2(ces_14_7_io_ins_2),
    .io_ins_3(ces_14_7_io_ins_3),
    .io_outs_0(ces_14_7_io_outs_0),
    .io_outs_1(ces_14_7_io_outs_1),
    .io_outs_2(ces_14_7_io_outs_2),
    .io_outs_3(ces_14_7_io_outs_3)
  );
  Element ces_14_8 ( // @[MockArray.scala 36:52]
    .clock(ces_14_8_clock),
    .io_ins_0(ces_14_8_io_ins_0),
    .io_ins_1(ces_14_8_io_ins_1),
    .io_ins_2(ces_14_8_io_ins_2),
    .io_ins_3(ces_14_8_io_ins_3),
    .io_outs_0(ces_14_8_io_outs_0),
    .io_outs_1(ces_14_8_io_outs_1),
    .io_outs_2(ces_14_8_io_outs_2),
    .io_outs_3(ces_14_8_io_outs_3)
  );
  Element ces_14_9 ( // @[MockArray.scala 36:52]
    .clock(ces_14_9_clock),
    .io_ins_0(ces_14_9_io_ins_0),
    .io_ins_1(ces_14_9_io_ins_1),
    .io_ins_2(ces_14_9_io_ins_2),
    .io_ins_3(ces_14_9_io_ins_3),
    .io_outs_0(ces_14_9_io_outs_0),
    .io_outs_1(ces_14_9_io_outs_1),
    .io_outs_2(ces_14_9_io_outs_2),
    .io_outs_3(ces_14_9_io_outs_3)
  );
  Element ces_14_10 ( // @[MockArray.scala 36:52]
    .clock(ces_14_10_clock),
    .io_ins_0(ces_14_10_io_ins_0),
    .io_ins_1(ces_14_10_io_ins_1),
    .io_ins_2(ces_14_10_io_ins_2),
    .io_ins_3(ces_14_10_io_ins_3),
    .io_outs_0(ces_14_10_io_outs_0),
    .io_outs_1(ces_14_10_io_outs_1),
    .io_outs_2(ces_14_10_io_outs_2),
    .io_outs_3(ces_14_10_io_outs_3)
  );
  Element ces_14_11 ( // @[MockArray.scala 36:52]
    .clock(ces_14_11_clock),
    .io_ins_0(ces_14_11_io_ins_0),
    .io_ins_1(ces_14_11_io_ins_1),
    .io_ins_2(ces_14_11_io_ins_2),
    .io_ins_3(ces_14_11_io_ins_3),
    .io_outs_0(ces_14_11_io_outs_0),
    .io_outs_1(ces_14_11_io_outs_1),
    .io_outs_2(ces_14_11_io_outs_2),
    .io_outs_3(ces_14_11_io_outs_3)
  );
  Element ces_14_12 ( // @[MockArray.scala 36:52]
    .clock(ces_14_12_clock),
    .io_ins_0(ces_14_12_io_ins_0),
    .io_ins_1(ces_14_12_io_ins_1),
    .io_ins_2(ces_14_12_io_ins_2),
    .io_ins_3(ces_14_12_io_ins_3),
    .io_outs_0(ces_14_12_io_outs_0),
    .io_outs_1(ces_14_12_io_outs_1),
    .io_outs_2(ces_14_12_io_outs_2),
    .io_outs_3(ces_14_12_io_outs_3)
  );
  Element ces_14_13 ( // @[MockArray.scala 36:52]
    .clock(ces_14_13_clock),
    .io_ins_0(ces_14_13_io_ins_0),
    .io_ins_1(ces_14_13_io_ins_1),
    .io_ins_2(ces_14_13_io_ins_2),
    .io_ins_3(ces_14_13_io_ins_3),
    .io_outs_0(ces_14_13_io_outs_0),
    .io_outs_1(ces_14_13_io_outs_1),
    .io_outs_2(ces_14_13_io_outs_2),
    .io_outs_3(ces_14_13_io_outs_3)
  );
  Element ces_14_14 ( // @[MockArray.scala 36:52]
    .clock(ces_14_14_clock),
    .io_ins_0(ces_14_14_io_ins_0),
    .io_ins_1(ces_14_14_io_ins_1),
    .io_ins_2(ces_14_14_io_ins_2),
    .io_ins_3(ces_14_14_io_ins_3),
    .io_outs_0(ces_14_14_io_outs_0),
    .io_outs_1(ces_14_14_io_outs_1),
    .io_outs_2(ces_14_14_io_outs_2),
    .io_outs_3(ces_14_14_io_outs_3)
  );
  Element ces_14_15 ( // @[MockArray.scala 36:52]
    .clock(ces_14_15_clock),
    .io_ins_0(ces_14_15_io_ins_0),
    .io_ins_1(ces_14_15_io_ins_1),
    .io_ins_2(ces_14_15_io_ins_2),
    .io_ins_3(ces_14_15_io_ins_3),
    .io_outs_0(ces_14_15_io_outs_0),
    .io_outs_1(ces_14_15_io_outs_1),
    .io_outs_2(ces_14_15_io_outs_2),
    .io_outs_3(ces_14_15_io_outs_3)
  );
  Element ces_14_16 ( // @[MockArray.scala 36:52]
    .clock(ces_14_16_clock),
    .io_ins_0(ces_14_16_io_ins_0),
    .io_ins_1(ces_14_16_io_ins_1),
    .io_ins_2(ces_14_16_io_ins_2),
    .io_ins_3(ces_14_16_io_ins_3),
    .io_outs_0(ces_14_16_io_outs_0),
    .io_outs_1(ces_14_16_io_outs_1),
    .io_outs_2(ces_14_16_io_outs_2),
    .io_outs_3(ces_14_16_io_outs_3)
  );
  Element ces_14_17 ( // @[MockArray.scala 36:52]
    .clock(ces_14_17_clock),
    .io_ins_0(ces_14_17_io_ins_0),
    .io_ins_1(ces_14_17_io_ins_1),
    .io_ins_2(ces_14_17_io_ins_2),
    .io_ins_3(ces_14_17_io_ins_3),
    .io_outs_0(ces_14_17_io_outs_0),
    .io_outs_1(ces_14_17_io_outs_1),
    .io_outs_2(ces_14_17_io_outs_2),
    .io_outs_3(ces_14_17_io_outs_3)
  );
  Element ces_14_18 ( // @[MockArray.scala 36:52]
    .clock(ces_14_18_clock),
    .io_ins_0(ces_14_18_io_ins_0),
    .io_ins_1(ces_14_18_io_ins_1),
    .io_ins_2(ces_14_18_io_ins_2),
    .io_ins_3(ces_14_18_io_ins_3),
    .io_outs_0(ces_14_18_io_outs_0),
    .io_outs_1(ces_14_18_io_outs_1),
    .io_outs_2(ces_14_18_io_outs_2),
    .io_outs_3(ces_14_18_io_outs_3)
  );
  Element ces_14_19 ( // @[MockArray.scala 36:52]
    .clock(ces_14_19_clock),
    .io_ins_0(ces_14_19_io_ins_0),
    .io_ins_1(ces_14_19_io_ins_1),
    .io_ins_2(ces_14_19_io_ins_2),
    .io_ins_3(ces_14_19_io_ins_3),
    .io_outs_0(ces_14_19_io_outs_0),
    .io_outs_1(ces_14_19_io_outs_1),
    .io_outs_2(ces_14_19_io_outs_2),
    .io_outs_3(ces_14_19_io_outs_3)
  );
  Element ces_14_20 ( // @[MockArray.scala 36:52]
    .clock(ces_14_20_clock),
    .io_ins_0(ces_14_20_io_ins_0),
    .io_ins_1(ces_14_20_io_ins_1),
    .io_ins_2(ces_14_20_io_ins_2),
    .io_ins_3(ces_14_20_io_ins_3),
    .io_outs_0(ces_14_20_io_outs_0),
    .io_outs_1(ces_14_20_io_outs_1),
    .io_outs_2(ces_14_20_io_outs_2),
    .io_outs_3(ces_14_20_io_outs_3)
  );
  Element ces_14_21 ( // @[MockArray.scala 36:52]
    .clock(ces_14_21_clock),
    .io_ins_0(ces_14_21_io_ins_0),
    .io_ins_1(ces_14_21_io_ins_1),
    .io_ins_2(ces_14_21_io_ins_2),
    .io_ins_3(ces_14_21_io_ins_3),
    .io_outs_0(ces_14_21_io_outs_0),
    .io_outs_1(ces_14_21_io_outs_1),
    .io_outs_2(ces_14_21_io_outs_2),
    .io_outs_3(ces_14_21_io_outs_3)
  );
  Element ces_14_22 ( // @[MockArray.scala 36:52]
    .clock(ces_14_22_clock),
    .io_ins_0(ces_14_22_io_ins_0),
    .io_ins_1(ces_14_22_io_ins_1),
    .io_ins_2(ces_14_22_io_ins_2),
    .io_ins_3(ces_14_22_io_ins_3),
    .io_outs_0(ces_14_22_io_outs_0),
    .io_outs_1(ces_14_22_io_outs_1),
    .io_outs_2(ces_14_22_io_outs_2),
    .io_outs_3(ces_14_22_io_outs_3)
  );
  Element ces_14_23 ( // @[MockArray.scala 36:52]
    .clock(ces_14_23_clock),
    .io_ins_0(ces_14_23_io_ins_0),
    .io_ins_1(ces_14_23_io_ins_1),
    .io_ins_2(ces_14_23_io_ins_2),
    .io_ins_3(ces_14_23_io_ins_3),
    .io_outs_0(ces_14_23_io_outs_0),
    .io_outs_1(ces_14_23_io_outs_1),
    .io_outs_2(ces_14_23_io_outs_2),
    .io_outs_3(ces_14_23_io_outs_3)
  );
  Element ces_14_24 ( // @[MockArray.scala 36:52]
    .clock(ces_14_24_clock),
    .io_ins_0(ces_14_24_io_ins_0),
    .io_ins_1(ces_14_24_io_ins_1),
    .io_ins_2(ces_14_24_io_ins_2),
    .io_ins_3(ces_14_24_io_ins_3),
    .io_outs_0(ces_14_24_io_outs_0),
    .io_outs_1(ces_14_24_io_outs_1),
    .io_outs_2(ces_14_24_io_outs_2),
    .io_outs_3(ces_14_24_io_outs_3)
  );
  Element ces_14_25 ( // @[MockArray.scala 36:52]
    .clock(ces_14_25_clock),
    .io_ins_0(ces_14_25_io_ins_0),
    .io_ins_1(ces_14_25_io_ins_1),
    .io_ins_2(ces_14_25_io_ins_2),
    .io_ins_3(ces_14_25_io_ins_3),
    .io_outs_0(ces_14_25_io_outs_0),
    .io_outs_1(ces_14_25_io_outs_1),
    .io_outs_2(ces_14_25_io_outs_2),
    .io_outs_3(ces_14_25_io_outs_3)
  );
  Element ces_14_26 ( // @[MockArray.scala 36:52]
    .clock(ces_14_26_clock),
    .io_ins_0(ces_14_26_io_ins_0),
    .io_ins_1(ces_14_26_io_ins_1),
    .io_ins_2(ces_14_26_io_ins_2),
    .io_ins_3(ces_14_26_io_ins_3),
    .io_outs_0(ces_14_26_io_outs_0),
    .io_outs_1(ces_14_26_io_outs_1),
    .io_outs_2(ces_14_26_io_outs_2),
    .io_outs_3(ces_14_26_io_outs_3)
  );
  Element ces_14_27 ( // @[MockArray.scala 36:52]
    .clock(ces_14_27_clock),
    .io_ins_0(ces_14_27_io_ins_0),
    .io_ins_1(ces_14_27_io_ins_1),
    .io_ins_2(ces_14_27_io_ins_2),
    .io_ins_3(ces_14_27_io_ins_3),
    .io_outs_0(ces_14_27_io_outs_0),
    .io_outs_1(ces_14_27_io_outs_1),
    .io_outs_2(ces_14_27_io_outs_2),
    .io_outs_3(ces_14_27_io_outs_3)
  );
  Element ces_14_28 ( // @[MockArray.scala 36:52]
    .clock(ces_14_28_clock),
    .io_ins_0(ces_14_28_io_ins_0),
    .io_ins_1(ces_14_28_io_ins_1),
    .io_ins_2(ces_14_28_io_ins_2),
    .io_ins_3(ces_14_28_io_ins_3),
    .io_outs_0(ces_14_28_io_outs_0),
    .io_outs_1(ces_14_28_io_outs_1),
    .io_outs_2(ces_14_28_io_outs_2),
    .io_outs_3(ces_14_28_io_outs_3)
  );
  Element ces_14_29 ( // @[MockArray.scala 36:52]
    .clock(ces_14_29_clock),
    .io_ins_0(ces_14_29_io_ins_0),
    .io_ins_1(ces_14_29_io_ins_1),
    .io_ins_2(ces_14_29_io_ins_2),
    .io_ins_3(ces_14_29_io_ins_3),
    .io_outs_0(ces_14_29_io_outs_0),
    .io_outs_1(ces_14_29_io_outs_1),
    .io_outs_2(ces_14_29_io_outs_2),
    .io_outs_3(ces_14_29_io_outs_3)
  );
  Element ces_14_30 ( // @[MockArray.scala 36:52]
    .clock(ces_14_30_clock),
    .io_ins_0(ces_14_30_io_ins_0),
    .io_ins_1(ces_14_30_io_ins_1),
    .io_ins_2(ces_14_30_io_ins_2),
    .io_ins_3(ces_14_30_io_ins_3),
    .io_outs_0(ces_14_30_io_outs_0),
    .io_outs_1(ces_14_30_io_outs_1),
    .io_outs_2(ces_14_30_io_outs_2),
    .io_outs_3(ces_14_30_io_outs_3)
  );
  Element ces_14_31 ( // @[MockArray.scala 36:52]
    .clock(ces_14_31_clock),
    .io_ins_0(ces_14_31_io_ins_0),
    .io_ins_1(ces_14_31_io_ins_1),
    .io_ins_2(ces_14_31_io_ins_2),
    .io_ins_3(ces_14_31_io_ins_3),
    .io_outs_0(ces_14_31_io_outs_0),
    .io_outs_1(ces_14_31_io_outs_1),
    .io_outs_2(ces_14_31_io_outs_2),
    .io_outs_3(ces_14_31_io_outs_3)
  );
  Element ces_15_0 ( // @[MockArray.scala 36:52]
    .clock(ces_15_0_clock),
    .io_ins_0(ces_15_0_io_ins_0),
    .io_ins_1(ces_15_0_io_ins_1),
    .io_ins_2(ces_15_0_io_ins_2),
    .io_ins_3(ces_15_0_io_ins_3),
    .io_outs_0(ces_15_0_io_outs_0),
    .io_outs_1(ces_15_0_io_outs_1),
    .io_outs_2(ces_15_0_io_outs_2),
    .io_outs_3(ces_15_0_io_outs_3)
  );
  Element ces_15_1 ( // @[MockArray.scala 36:52]
    .clock(ces_15_1_clock),
    .io_ins_0(ces_15_1_io_ins_0),
    .io_ins_1(ces_15_1_io_ins_1),
    .io_ins_2(ces_15_1_io_ins_2),
    .io_ins_3(ces_15_1_io_ins_3),
    .io_outs_0(ces_15_1_io_outs_0),
    .io_outs_1(ces_15_1_io_outs_1),
    .io_outs_2(ces_15_1_io_outs_2),
    .io_outs_3(ces_15_1_io_outs_3)
  );
  Element ces_15_2 ( // @[MockArray.scala 36:52]
    .clock(ces_15_2_clock),
    .io_ins_0(ces_15_2_io_ins_0),
    .io_ins_1(ces_15_2_io_ins_1),
    .io_ins_2(ces_15_2_io_ins_2),
    .io_ins_3(ces_15_2_io_ins_3),
    .io_outs_0(ces_15_2_io_outs_0),
    .io_outs_1(ces_15_2_io_outs_1),
    .io_outs_2(ces_15_2_io_outs_2),
    .io_outs_3(ces_15_2_io_outs_3)
  );
  Element ces_15_3 ( // @[MockArray.scala 36:52]
    .clock(ces_15_3_clock),
    .io_ins_0(ces_15_3_io_ins_0),
    .io_ins_1(ces_15_3_io_ins_1),
    .io_ins_2(ces_15_3_io_ins_2),
    .io_ins_3(ces_15_3_io_ins_3),
    .io_outs_0(ces_15_3_io_outs_0),
    .io_outs_1(ces_15_3_io_outs_1),
    .io_outs_2(ces_15_3_io_outs_2),
    .io_outs_3(ces_15_3_io_outs_3)
  );
  Element ces_15_4 ( // @[MockArray.scala 36:52]
    .clock(ces_15_4_clock),
    .io_ins_0(ces_15_4_io_ins_0),
    .io_ins_1(ces_15_4_io_ins_1),
    .io_ins_2(ces_15_4_io_ins_2),
    .io_ins_3(ces_15_4_io_ins_3),
    .io_outs_0(ces_15_4_io_outs_0),
    .io_outs_1(ces_15_4_io_outs_1),
    .io_outs_2(ces_15_4_io_outs_2),
    .io_outs_3(ces_15_4_io_outs_3)
  );
  Element ces_15_5 ( // @[MockArray.scala 36:52]
    .clock(ces_15_5_clock),
    .io_ins_0(ces_15_5_io_ins_0),
    .io_ins_1(ces_15_5_io_ins_1),
    .io_ins_2(ces_15_5_io_ins_2),
    .io_ins_3(ces_15_5_io_ins_3),
    .io_outs_0(ces_15_5_io_outs_0),
    .io_outs_1(ces_15_5_io_outs_1),
    .io_outs_2(ces_15_5_io_outs_2),
    .io_outs_3(ces_15_5_io_outs_3)
  );
  Element ces_15_6 ( // @[MockArray.scala 36:52]
    .clock(ces_15_6_clock),
    .io_ins_0(ces_15_6_io_ins_0),
    .io_ins_1(ces_15_6_io_ins_1),
    .io_ins_2(ces_15_6_io_ins_2),
    .io_ins_3(ces_15_6_io_ins_3),
    .io_outs_0(ces_15_6_io_outs_0),
    .io_outs_1(ces_15_6_io_outs_1),
    .io_outs_2(ces_15_6_io_outs_2),
    .io_outs_3(ces_15_6_io_outs_3)
  );
  Element ces_15_7 ( // @[MockArray.scala 36:52]
    .clock(ces_15_7_clock),
    .io_ins_0(ces_15_7_io_ins_0),
    .io_ins_1(ces_15_7_io_ins_1),
    .io_ins_2(ces_15_7_io_ins_2),
    .io_ins_3(ces_15_7_io_ins_3),
    .io_outs_0(ces_15_7_io_outs_0),
    .io_outs_1(ces_15_7_io_outs_1),
    .io_outs_2(ces_15_7_io_outs_2),
    .io_outs_3(ces_15_7_io_outs_3)
  );
  Element ces_15_8 ( // @[MockArray.scala 36:52]
    .clock(ces_15_8_clock),
    .io_ins_0(ces_15_8_io_ins_0),
    .io_ins_1(ces_15_8_io_ins_1),
    .io_ins_2(ces_15_8_io_ins_2),
    .io_ins_3(ces_15_8_io_ins_3),
    .io_outs_0(ces_15_8_io_outs_0),
    .io_outs_1(ces_15_8_io_outs_1),
    .io_outs_2(ces_15_8_io_outs_2),
    .io_outs_3(ces_15_8_io_outs_3)
  );
  Element ces_15_9 ( // @[MockArray.scala 36:52]
    .clock(ces_15_9_clock),
    .io_ins_0(ces_15_9_io_ins_0),
    .io_ins_1(ces_15_9_io_ins_1),
    .io_ins_2(ces_15_9_io_ins_2),
    .io_ins_3(ces_15_9_io_ins_3),
    .io_outs_0(ces_15_9_io_outs_0),
    .io_outs_1(ces_15_9_io_outs_1),
    .io_outs_2(ces_15_9_io_outs_2),
    .io_outs_3(ces_15_9_io_outs_3)
  );
  Element ces_15_10 ( // @[MockArray.scala 36:52]
    .clock(ces_15_10_clock),
    .io_ins_0(ces_15_10_io_ins_0),
    .io_ins_1(ces_15_10_io_ins_1),
    .io_ins_2(ces_15_10_io_ins_2),
    .io_ins_3(ces_15_10_io_ins_3),
    .io_outs_0(ces_15_10_io_outs_0),
    .io_outs_1(ces_15_10_io_outs_1),
    .io_outs_2(ces_15_10_io_outs_2),
    .io_outs_3(ces_15_10_io_outs_3)
  );
  Element ces_15_11 ( // @[MockArray.scala 36:52]
    .clock(ces_15_11_clock),
    .io_ins_0(ces_15_11_io_ins_0),
    .io_ins_1(ces_15_11_io_ins_1),
    .io_ins_2(ces_15_11_io_ins_2),
    .io_ins_3(ces_15_11_io_ins_3),
    .io_outs_0(ces_15_11_io_outs_0),
    .io_outs_1(ces_15_11_io_outs_1),
    .io_outs_2(ces_15_11_io_outs_2),
    .io_outs_3(ces_15_11_io_outs_3)
  );
  Element ces_15_12 ( // @[MockArray.scala 36:52]
    .clock(ces_15_12_clock),
    .io_ins_0(ces_15_12_io_ins_0),
    .io_ins_1(ces_15_12_io_ins_1),
    .io_ins_2(ces_15_12_io_ins_2),
    .io_ins_3(ces_15_12_io_ins_3),
    .io_outs_0(ces_15_12_io_outs_0),
    .io_outs_1(ces_15_12_io_outs_1),
    .io_outs_2(ces_15_12_io_outs_2),
    .io_outs_3(ces_15_12_io_outs_3)
  );
  Element ces_15_13 ( // @[MockArray.scala 36:52]
    .clock(ces_15_13_clock),
    .io_ins_0(ces_15_13_io_ins_0),
    .io_ins_1(ces_15_13_io_ins_1),
    .io_ins_2(ces_15_13_io_ins_2),
    .io_ins_3(ces_15_13_io_ins_3),
    .io_outs_0(ces_15_13_io_outs_0),
    .io_outs_1(ces_15_13_io_outs_1),
    .io_outs_2(ces_15_13_io_outs_2),
    .io_outs_3(ces_15_13_io_outs_3)
  );
  Element ces_15_14 ( // @[MockArray.scala 36:52]
    .clock(ces_15_14_clock),
    .io_ins_0(ces_15_14_io_ins_0),
    .io_ins_1(ces_15_14_io_ins_1),
    .io_ins_2(ces_15_14_io_ins_2),
    .io_ins_3(ces_15_14_io_ins_3),
    .io_outs_0(ces_15_14_io_outs_0),
    .io_outs_1(ces_15_14_io_outs_1),
    .io_outs_2(ces_15_14_io_outs_2),
    .io_outs_3(ces_15_14_io_outs_3)
  );
  Element ces_15_15 ( // @[MockArray.scala 36:52]
    .clock(ces_15_15_clock),
    .io_ins_0(ces_15_15_io_ins_0),
    .io_ins_1(ces_15_15_io_ins_1),
    .io_ins_2(ces_15_15_io_ins_2),
    .io_ins_3(ces_15_15_io_ins_3),
    .io_outs_0(ces_15_15_io_outs_0),
    .io_outs_1(ces_15_15_io_outs_1),
    .io_outs_2(ces_15_15_io_outs_2),
    .io_outs_3(ces_15_15_io_outs_3)
  );
  Element ces_15_16 ( // @[MockArray.scala 36:52]
    .clock(ces_15_16_clock),
    .io_ins_0(ces_15_16_io_ins_0),
    .io_ins_1(ces_15_16_io_ins_1),
    .io_ins_2(ces_15_16_io_ins_2),
    .io_ins_3(ces_15_16_io_ins_3),
    .io_outs_0(ces_15_16_io_outs_0),
    .io_outs_1(ces_15_16_io_outs_1),
    .io_outs_2(ces_15_16_io_outs_2),
    .io_outs_3(ces_15_16_io_outs_3)
  );
  Element ces_15_17 ( // @[MockArray.scala 36:52]
    .clock(ces_15_17_clock),
    .io_ins_0(ces_15_17_io_ins_0),
    .io_ins_1(ces_15_17_io_ins_1),
    .io_ins_2(ces_15_17_io_ins_2),
    .io_ins_3(ces_15_17_io_ins_3),
    .io_outs_0(ces_15_17_io_outs_0),
    .io_outs_1(ces_15_17_io_outs_1),
    .io_outs_2(ces_15_17_io_outs_2),
    .io_outs_3(ces_15_17_io_outs_3)
  );
  Element ces_15_18 ( // @[MockArray.scala 36:52]
    .clock(ces_15_18_clock),
    .io_ins_0(ces_15_18_io_ins_0),
    .io_ins_1(ces_15_18_io_ins_1),
    .io_ins_2(ces_15_18_io_ins_2),
    .io_ins_3(ces_15_18_io_ins_3),
    .io_outs_0(ces_15_18_io_outs_0),
    .io_outs_1(ces_15_18_io_outs_1),
    .io_outs_2(ces_15_18_io_outs_2),
    .io_outs_3(ces_15_18_io_outs_3)
  );
  Element ces_15_19 ( // @[MockArray.scala 36:52]
    .clock(ces_15_19_clock),
    .io_ins_0(ces_15_19_io_ins_0),
    .io_ins_1(ces_15_19_io_ins_1),
    .io_ins_2(ces_15_19_io_ins_2),
    .io_ins_3(ces_15_19_io_ins_3),
    .io_outs_0(ces_15_19_io_outs_0),
    .io_outs_1(ces_15_19_io_outs_1),
    .io_outs_2(ces_15_19_io_outs_2),
    .io_outs_3(ces_15_19_io_outs_3)
  );
  Element ces_15_20 ( // @[MockArray.scala 36:52]
    .clock(ces_15_20_clock),
    .io_ins_0(ces_15_20_io_ins_0),
    .io_ins_1(ces_15_20_io_ins_1),
    .io_ins_2(ces_15_20_io_ins_2),
    .io_ins_3(ces_15_20_io_ins_3),
    .io_outs_0(ces_15_20_io_outs_0),
    .io_outs_1(ces_15_20_io_outs_1),
    .io_outs_2(ces_15_20_io_outs_2),
    .io_outs_3(ces_15_20_io_outs_3)
  );
  Element ces_15_21 ( // @[MockArray.scala 36:52]
    .clock(ces_15_21_clock),
    .io_ins_0(ces_15_21_io_ins_0),
    .io_ins_1(ces_15_21_io_ins_1),
    .io_ins_2(ces_15_21_io_ins_2),
    .io_ins_3(ces_15_21_io_ins_3),
    .io_outs_0(ces_15_21_io_outs_0),
    .io_outs_1(ces_15_21_io_outs_1),
    .io_outs_2(ces_15_21_io_outs_2),
    .io_outs_3(ces_15_21_io_outs_3)
  );
  Element ces_15_22 ( // @[MockArray.scala 36:52]
    .clock(ces_15_22_clock),
    .io_ins_0(ces_15_22_io_ins_0),
    .io_ins_1(ces_15_22_io_ins_1),
    .io_ins_2(ces_15_22_io_ins_2),
    .io_ins_3(ces_15_22_io_ins_3),
    .io_outs_0(ces_15_22_io_outs_0),
    .io_outs_1(ces_15_22_io_outs_1),
    .io_outs_2(ces_15_22_io_outs_2),
    .io_outs_3(ces_15_22_io_outs_3)
  );
  Element ces_15_23 ( // @[MockArray.scala 36:52]
    .clock(ces_15_23_clock),
    .io_ins_0(ces_15_23_io_ins_0),
    .io_ins_1(ces_15_23_io_ins_1),
    .io_ins_2(ces_15_23_io_ins_2),
    .io_ins_3(ces_15_23_io_ins_3),
    .io_outs_0(ces_15_23_io_outs_0),
    .io_outs_1(ces_15_23_io_outs_1),
    .io_outs_2(ces_15_23_io_outs_2),
    .io_outs_3(ces_15_23_io_outs_3)
  );
  Element ces_15_24 ( // @[MockArray.scala 36:52]
    .clock(ces_15_24_clock),
    .io_ins_0(ces_15_24_io_ins_0),
    .io_ins_1(ces_15_24_io_ins_1),
    .io_ins_2(ces_15_24_io_ins_2),
    .io_ins_3(ces_15_24_io_ins_3),
    .io_outs_0(ces_15_24_io_outs_0),
    .io_outs_1(ces_15_24_io_outs_1),
    .io_outs_2(ces_15_24_io_outs_2),
    .io_outs_3(ces_15_24_io_outs_3)
  );
  Element ces_15_25 ( // @[MockArray.scala 36:52]
    .clock(ces_15_25_clock),
    .io_ins_0(ces_15_25_io_ins_0),
    .io_ins_1(ces_15_25_io_ins_1),
    .io_ins_2(ces_15_25_io_ins_2),
    .io_ins_3(ces_15_25_io_ins_3),
    .io_outs_0(ces_15_25_io_outs_0),
    .io_outs_1(ces_15_25_io_outs_1),
    .io_outs_2(ces_15_25_io_outs_2),
    .io_outs_3(ces_15_25_io_outs_3)
  );
  Element ces_15_26 ( // @[MockArray.scala 36:52]
    .clock(ces_15_26_clock),
    .io_ins_0(ces_15_26_io_ins_0),
    .io_ins_1(ces_15_26_io_ins_1),
    .io_ins_2(ces_15_26_io_ins_2),
    .io_ins_3(ces_15_26_io_ins_3),
    .io_outs_0(ces_15_26_io_outs_0),
    .io_outs_1(ces_15_26_io_outs_1),
    .io_outs_2(ces_15_26_io_outs_2),
    .io_outs_3(ces_15_26_io_outs_3)
  );
  Element ces_15_27 ( // @[MockArray.scala 36:52]
    .clock(ces_15_27_clock),
    .io_ins_0(ces_15_27_io_ins_0),
    .io_ins_1(ces_15_27_io_ins_1),
    .io_ins_2(ces_15_27_io_ins_2),
    .io_ins_3(ces_15_27_io_ins_3),
    .io_outs_0(ces_15_27_io_outs_0),
    .io_outs_1(ces_15_27_io_outs_1),
    .io_outs_2(ces_15_27_io_outs_2),
    .io_outs_3(ces_15_27_io_outs_3)
  );
  Element ces_15_28 ( // @[MockArray.scala 36:52]
    .clock(ces_15_28_clock),
    .io_ins_0(ces_15_28_io_ins_0),
    .io_ins_1(ces_15_28_io_ins_1),
    .io_ins_2(ces_15_28_io_ins_2),
    .io_ins_3(ces_15_28_io_ins_3),
    .io_outs_0(ces_15_28_io_outs_0),
    .io_outs_1(ces_15_28_io_outs_1),
    .io_outs_2(ces_15_28_io_outs_2),
    .io_outs_3(ces_15_28_io_outs_3)
  );
  Element ces_15_29 ( // @[MockArray.scala 36:52]
    .clock(ces_15_29_clock),
    .io_ins_0(ces_15_29_io_ins_0),
    .io_ins_1(ces_15_29_io_ins_1),
    .io_ins_2(ces_15_29_io_ins_2),
    .io_ins_3(ces_15_29_io_ins_3),
    .io_outs_0(ces_15_29_io_outs_0),
    .io_outs_1(ces_15_29_io_outs_1),
    .io_outs_2(ces_15_29_io_outs_2),
    .io_outs_3(ces_15_29_io_outs_3)
  );
  Element ces_15_30 ( // @[MockArray.scala 36:52]
    .clock(ces_15_30_clock),
    .io_ins_0(ces_15_30_io_ins_0),
    .io_ins_1(ces_15_30_io_ins_1),
    .io_ins_2(ces_15_30_io_ins_2),
    .io_ins_3(ces_15_30_io_ins_3),
    .io_outs_0(ces_15_30_io_outs_0),
    .io_outs_1(ces_15_30_io_outs_1),
    .io_outs_2(ces_15_30_io_outs_2),
    .io_outs_3(ces_15_30_io_outs_3)
  );
  Element ces_15_31 ( // @[MockArray.scala 36:52]
    .clock(ces_15_31_clock),
    .io_ins_0(ces_15_31_io_ins_0),
    .io_ins_1(ces_15_31_io_ins_1),
    .io_ins_2(ces_15_31_io_ins_2),
    .io_ins_3(ces_15_31_io_ins_3),
    .io_outs_0(ces_15_31_io_outs_0),
    .io_outs_1(ces_15_31_io_outs_1),
    .io_outs_2(ces_15_31_io_outs_2),
    .io_outs_3(ces_15_31_io_outs_3)
  );
  Element ces_16_0 ( // @[MockArray.scala 36:52]
    .clock(ces_16_0_clock),
    .io_ins_0(ces_16_0_io_ins_0),
    .io_ins_1(ces_16_0_io_ins_1),
    .io_ins_2(ces_16_0_io_ins_2),
    .io_ins_3(ces_16_0_io_ins_3),
    .io_outs_0(ces_16_0_io_outs_0),
    .io_outs_1(ces_16_0_io_outs_1),
    .io_outs_2(ces_16_0_io_outs_2),
    .io_outs_3(ces_16_0_io_outs_3)
  );
  Element ces_16_1 ( // @[MockArray.scala 36:52]
    .clock(ces_16_1_clock),
    .io_ins_0(ces_16_1_io_ins_0),
    .io_ins_1(ces_16_1_io_ins_1),
    .io_ins_2(ces_16_1_io_ins_2),
    .io_ins_3(ces_16_1_io_ins_3),
    .io_outs_0(ces_16_1_io_outs_0),
    .io_outs_1(ces_16_1_io_outs_1),
    .io_outs_2(ces_16_1_io_outs_2),
    .io_outs_3(ces_16_1_io_outs_3)
  );
  Element ces_16_2 ( // @[MockArray.scala 36:52]
    .clock(ces_16_2_clock),
    .io_ins_0(ces_16_2_io_ins_0),
    .io_ins_1(ces_16_2_io_ins_1),
    .io_ins_2(ces_16_2_io_ins_2),
    .io_ins_3(ces_16_2_io_ins_3),
    .io_outs_0(ces_16_2_io_outs_0),
    .io_outs_1(ces_16_2_io_outs_1),
    .io_outs_2(ces_16_2_io_outs_2),
    .io_outs_3(ces_16_2_io_outs_3)
  );
  Element ces_16_3 ( // @[MockArray.scala 36:52]
    .clock(ces_16_3_clock),
    .io_ins_0(ces_16_3_io_ins_0),
    .io_ins_1(ces_16_3_io_ins_1),
    .io_ins_2(ces_16_3_io_ins_2),
    .io_ins_3(ces_16_3_io_ins_3),
    .io_outs_0(ces_16_3_io_outs_0),
    .io_outs_1(ces_16_3_io_outs_1),
    .io_outs_2(ces_16_3_io_outs_2),
    .io_outs_3(ces_16_3_io_outs_3)
  );
  Element ces_16_4 ( // @[MockArray.scala 36:52]
    .clock(ces_16_4_clock),
    .io_ins_0(ces_16_4_io_ins_0),
    .io_ins_1(ces_16_4_io_ins_1),
    .io_ins_2(ces_16_4_io_ins_2),
    .io_ins_3(ces_16_4_io_ins_3),
    .io_outs_0(ces_16_4_io_outs_0),
    .io_outs_1(ces_16_4_io_outs_1),
    .io_outs_2(ces_16_4_io_outs_2),
    .io_outs_3(ces_16_4_io_outs_3)
  );
  Element ces_16_5 ( // @[MockArray.scala 36:52]
    .clock(ces_16_5_clock),
    .io_ins_0(ces_16_5_io_ins_0),
    .io_ins_1(ces_16_5_io_ins_1),
    .io_ins_2(ces_16_5_io_ins_2),
    .io_ins_3(ces_16_5_io_ins_3),
    .io_outs_0(ces_16_5_io_outs_0),
    .io_outs_1(ces_16_5_io_outs_1),
    .io_outs_2(ces_16_5_io_outs_2),
    .io_outs_3(ces_16_5_io_outs_3)
  );
  Element ces_16_6 ( // @[MockArray.scala 36:52]
    .clock(ces_16_6_clock),
    .io_ins_0(ces_16_6_io_ins_0),
    .io_ins_1(ces_16_6_io_ins_1),
    .io_ins_2(ces_16_6_io_ins_2),
    .io_ins_3(ces_16_6_io_ins_3),
    .io_outs_0(ces_16_6_io_outs_0),
    .io_outs_1(ces_16_6_io_outs_1),
    .io_outs_2(ces_16_6_io_outs_2),
    .io_outs_3(ces_16_6_io_outs_3)
  );
  Element ces_16_7 ( // @[MockArray.scala 36:52]
    .clock(ces_16_7_clock),
    .io_ins_0(ces_16_7_io_ins_0),
    .io_ins_1(ces_16_7_io_ins_1),
    .io_ins_2(ces_16_7_io_ins_2),
    .io_ins_3(ces_16_7_io_ins_3),
    .io_outs_0(ces_16_7_io_outs_0),
    .io_outs_1(ces_16_7_io_outs_1),
    .io_outs_2(ces_16_7_io_outs_2),
    .io_outs_3(ces_16_7_io_outs_3)
  );
  Element ces_16_8 ( // @[MockArray.scala 36:52]
    .clock(ces_16_8_clock),
    .io_ins_0(ces_16_8_io_ins_0),
    .io_ins_1(ces_16_8_io_ins_1),
    .io_ins_2(ces_16_8_io_ins_2),
    .io_ins_3(ces_16_8_io_ins_3),
    .io_outs_0(ces_16_8_io_outs_0),
    .io_outs_1(ces_16_8_io_outs_1),
    .io_outs_2(ces_16_8_io_outs_2),
    .io_outs_3(ces_16_8_io_outs_3)
  );
  Element ces_16_9 ( // @[MockArray.scala 36:52]
    .clock(ces_16_9_clock),
    .io_ins_0(ces_16_9_io_ins_0),
    .io_ins_1(ces_16_9_io_ins_1),
    .io_ins_2(ces_16_9_io_ins_2),
    .io_ins_3(ces_16_9_io_ins_3),
    .io_outs_0(ces_16_9_io_outs_0),
    .io_outs_1(ces_16_9_io_outs_1),
    .io_outs_2(ces_16_9_io_outs_2),
    .io_outs_3(ces_16_9_io_outs_3)
  );
  Element ces_16_10 ( // @[MockArray.scala 36:52]
    .clock(ces_16_10_clock),
    .io_ins_0(ces_16_10_io_ins_0),
    .io_ins_1(ces_16_10_io_ins_1),
    .io_ins_2(ces_16_10_io_ins_2),
    .io_ins_3(ces_16_10_io_ins_3),
    .io_outs_0(ces_16_10_io_outs_0),
    .io_outs_1(ces_16_10_io_outs_1),
    .io_outs_2(ces_16_10_io_outs_2),
    .io_outs_3(ces_16_10_io_outs_3)
  );
  Element ces_16_11 ( // @[MockArray.scala 36:52]
    .clock(ces_16_11_clock),
    .io_ins_0(ces_16_11_io_ins_0),
    .io_ins_1(ces_16_11_io_ins_1),
    .io_ins_2(ces_16_11_io_ins_2),
    .io_ins_3(ces_16_11_io_ins_3),
    .io_outs_0(ces_16_11_io_outs_0),
    .io_outs_1(ces_16_11_io_outs_1),
    .io_outs_2(ces_16_11_io_outs_2),
    .io_outs_3(ces_16_11_io_outs_3)
  );
  Element ces_16_12 ( // @[MockArray.scala 36:52]
    .clock(ces_16_12_clock),
    .io_ins_0(ces_16_12_io_ins_0),
    .io_ins_1(ces_16_12_io_ins_1),
    .io_ins_2(ces_16_12_io_ins_2),
    .io_ins_3(ces_16_12_io_ins_3),
    .io_outs_0(ces_16_12_io_outs_0),
    .io_outs_1(ces_16_12_io_outs_1),
    .io_outs_2(ces_16_12_io_outs_2),
    .io_outs_3(ces_16_12_io_outs_3)
  );
  Element ces_16_13 ( // @[MockArray.scala 36:52]
    .clock(ces_16_13_clock),
    .io_ins_0(ces_16_13_io_ins_0),
    .io_ins_1(ces_16_13_io_ins_1),
    .io_ins_2(ces_16_13_io_ins_2),
    .io_ins_3(ces_16_13_io_ins_3),
    .io_outs_0(ces_16_13_io_outs_0),
    .io_outs_1(ces_16_13_io_outs_1),
    .io_outs_2(ces_16_13_io_outs_2),
    .io_outs_3(ces_16_13_io_outs_3)
  );
  Element ces_16_14 ( // @[MockArray.scala 36:52]
    .clock(ces_16_14_clock),
    .io_ins_0(ces_16_14_io_ins_0),
    .io_ins_1(ces_16_14_io_ins_1),
    .io_ins_2(ces_16_14_io_ins_2),
    .io_ins_3(ces_16_14_io_ins_3),
    .io_outs_0(ces_16_14_io_outs_0),
    .io_outs_1(ces_16_14_io_outs_1),
    .io_outs_2(ces_16_14_io_outs_2),
    .io_outs_3(ces_16_14_io_outs_3)
  );
  Element ces_16_15 ( // @[MockArray.scala 36:52]
    .clock(ces_16_15_clock),
    .io_ins_0(ces_16_15_io_ins_0),
    .io_ins_1(ces_16_15_io_ins_1),
    .io_ins_2(ces_16_15_io_ins_2),
    .io_ins_3(ces_16_15_io_ins_3),
    .io_outs_0(ces_16_15_io_outs_0),
    .io_outs_1(ces_16_15_io_outs_1),
    .io_outs_2(ces_16_15_io_outs_2),
    .io_outs_3(ces_16_15_io_outs_3)
  );
  Element ces_16_16 ( // @[MockArray.scala 36:52]
    .clock(ces_16_16_clock),
    .io_ins_0(ces_16_16_io_ins_0),
    .io_ins_1(ces_16_16_io_ins_1),
    .io_ins_2(ces_16_16_io_ins_2),
    .io_ins_3(ces_16_16_io_ins_3),
    .io_outs_0(ces_16_16_io_outs_0),
    .io_outs_1(ces_16_16_io_outs_1),
    .io_outs_2(ces_16_16_io_outs_2),
    .io_outs_3(ces_16_16_io_outs_3)
  );
  Element ces_16_17 ( // @[MockArray.scala 36:52]
    .clock(ces_16_17_clock),
    .io_ins_0(ces_16_17_io_ins_0),
    .io_ins_1(ces_16_17_io_ins_1),
    .io_ins_2(ces_16_17_io_ins_2),
    .io_ins_3(ces_16_17_io_ins_3),
    .io_outs_0(ces_16_17_io_outs_0),
    .io_outs_1(ces_16_17_io_outs_1),
    .io_outs_2(ces_16_17_io_outs_2),
    .io_outs_3(ces_16_17_io_outs_3)
  );
  Element ces_16_18 ( // @[MockArray.scala 36:52]
    .clock(ces_16_18_clock),
    .io_ins_0(ces_16_18_io_ins_0),
    .io_ins_1(ces_16_18_io_ins_1),
    .io_ins_2(ces_16_18_io_ins_2),
    .io_ins_3(ces_16_18_io_ins_3),
    .io_outs_0(ces_16_18_io_outs_0),
    .io_outs_1(ces_16_18_io_outs_1),
    .io_outs_2(ces_16_18_io_outs_2),
    .io_outs_3(ces_16_18_io_outs_3)
  );
  Element ces_16_19 ( // @[MockArray.scala 36:52]
    .clock(ces_16_19_clock),
    .io_ins_0(ces_16_19_io_ins_0),
    .io_ins_1(ces_16_19_io_ins_1),
    .io_ins_2(ces_16_19_io_ins_2),
    .io_ins_3(ces_16_19_io_ins_3),
    .io_outs_0(ces_16_19_io_outs_0),
    .io_outs_1(ces_16_19_io_outs_1),
    .io_outs_2(ces_16_19_io_outs_2),
    .io_outs_3(ces_16_19_io_outs_3)
  );
  Element ces_16_20 ( // @[MockArray.scala 36:52]
    .clock(ces_16_20_clock),
    .io_ins_0(ces_16_20_io_ins_0),
    .io_ins_1(ces_16_20_io_ins_1),
    .io_ins_2(ces_16_20_io_ins_2),
    .io_ins_3(ces_16_20_io_ins_3),
    .io_outs_0(ces_16_20_io_outs_0),
    .io_outs_1(ces_16_20_io_outs_1),
    .io_outs_2(ces_16_20_io_outs_2),
    .io_outs_3(ces_16_20_io_outs_3)
  );
  Element ces_16_21 ( // @[MockArray.scala 36:52]
    .clock(ces_16_21_clock),
    .io_ins_0(ces_16_21_io_ins_0),
    .io_ins_1(ces_16_21_io_ins_1),
    .io_ins_2(ces_16_21_io_ins_2),
    .io_ins_3(ces_16_21_io_ins_3),
    .io_outs_0(ces_16_21_io_outs_0),
    .io_outs_1(ces_16_21_io_outs_1),
    .io_outs_2(ces_16_21_io_outs_2),
    .io_outs_3(ces_16_21_io_outs_3)
  );
  Element ces_16_22 ( // @[MockArray.scala 36:52]
    .clock(ces_16_22_clock),
    .io_ins_0(ces_16_22_io_ins_0),
    .io_ins_1(ces_16_22_io_ins_1),
    .io_ins_2(ces_16_22_io_ins_2),
    .io_ins_3(ces_16_22_io_ins_3),
    .io_outs_0(ces_16_22_io_outs_0),
    .io_outs_1(ces_16_22_io_outs_1),
    .io_outs_2(ces_16_22_io_outs_2),
    .io_outs_3(ces_16_22_io_outs_3)
  );
  Element ces_16_23 ( // @[MockArray.scala 36:52]
    .clock(ces_16_23_clock),
    .io_ins_0(ces_16_23_io_ins_0),
    .io_ins_1(ces_16_23_io_ins_1),
    .io_ins_2(ces_16_23_io_ins_2),
    .io_ins_3(ces_16_23_io_ins_3),
    .io_outs_0(ces_16_23_io_outs_0),
    .io_outs_1(ces_16_23_io_outs_1),
    .io_outs_2(ces_16_23_io_outs_2),
    .io_outs_3(ces_16_23_io_outs_3)
  );
  Element ces_16_24 ( // @[MockArray.scala 36:52]
    .clock(ces_16_24_clock),
    .io_ins_0(ces_16_24_io_ins_0),
    .io_ins_1(ces_16_24_io_ins_1),
    .io_ins_2(ces_16_24_io_ins_2),
    .io_ins_3(ces_16_24_io_ins_3),
    .io_outs_0(ces_16_24_io_outs_0),
    .io_outs_1(ces_16_24_io_outs_1),
    .io_outs_2(ces_16_24_io_outs_2),
    .io_outs_3(ces_16_24_io_outs_3)
  );
  Element ces_16_25 ( // @[MockArray.scala 36:52]
    .clock(ces_16_25_clock),
    .io_ins_0(ces_16_25_io_ins_0),
    .io_ins_1(ces_16_25_io_ins_1),
    .io_ins_2(ces_16_25_io_ins_2),
    .io_ins_3(ces_16_25_io_ins_3),
    .io_outs_0(ces_16_25_io_outs_0),
    .io_outs_1(ces_16_25_io_outs_1),
    .io_outs_2(ces_16_25_io_outs_2),
    .io_outs_3(ces_16_25_io_outs_3)
  );
  Element ces_16_26 ( // @[MockArray.scala 36:52]
    .clock(ces_16_26_clock),
    .io_ins_0(ces_16_26_io_ins_0),
    .io_ins_1(ces_16_26_io_ins_1),
    .io_ins_2(ces_16_26_io_ins_2),
    .io_ins_3(ces_16_26_io_ins_3),
    .io_outs_0(ces_16_26_io_outs_0),
    .io_outs_1(ces_16_26_io_outs_1),
    .io_outs_2(ces_16_26_io_outs_2),
    .io_outs_3(ces_16_26_io_outs_3)
  );
  Element ces_16_27 ( // @[MockArray.scala 36:52]
    .clock(ces_16_27_clock),
    .io_ins_0(ces_16_27_io_ins_0),
    .io_ins_1(ces_16_27_io_ins_1),
    .io_ins_2(ces_16_27_io_ins_2),
    .io_ins_3(ces_16_27_io_ins_3),
    .io_outs_0(ces_16_27_io_outs_0),
    .io_outs_1(ces_16_27_io_outs_1),
    .io_outs_2(ces_16_27_io_outs_2),
    .io_outs_3(ces_16_27_io_outs_3)
  );
  Element ces_16_28 ( // @[MockArray.scala 36:52]
    .clock(ces_16_28_clock),
    .io_ins_0(ces_16_28_io_ins_0),
    .io_ins_1(ces_16_28_io_ins_1),
    .io_ins_2(ces_16_28_io_ins_2),
    .io_ins_3(ces_16_28_io_ins_3),
    .io_outs_0(ces_16_28_io_outs_0),
    .io_outs_1(ces_16_28_io_outs_1),
    .io_outs_2(ces_16_28_io_outs_2),
    .io_outs_3(ces_16_28_io_outs_3)
  );
  Element ces_16_29 ( // @[MockArray.scala 36:52]
    .clock(ces_16_29_clock),
    .io_ins_0(ces_16_29_io_ins_0),
    .io_ins_1(ces_16_29_io_ins_1),
    .io_ins_2(ces_16_29_io_ins_2),
    .io_ins_3(ces_16_29_io_ins_3),
    .io_outs_0(ces_16_29_io_outs_0),
    .io_outs_1(ces_16_29_io_outs_1),
    .io_outs_2(ces_16_29_io_outs_2),
    .io_outs_3(ces_16_29_io_outs_3)
  );
  Element ces_16_30 ( // @[MockArray.scala 36:52]
    .clock(ces_16_30_clock),
    .io_ins_0(ces_16_30_io_ins_0),
    .io_ins_1(ces_16_30_io_ins_1),
    .io_ins_2(ces_16_30_io_ins_2),
    .io_ins_3(ces_16_30_io_ins_3),
    .io_outs_0(ces_16_30_io_outs_0),
    .io_outs_1(ces_16_30_io_outs_1),
    .io_outs_2(ces_16_30_io_outs_2),
    .io_outs_3(ces_16_30_io_outs_3)
  );
  Element ces_16_31 ( // @[MockArray.scala 36:52]
    .clock(ces_16_31_clock),
    .io_ins_0(ces_16_31_io_ins_0),
    .io_ins_1(ces_16_31_io_ins_1),
    .io_ins_2(ces_16_31_io_ins_2),
    .io_ins_3(ces_16_31_io_ins_3),
    .io_outs_0(ces_16_31_io_outs_0),
    .io_outs_1(ces_16_31_io_outs_1),
    .io_outs_2(ces_16_31_io_outs_2),
    .io_outs_3(ces_16_31_io_outs_3)
  );
  Element ces_17_0 ( // @[MockArray.scala 36:52]
    .clock(ces_17_0_clock),
    .io_ins_0(ces_17_0_io_ins_0),
    .io_ins_1(ces_17_0_io_ins_1),
    .io_ins_2(ces_17_0_io_ins_2),
    .io_ins_3(ces_17_0_io_ins_3),
    .io_outs_0(ces_17_0_io_outs_0),
    .io_outs_1(ces_17_0_io_outs_1),
    .io_outs_2(ces_17_0_io_outs_2),
    .io_outs_3(ces_17_0_io_outs_3)
  );
  Element ces_17_1 ( // @[MockArray.scala 36:52]
    .clock(ces_17_1_clock),
    .io_ins_0(ces_17_1_io_ins_0),
    .io_ins_1(ces_17_1_io_ins_1),
    .io_ins_2(ces_17_1_io_ins_2),
    .io_ins_3(ces_17_1_io_ins_3),
    .io_outs_0(ces_17_1_io_outs_0),
    .io_outs_1(ces_17_1_io_outs_1),
    .io_outs_2(ces_17_1_io_outs_2),
    .io_outs_3(ces_17_1_io_outs_3)
  );
  Element ces_17_2 ( // @[MockArray.scala 36:52]
    .clock(ces_17_2_clock),
    .io_ins_0(ces_17_2_io_ins_0),
    .io_ins_1(ces_17_2_io_ins_1),
    .io_ins_2(ces_17_2_io_ins_2),
    .io_ins_3(ces_17_2_io_ins_3),
    .io_outs_0(ces_17_2_io_outs_0),
    .io_outs_1(ces_17_2_io_outs_1),
    .io_outs_2(ces_17_2_io_outs_2),
    .io_outs_3(ces_17_2_io_outs_3)
  );
  Element ces_17_3 ( // @[MockArray.scala 36:52]
    .clock(ces_17_3_clock),
    .io_ins_0(ces_17_3_io_ins_0),
    .io_ins_1(ces_17_3_io_ins_1),
    .io_ins_2(ces_17_3_io_ins_2),
    .io_ins_3(ces_17_3_io_ins_3),
    .io_outs_0(ces_17_3_io_outs_0),
    .io_outs_1(ces_17_3_io_outs_1),
    .io_outs_2(ces_17_3_io_outs_2),
    .io_outs_3(ces_17_3_io_outs_3)
  );
  Element ces_17_4 ( // @[MockArray.scala 36:52]
    .clock(ces_17_4_clock),
    .io_ins_0(ces_17_4_io_ins_0),
    .io_ins_1(ces_17_4_io_ins_1),
    .io_ins_2(ces_17_4_io_ins_2),
    .io_ins_3(ces_17_4_io_ins_3),
    .io_outs_0(ces_17_4_io_outs_0),
    .io_outs_1(ces_17_4_io_outs_1),
    .io_outs_2(ces_17_4_io_outs_2),
    .io_outs_3(ces_17_4_io_outs_3)
  );
  Element ces_17_5 ( // @[MockArray.scala 36:52]
    .clock(ces_17_5_clock),
    .io_ins_0(ces_17_5_io_ins_0),
    .io_ins_1(ces_17_5_io_ins_1),
    .io_ins_2(ces_17_5_io_ins_2),
    .io_ins_3(ces_17_5_io_ins_3),
    .io_outs_0(ces_17_5_io_outs_0),
    .io_outs_1(ces_17_5_io_outs_1),
    .io_outs_2(ces_17_5_io_outs_2),
    .io_outs_3(ces_17_5_io_outs_3)
  );
  Element ces_17_6 ( // @[MockArray.scala 36:52]
    .clock(ces_17_6_clock),
    .io_ins_0(ces_17_6_io_ins_0),
    .io_ins_1(ces_17_6_io_ins_1),
    .io_ins_2(ces_17_6_io_ins_2),
    .io_ins_3(ces_17_6_io_ins_3),
    .io_outs_0(ces_17_6_io_outs_0),
    .io_outs_1(ces_17_6_io_outs_1),
    .io_outs_2(ces_17_6_io_outs_2),
    .io_outs_3(ces_17_6_io_outs_3)
  );
  Element ces_17_7 ( // @[MockArray.scala 36:52]
    .clock(ces_17_7_clock),
    .io_ins_0(ces_17_7_io_ins_0),
    .io_ins_1(ces_17_7_io_ins_1),
    .io_ins_2(ces_17_7_io_ins_2),
    .io_ins_3(ces_17_7_io_ins_3),
    .io_outs_0(ces_17_7_io_outs_0),
    .io_outs_1(ces_17_7_io_outs_1),
    .io_outs_2(ces_17_7_io_outs_2),
    .io_outs_3(ces_17_7_io_outs_3)
  );
  Element ces_17_8 ( // @[MockArray.scala 36:52]
    .clock(ces_17_8_clock),
    .io_ins_0(ces_17_8_io_ins_0),
    .io_ins_1(ces_17_8_io_ins_1),
    .io_ins_2(ces_17_8_io_ins_2),
    .io_ins_3(ces_17_8_io_ins_3),
    .io_outs_0(ces_17_8_io_outs_0),
    .io_outs_1(ces_17_8_io_outs_1),
    .io_outs_2(ces_17_8_io_outs_2),
    .io_outs_3(ces_17_8_io_outs_3)
  );
  Element ces_17_9 ( // @[MockArray.scala 36:52]
    .clock(ces_17_9_clock),
    .io_ins_0(ces_17_9_io_ins_0),
    .io_ins_1(ces_17_9_io_ins_1),
    .io_ins_2(ces_17_9_io_ins_2),
    .io_ins_3(ces_17_9_io_ins_3),
    .io_outs_0(ces_17_9_io_outs_0),
    .io_outs_1(ces_17_9_io_outs_1),
    .io_outs_2(ces_17_9_io_outs_2),
    .io_outs_3(ces_17_9_io_outs_3)
  );
  Element ces_17_10 ( // @[MockArray.scala 36:52]
    .clock(ces_17_10_clock),
    .io_ins_0(ces_17_10_io_ins_0),
    .io_ins_1(ces_17_10_io_ins_1),
    .io_ins_2(ces_17_10_io_ins_2),
    .io_ins_3(ces_17_10_io_ins_3),
    .io_outs_0(ces_17_10_io_outs_0),
    .io_outs_1(ces_17_10_io_outs_1),
    .io_outs_2(ces_17_10_io_outs_2),
    .io_outs_3(ces_17_10_io_outs_3)
  );
  Element ces_17_11 ( // @[MockArray.scala 36:52]
    .clock(ces_17_11_clock),
    .io_ins_0(ces_17_11_io_ins_0),
    .io_ins_1(ces_17_11_io_ins_1),
    .io_ins_2(ces_17_11_io_ins_2),
    .io_ins_3(ces_17_11_io_ins_3),
    .io_outs_0(ces_17_11_io_outs_0),
    .io_outs_1(ces_17_11_io_outs_1),
    .io_outs_2(ces_17_11_io_outs_2),
    .io_outs_3(ces_17_11_io_outs_3)
  );
  Element ces_17_12 ( // @[MockArray.scala 36:52]
    .clock(ces_17_12_clock),
    .io_ins_0(ces_17_12_io_ins_0),
    .io_ins_1(ces_17_12_io_ins_1),
    .io_ins_2(ces_17_12_io_ins_2),
    .io_ins_3(ces_17_12_io_ins_3),
    .io_outs_0(ces_17_12_io_outs_0),
    .io_outs_1(ces_17_12_io_outs_1),
    .io_outs_2(ces_17_12_io_outs_2),
    .io_outs_3(ces_17_12_io_outs_3)
  );
  Element ces_17_13 ( // @[MockArray.scala 36:52]
    .clock(ces_17_13_clock),
    .io_ins_0(ces_17_13_io_ins_0),
    .io_ins_1(ces_17_13_io_ins_1),
    .io_ins_2(ces_17_13_io_ins_2),
    .io_ins_3(ces_17_13_io_ins_3),
    .io_outs_0(ces_17_13_io_outs_0),
    .io_outs_1(ces_17_13_io_outs_1),
    .io_outs_2(ces_17_13_io_outs_2),
    .io_outs_3(ces_17_13_io_outs_3)
  );
  Element ces_17_14 ( // @[MockArray.scala 36:52]
    .clock(ces_17_14_clock),
    .io_ins_0(ces_17_14_io_ins_0),
    .io_ins_1(ces_17_14_io_ins_1),
    .io_ins_2(ces_17_14_io_ins_2),
    .io_ins_3(ces_17_14_io_ins_3),
    .io_outs_0(ces_17_14_io_outs_0),
    .io_outs_1(ces_17_14_io_outs_1),
    .io_outs_2(ces_17_14_io_outs_2),
    .io_outs_3(ces_17_14_io_outs_3)
  );
  Element ces_17_15 ( // @[MockArray.scala 36:52]
    .clock(ces_17_15_clock),
    .io_ins_0(ces_17_15_io_ins_0),
    .io_ins_1(ces_17_15_io_ins_1),
    .io_ins_2(ces_17_15_io_ins_2),
    .io_ins_3(ces_17_15_io_ins_3),
    .io_outs_0(ces_17_15_io_outs_0),
    .io_outs_1(ces_17_15_io_outs_1),
    .io_outs_2(ces_17_15_io_outs_2),
    .io_outs_3(ces_17_15_io_outs_3)
  );
  Element ces_17_16 ( // @[MockArray.scala 36:52]
    .clock(ces_17_16_clock),
    .io_ins_0(ces_17_16_io_ins_0),
    .io_ins_1(ces_17_16_io_ins_1),
    .io_ins_2(ces_17_16_io_ins_2),
    .io_ins_3(ces_17_16_io_ins_3),
    .io_outs_0(ces_17_16_io_outs_0),
    .io_outs_1(ces_17_16_io_outs_1),
    .io_outs_2(ces_17_16_io_outs_2),
    .io_outs_3(ces_17_16_io_outs_3)
  );
  Element ces_17_17 ( // @[MockArray.scala 36:52]
    .clock(ces_17_17_clock),
    .io_ins_0(ces_17_17_io_ins_0),
    .io_ins_1(ces_17_17_io_ins_1),
    .io_ins_2(ces_17_17_io_ins_2),
    .io_ins_3(ces_17_17_io_ins_3),
    .io_outs_0(ces_17_17_io_outs_0),
    .io_outs_1(ces_17_17_io_outs_1),
    .io_outs_2(ces_17_17_io_outs_2),
    .io_outs_3(ces_17_17_io_outs_3)
  );
  Element ces_17_18 ( // @[MockArray.scala 36:52]
    .clock(ces_17_18_clock),
    .io_ins_0(ces_17_18_io_ins_0),
    .io_ins_1(ces_17_18_io_ins_1),
    .io_ins_2(ces_17_18_io_ins_2),
    .io_ins_3(ces_17_18_io_ins_3),
    .io_outs_0(ces_17_18_io_outs_0),
    .io_outs_1(ces_17_18_io_outs_1),
    .io_outs_2(ces_17_18_io_outs_2),
    .io_outs_3(ces_17_18_io_outs_3)
  );
  Element ces_17_19 ( // @[MockArray.scala 36:52]
    .clock(ces_17_19_clock),
    .io_ins_0(ces_17_19_io_ins_0),
    .io_ins_1(ces_17_19_io_ins_1),
    .io_ins_2(ces_17_19_io_ins_2),
    .io_ins_3(ces_17_19_io_ins_3),
    .io_outs_0(ces_17_19_io_outs_0),
    .io_outs_1(ces_17_19_io_outs_1),
    .io_outs_2(ces_17_19_io_outs_2),
    .io_outs_3(ces_17_19_io_outs_3)
  );
  Element ces_17_20 ( // @[MockArray.scala 36:52]
    .clock(ces_17_20_clock),
    .io_ins_0(ces_17_20_io_ins_0),
    .io_ins_1(ces_17_20_io_ins_1),
    .io_ins_2(ces_17_20_io_ins_2),
    .io_ins_3(ces_17_20_io_ins_3),
    .io_outs_0(ces_17_20_io_outs_0),
    .io_outs_1(ces_17_20_io_outs_1),
    .io_outs_2(ces_17_20_io_outs_2),
    .io_outs_3(ces_17_20_io_outs_3)
  );
  Element ces_17_21 ( // @[MockArray.scala 36:52]
    .clock(ces_17_21_clock),
    .io_ins_0(ces_17_21_io_ins_0),
    .io_ins_1(ces_17_21_io_ins_1),
    .io_ins_2(ces_17_21_io_ins_2),
    .io_ins_3(ces_17_21_io_ins_3),
    .io_outs_0(ces_17_21_io_outs_0),
    .io_outs_1(ces_17_21_io_outs_1),
    .io_outs_2(ces_17_21_io_outs_2),
    .io_outs_3(ces_17_21_io_outs_3)
  );
  Element ces_17_22 ( // @[MockArray.scala 36:52]
    .clock(ces_17_22_clock),
    .io_ins_0(ces_17_22_io_ins_0),
    .io_ins_1(ces_17_22_io_ins_1),
    .io_ins_2(ces_17_22_io_ins_2),
    .io_ins_3(ces_17_22_io_ins_3),
    .io_outs_0(ces_17_22_io_outs_0),
    .io_outs_1(ces_17_22_io_outs_1),
    .io_outs_2(ces_17_22_io_outs_2),
    .io_outs_3(ces_17_22_io_outs_3)
  );
  Element ces_17_23 ( // @[MockArray.scala 36:52]
    .clock(ces_17_23_clock),
    .io_ins_0(ces_17_23_io_ins_0),
    .io_ins_1(ces_17_23_io_ins_1),
    .io_ins_2(ces_17_23_io_ins_2),
    .io_ins_3(ces_17_23_io_ins_3),
    .io_outs_0(ces_17_23_io_outs_0),
    .io_outs_1(ces_17_23_io_outs_1),
    .io_outs_2(ces_17_23_io_outs_2),
    .io_outs_3(ces_17_23_io_outs_3)
  );
  Element ces_17_24 ( // @[MockArray.scala 36:52]
    .clock(ces_17_24_clock),
    .io_ins_0(ces_17_24_io_ins_0),
    .io_ins_1(ces_17_24_io_ins_1),
    .io_ins_2(ces_17_24_io_ins_2),
    .io_ins_3(ces_17_24_io_ins_3),
    .io_outs_0(ces_17_24_io_outs_0),
    .io_outs_1(ces_17_24_io_outs_1),
    .io_outs_2(ces_17_24_io_outs_2),
    .io_outs_3(ces_17_24_io_outs_3)
  );
  Element ces_17_25 ( // @[MockArray.scala 36:52]
    .clock(ces_17_25_clock),
    .io_ins_0(ces_17_25_io_ins_0),
    .io_ins_1(ces_17_25_io_ins_1),
    .io_ins_2(ces_17_25_io_ins_2),
    .io_ins_3(ces_17_25_io_ins_3),
    .io_outs_0(ces_17_25_io_outs_0),
    .io_outs_1(ces_17_25_io_outs_1),
    .io_outs_2(ces_17_25_io_outs_2),
    .io_outs_3(ces_17_25_io_outs_3)
  );
  Element ces_17_26 ( // @[MockArray.scala 36:52]
    .clock(ces_17_26_clock),
    .io_ins_0(ces_17_26_io_ins_0),
    .io_ins_1(ces_17_26_io_ins_1),
    .io_ins_2(ces_17_26_io_ins_2),
    .io_ins_3(ces_17_26_io_ins_3),
    .io_outs_0(ces_17_26_io_outs_0),
    .io_outs_1(ces_17_26_io_outs_1),
    .io_outs_2(ces_17_26_io_outs_2),
    .io_outs_3(ces_17_26_io_outs_3)
  );
  Element ces_17_27 ( // @[MockArray.scala 36:52]
    .clock(ces_17_27_clock),
    .io_ins_0(ces_17_27_io_ins_0),
    .io_ins_1(ces_17_27_io_ins_1),
    .io_ins_2(ces_17_27_io_ins_2),
    .io_ins_3(ces_17_27_io_ins_3),
    .io_outs_0(ces_17_27_io_outs_0),
    .io_outs_1(ces_17_27_io_outs_1),
    .io_outs_2(ces_17_27_io_outs_2),
    .io_outs_3(ces_17_27_io_outs_3)
  );
  Element ces_17_28 ( // @[MockArray.scala 36:52]
    .clock(ces_17_28_clock),
    .io_ins_0(ces_17_28_io_ins_0),
    .io_ins_1(ces_17_28_io_ins_1),
    .io_ins_2(ces_17_28_io_ins_2),
    .io_ins_3(ces_17_28_io_ins_3),
    .io_outs_0(ces_17_28_io_outs_0),
    .io_outs_1(ces_17_28_io_outs_1),
    .io_outs_2(ces_17_28_io_outs_2),
    .io_outs_3(ces_17_28_io_outs_3)
  );
  Element ces_17_29 ( // @[MockArray.scala 36:52]
    .clock(ces_17_29_clock),
    .io_ins_0(ces_17_29_io_ins_0),
    .io_ins_1(ces_17_29_io_ins_1),
    .io_ins_2(ces_17_29_io_ins_2),
    .io_ins_3(ces_17_29_io_ins_3),
    .io_outs_0(ces_17_29_io_outs_0),
    .io_outs_1(ces_17_29_io_outs_1),
    .io_outs_2(ces_17_29_io_outs_2),
    .io_outs_3(ces_17_29_io_outs_3)
  );
  Element ces_17_30 ( // @[MockArray.scala 36:52]
    .clock(ces_17_30_clock),
    .io_ins_0(ces_17_30_io_ins_0),
    .io_ins_1(ces_17_30_io_ins_1),
    .io_ins_2(ces_17_30_io_ins_2),
    .io_ins_3(ces_17_30_io_ins_3),
    .io_outs_0(ces_17_30_io_outs_0),
    .io_outs_1(ces_17_30_io_outs_1),
    .io_outs_2(ces_17_30_io_outs_2),
    .io_outs_3(ces_17_30_io_outs_3)
  );
  Element ces_17_31 ( // @[MockArray.scala 36:52]
    .clock(ces_17_31_clock),
    .io_ins_0(ces_17_31_io_ins_0),
    .io_ins_1(ces_17_31_io_ins_1),
    .io_ins_2(ces_17_31_io_ins_2),
    .io_ins_3(ces_17_31_io_ins_3),
    .io_outs_0(ces_17_31_io_outs_0),
    .io_outs_1(ces_17_31_io_outs_1),
    .io_outs_2(ces_17_31_io_outs_2),
    .io_outs_3(ces_17_31_io_outs_3)
  );
  Element ces_18_0 ( // @[MockArray.scala 36:52]
    .clock(ces_18_0_clock),
    .io_ins_0(ces_18_0_io_ins_0),
    .io_ins_1(ces_18_0_io_ins_1),
    .io_ins_2(ces_18_0_io_ins_2),
    .io_ins_3(ces_18_0_io_ins_3),
    .io_outs_0(ces_18_0_io_outs_0),
    .io_outs_1(ces_18_0_io_outs_1),
    .io_outs_2(ces_18_0_io_outs_2),
    .io_outs_3(ces_18_0_io_outs_3)
  );
  Element ces_18_1 ( // @[MockArray.scala 36:52]
    .clock(ces_18_1_clock),
    .io_ins_0(ces_18_1_io_ins_0),
    .io_ins_1(ces_18_1_io_ins_1),
    .io_ins_2(ces_18_1_io_ins_2),
    .io_ins_3(ces_18_1_io_ins_3),
    .io_outs_0(ces_18_1_io_outs_0),
    .io_outs_1(ces_18_1_io_outs_1),
    .io_outs_2(ces_18_1_io_outs_2),
    .io_outs_3(ces_18_1_io_outs_3)
  );
  Element ces_18_2 ( // @[MockArray.scala 36:52]
    .clock(ces_18_2_clock),
    .io_ins_0(ces_18_2_io_ins_0),
    .io_ins_1(ces_18_2_io_ins_1),
    .io_ins_2(ces_18_2_io_ins_2),
    .io_ins_3(ces_18_2_io_ins_3),
    .io_outs_0(ces_18_2_io_outs_0),
    .io_outs_1(ces_18_2_io_outs_1),
    .io_outs_2(ces_18_2_io_outs_2),
    .io_outs_3(ces_18_2_io_outs_3)
  );
  Element ces_18_3 ( // @[MockArray.scala 36:52]
    .clock(ces_18_3_clock),
    .io_ins_0(ces_18_3_io_ins_0),
    .io_ins_1(ces_18_3_io_ins_1),
    .io_ins_2(ces_18_3_io_ins_2),
    .io_ins_3(ces_18_3_io_ins_3),
    .io_outs_0(ces_18_3_io_outs_0),
    .io_outs_1(ces_18_3_io_outs_1),
    .io_outs_2(ces_18_3_io_outs_2),
    .io_outs_3(ces_18_3_io_outs_3)
  );
  Element ces_18_4 ( // @[MockArray.scala 36:52]
    .clock(ces_18_4_clock),
    .io_ins_0(ces_18_4_io_ins_0),
    .io_ins_1(ces_18_4_io_ins_1),
    .io_ins_2(ces_18_4_io_ins_2),
    .io_ins_3(ces_18_4_io_ins_3),
    .io_outs_0(ces_18_4_io_outs_0),
    .io_outs_1(ces_18_4_io_outs_1),
    .io_outs_2(ces_18_4_io_outs_2),
    .io_outs_3(ces_18_4_io_outs_3)
  );
  Element ces_18_5 ( // @[MockArray.scala 36:52]
    .clock(ces_18_5_clock),
    .io_ins_0(ces_18_5_io_ins_0),
    .io_ins_1(ces_18_5_io_ins_1),
    .io_ins_2(ces_18_5_io_ins_2),
    .io_ins_3(ces_18_5_io_ins_3),
    .io_outs_0(ces_18_5_io_outs_0),
    .io_outs_1(ces_18_5_io_outs_1),
    .io_outs_2(ces_18_5_io_outs_2),
    .io_outs_3(ces_18_5_io_outs_3)
  );
  Element ces_18_6 ( // @[MockArray.scala 36:52]
    .clock(ces_18_6_clock),
    .io_ins_0(ces_18_6_io_ins_0),
    .io_ins_1(ces_18_6_io_ins_1),
    .io_ins_2(ces_18_6_io_ins_2),
    .io_ins_3(ces_18_6_io_ins_3),
    .io_outs_0(ces_18_6_io_outs_0),
    .io_outs_1(ces_18_6_io_outs_1),
    .io_outs_2(ces_18_6_io_outs_2),
    .io_outs_3(ces_18_6_io_outs_3)
  );
  Element ces_18_7 ( // @[MockArray.scala 36:52]
    .clock(ces_18_7_clock),
    .io_ins_0(ces_18_7_io_ins_0),
    .io_ins_1(ces_18_7_io_ins_1),
    .io_ins_2(ces_18_7_io_ins_2),
    .io_ins_3(ces_18_7_io_ins_3),
    .io_outs_0(ces_18_7_io_outs_0),
    .io_outs_1(ces_18_7_io_outs_1),
    .io_outs_2(ces_18_7_io_outs_2),
    .io_outs_3(ces_18_7_io_outs_3)
  );
  Element ces_18_8 ( // @[MockArray.scala 36:52]
    .clock(ces_18_8_clock),
    .io_ins_0(ces_18_8_io_ins_0),
    .io_ins_1(ces_18_8_io_ins_1),
    .io_ins_2(ces_18_8_io_ins_2),
    .io_ins_3(ces_18_8_io_ins_3),
    .io_outs_0(ces_18_8_io_outs_0),
    .io_outs_1(ces_18_8_io_outs_1),
    .io_outs_2(ces_18_8_io_outs_2),
    .io_outs_3(ces_18_8_io_outs_3)
  );
  Element ces_18_9 ( // @[MockArray.scala 36:52]
    .clock(ces_18_9_clock),
    .io_ins_0(ces_18_9_io_ins_0),
    .io_ins_1(ces_18_9_io_ins_1),
    .io_ins_2(ces_18_9_io_ins_2),
    .io_ins_3(ces_18_9_io_ins_3),
    .io_outs_0(ces_18_9_io_outs_0),
    .io_outs_1(ces_18_9_io_outs_1),
    .io_outs_2(ces_18_9_io_outs_2),
    .io_outs_3(ces_18_9_io_outs_3)
  );
  Element ces_18_10 ( // @[MockArray.scala 36:52]
    .clock(ces_18_10_clock),
    .io_ins_0(ces_18_10_io_ins_0),
    .io_ins_1(ces_18_10_io_ins_1),
    .io_ins_2(ces_18_10_io_ins_2),
    .io_ins_3(ces_18_10_io_ins_3),
    .io_outs_0(ces_18_10_io_outs_0),
    .io_outs_1(ces_18_10_io_outs_1),
    .io_outs_2(ces_18_10_io_outs_2),
    .io_outs_3(ces_18_10_io_outs_3)
  );
  Element ces_18_11 ( // @[MockArray.scala 36:52]
    .clock(ces_18_11_clock),
    .io_ins_0(ces_18_11_io_ins_0),
    .io_ins_1(ces_18_11_io_ins_1),
    .io_ins_2(ces_18_11_io_ins_2),
    .io_ins_3(ces_18_11_io_ins_3),
    .io_outs_0(ces_18_11_io_outs_0),
    .io_outs_1(ces_18_11_io_outs_1),
    .io_outs_2(ces_18_11_io_outs_2),
    .io_outs_3(ces_18_11_io_outs_3)
  );
  Element ces_18_12 ( // @[MockArray.scala 36:52]
    .clock(ces_18_12_clock),
    .io_ins_0(ces_18_12_io_ins_0),
    .io_ins_1(ces_18_12_io_ins_1),
    .io_ins_2(ces_18_12_io_ins_2),
    .io_ins_3(ces_18_12_io_ins_3),
    .io_outs_0(ces_18_12_io_outs_0),
    .io_outs_1(ces_18_12_io_outs_1),
    .io_outs_2(ces_18_12_io_outs_2),
    .io_outs_3(ces_18_12_io_outs_3)
  );
  Element ces_18_13 ( // @[MockArray.scala 36:52]
    .clock(ces_18_13_clock),
    .io_ins_0(ces_18_13_io_ins_0),
    .io_ins_1(ces_18_13_io_ins_1),
    .io_ins_2(ces_18_13_io_ins_2),
    .io_ins_3(ces_18_13_io_ins_3),
    .io_outs_0(ces_18_13_io_outs_0),
    .io_outs_1(ces_18_13_io_outs_1),
    .io_outs_2(ces_18_13_io_outs_2),
    .io_outs_3(ces_18_13_io_outs_3)
  );
  Element ces_18_14 ( // @[MockArray.scala 36:52]
    .clock(ces_18_14_clock),
    .io_ins_0(ces_18_14_io_ins_0),
    .io_ins_1(ces_18_14_io_ins_1),
    .io_ins_2(ces_18_14_io_ins_2),
    .io_ins_3(ces_18_14_io_ins_3),
    .io_outs_0(ces_18_14_io_outs_0),
    .io_outs_1(ces_18_14_io_outs_1),
    .io_outs_2(ces_18_14_io_outs_2),
    .io_outs_3(ces_18_14_io_outs_3)
  );
  Element ces_18_15 ( // @[MockArray.scala 36:52]
    .clock(ces_18_15_clock),
    .io_ins_0(ces_18_15_io_ins_0),
    .io_ins_1(ces_18_15_io_ins_1),
    .io_ins_2(ces_18_15_io_ins_2),
    .io_ins_3(ces_18_15_io_ins_3),
    .io_outs_0(ces_18_15_io_outs_0),
    .io_outs_1(ces_18_15_io_outs_1),
    .io_outs_2(ces_18_15_io_outs_2),
    .io_outs_3(ces_18_15_io_outs_3)
  );
  Element ces_18_16 ( // @[MockArray.scala 36:52]
    .clock(ces_18_16_clock),
    .io_ins_0(ces_18_16_io_ins_0),
    .io_ins_1(ces_18_16_io_ins_1),
    .io_ins_2(ces_18_16_io_ins_2),
    .io_ins_3(ces_18_16_io_ins_3),
    .io_outs_0(ces_18_16_io_outs_0),
    .io_outs_1(ces_18_16_io_outs_1),
    .io_outs_2(ces_18_16_io_outs_2),
    .io_outs_3(ces_18_16_io_outs_3)
  );
  Element ces_18_17 ( // @[MockArray.scala 36:52]
    .clock(ces_18_17_clock),
    .io_ins_0(ces_18_17_io_ins_0),
    .io_ins_1(ces_18_17_io_ins_1),
    .io_ins_2(ces_18_17_io_ins_2),
    .io_ins_3(ces_18_17_io_ins_3),
    .io_outs_0(ces_18_17_io_outs_0),
    .io_outs_1(ces_18_17_io_outs_1),
    .io_outs_2(ces_18_17_io_outs_2),
    .io_outs_3(ces_18_17_io_outs_3)
  );
  Element ces_18_18 ( // @[MockArray.scala 36:52]
    .clock(ces_18_18_clock),
    .io_ins_0(ces_18_18_io_ins_0),
    .io_ins_1(ces_18_18_io_ins_1),
    .io_ins_2(ces_18_18_io_ins_2),
    .io_ins_3(ces_18_18_io_ins_3),
    .io_outs_0(ces_18_18_io_outs_0),
    .io_outs_1(ces_18_18_io_outs_1),
    .io_outs_2(ces_18_18_io_outs_2),
    .io_outs_3(ces_18_18_io_outs_3)
  );
  Element ces_18_19 ( // @[MockArray.scala 36:52]
    .clock(ces_18_19_clock),
    .io_ins_0(ces_18_19_io_ins_0),
    .io_ins_1(ces_18_19_io_ins_1),
    .io_ins_2(ces_18_19_io_ins_2),
    .io_ins_3(ces_18_19_io_ins_3),
    .io_outs_0(ces_18_19_io_outs_0),
    .io_outs_1(ces_18_19_io_outs_1),
    .io_outs_2(ces_18_19_io_outs_2),
    .io_outs_3(ces_18_19_io_outs_3)
  );
  Element ces_18_20 ( // @[MockArray.scala 36:52]
    .clock(ces_18_20_clock),
    .io_ins_0(ces_18_20_io_ins_0),
    .io_ins_1(ces_18_20_io_ins_1),
    .io_ins_2(ces_18_20_io_ins_2),
    .io_ins_3(ces_18_20_io_ins_3),
    .io_outs_0(ces_18_20_io_outs_0),
    .io_outs_1(ces_18_20_io_outs_1),
    .io_outs_2(ces_18_20_io_outs_2),
    .io_outs_3(ces_18_20_io_outs_3)
  );
  Element ces_18_21 ( // @[MockArray.scala 36:52]
    .clock(ces_18_21_clock),
    .io_ins_0(ces_18_21_io_ins_0),
    .io_ins_1(ces_18_21_io_ins_1),
    .io_ins_2(ces_18_21_io_ins_2),
    .io_ins_3(ces_18_21_io_ins_3),
    .io_outs_0(ces_18_21_io_outs_0),
    .io_outs_1(ces_18_21_io_outs_1),
    .io_outs_2(ces_18_21_io_outs_2),
    .io_outs_3(ces_18_21_io_outs_3)
  );
  Element ces_18_22 ( // @[MockArray.scala 36:52]
    .clock(ces_18_22_clock),
    .io_ins_0(ces_18_22_io_ins_0),
    .io_ins_1(ces_18_22_io_ins_1),
    .io_ins_2(ces_18_22_io_ins_2),
    .io_ins_3(ces_18_22_io_ins_3),
    .io_outs_0(ces_18_22_io_outs_0),
    .io_outs_1(ces_18_22_io_outs_1),
    .io_outs_2(ces_18_22_io_outs_2),
    .io_outs_3(ces_18_22_io_outs_3)
  );
  Element ces_18_23 ( // @[MockArray.scala 36:52]
    .clock(ces_18_23_clock),
    .io_ins_0(ces_18_23_io_ins_0),
    .io_ins_1(ces_18_23_io_ins_1),
    .io_ins_2(ces_18_23_io_ins_2),
    .io_ins_3(ces_18_23_io_ins_3),
    .io_outs_0(ces_18_23_io_outs_0),
    .io_outs_1(ces_18_23_io_outs_1),
    .io_outs_2(ces_18_23_io_outs_2),
    .io_outs_3(ces_18_23_io_outs_3)
  );
  Element ces_18_24 ( // @[MockArray.scala 36:52]
    .clock(ces_18_24_clock),
    .io_ins_0(ces_18_24_io_ins_0),
    .io_ins_1(ces_18_24_io_ins_1),
    .io_ins_2(ces_18_24_io_ins_2),
    .io_ins_3(ces_18_24_io_ins_3),
    .io_outs_0(ces_18_24_io_outs_0),
    .io_outs_1(ces_18_24_io_outs_1),
    .io_outs_2(ces_18_24_io_outs_2),
    .io_outs_3(ces_18_24_io_outs_3)
  );
  Element ces_18_25 ( // @[MockArray.scala 36:52]
    .clock(ces_18_25_clock),
    .io_ins_0(ces_18_25_io_ins_0),
    .io_ins_1(ces_18_25_io_ins_1),
    .io_ins_2(ces_18_25_io_ins_2),
    .io_ins_3(ces_18_25_io_ins_3),
    .io_outs_0(ces_18_25_io_outs_0),
    .io_outs_1(ces_18_25_io_outs_1),
    .io_outs_2(ces_18_25_io_outs_2),
    .io_outs_3(ces_18_25_io_outs_3)
  );
  Element ces_18_26 ( // @[MockArray.scala 36:52]
    .clock(ces_18_26_clock),
    .io_ins_0(ces_18_26_io_ins_0),
    .io_ins_1(ces_18_26_io_ins_1),
    .io_ins_2(ces_18_26_io_ins_2),
    .io_ins_3(ces_18_26_io_ins_3),
    .io_outs_0(ces_18_26_io_outs_0),
    .io_outs_1(ces_18_26_io_outs_1),
    .io_outs_2(ces_18_26_io_outs_2),
    .io_outs_3(ces_18_26_io_outs_3)
  );
  Element ces_18_27 ( // @[MockArray.scala 36:52]
    .clock(ces_18_27_clock),
    .io_ins_0(ces_18_27_io_ins_0),
    .io_ins_1(ces_18_27_io_ins_1),
    .io_ins_2(ces_18_27_io_ins_2),
    .io_ins_3(ces_18_27_io_ins_3),
    .io_outs_0(ces_18_27_io_outs_0),
    .io_outs_1(ces_18_27_io_outs_1),
    .io_outs_2(ces_18_27_io_outs_2),
    .io_outs_3(ces_18_27_io_outs_3)
  );
  Element ces_18_28 ( // @[MockArray.scala 36:52]
    .clock(ces_18_28_clock),
    .io_ins_0(ces_18_28_io_ins_0),
    .io_ins_1(ces_18_28_io_ins_1),
    .io_ins_2(ces_18_28_io_ins_2),
    .io_ins_3(ces_18_28_io_ins_3),
    .io_outs_0(ces_18_28_io_outs_0),
    .io_outs_1(ces_18_28_io_outs_1),
    .io_outs_2(ces_18_28_io_outs_2),
    .io_outs_3(ces_18_28_io_outs_3)
  );
  Element ces_18_29 ( // @[MockArray.scala 36:52]
    .clock(ces_18_29_clock),
    .io_ins_0(ces_18_29_io_ins_0),
    .io_ins_1(ces_18_29_io_ins_1),
    .io_ins_2(ces_18_29_io_ins_2),
    .io_ins_3(ces_18_29_io_ins_3),
    .io_outs_0(ces_18_29_io_outs_0),
    .io_outs_1(ces_18_29_io_outs_1),
    .io_outs_2(ces_18_29_io_outs_2),
    .io_outs_3(ces_18_29_io_outs_3)
  );
  Element ces_18_30 ( // @[MockArray.scala 36:52]
    .clock(ces_18_30_clock),
    .io_ins_0(ces_18_30_io_ins_0),
    .io_ins_1(ces_18_30_io_ins_1),
    .io_ins_2(ces_18_30_io_ins_2),
    .io_ins_3(ces_18_30_io_ins_3),
    .io_outs_0(ces_18_30_io_outs_0),
    .io_outs_1(ces_18_30_io_outs_1),
    .io_outs_2(ces_18_30_io_outs_2),
    .io_outs_3(ces_18_30_io_outs_3)
  );
  Element ces_18_31 ( // @[MockArray.scala 36:52]
    .clock(ces_18_31_clock),
    .io_ins_0(ces_18_31_io_ins_0),
    .io_ins_1(ces_18_31_io_ins_1),
    .io_ins_2(ces_18_31_io_ins_2),
    .io_ins_3(ces_18_31_io_ins_3),
    .io_outs_0(ces_18_31_io_outs_0),
    .io_outs_1(ces_18_31_io_outs_1),
    .io_outs_2(ces_18_31_io_outs_2),
    .io_outs_3(ces_18_31_io_outs_3)
  );
  Element ces_19_0 ( // @[MockArray.scala 36:52]
    .clock(ces_19_0_clock),
    .io_ins_0(ces_19_0_io_ins_0),
    .io_ins_1(ces_19_0_io_ins_1),
    .io_ins_2(ces_19_0_io_ins_2),
    .io_ins_3(ces_19_0_io_ins_3),
    .io_outs_0(ces_19_0_io_outs_0),
    .io_outs_1(ces_19_0_io_outs_1),
    .io_outs_2(ces_19_0_io_outs_2),
    .io_outs_3(ces_19_0_io_outs_3)
  );
  Element ces_19_1 ( // @[MockArray.scala 36:52]
    .clock(ces_19_1_clock),
    .io_ins_0(ces_19_1_io_ins_0),
    .io_ins_1(ces_19_1_io_ins_1),
    .io_ins_2(ces_19_1_io_ins_2),
    .io_ins_3(ces_19_1_io_ins_3),
    .io_outs_0(ces_19_1_io_outs_0),
    .io_outs_1(ces_19_1_io_outs_1),
    .io_outs_2(ces_19_1_io_outs_2),
    .io_outs_3(ces_19_1_io_outs_3)
  );
  Element ces_19_2 ( // @[MockArray.scala 36:52]
    .clock(ces_19_2_clock),
    .io_ins_0(ces_19_2_io_ins_0),
    .io_ins_1(ces_19_2_io_ins_1),
    .io_ins_2(ces_19_2_io_ins_2),
    .io_ins_3(ces_19_2_io_ins_3),
    .io_outs_0(ces_19_2_io_outs_0),
    .io_outs_1(ces_19_2_io_outs_1),
    .io_outs_2(ces_19_2_io_outs_2),
    .io_outs_3(ces_19_2_io_outs_3)
  );
  Element ces_19_3 ( // @[MockArray.scala 36:52]
    .clock(ces_19_3_clock),
    .io_ins_0(ces_19_3_io_ins_0),
    .io_ins_1(ces_19_3_io_ins_1),
    .io_ins_2(ces_19_3_io_ins_2),
    .io_ins_3(ces_19_3_io_ins_3),
    .io_outs_0(ces_19_3_io_outs_0),
    .io_outs_1(ces_19_3_io_outs_1),
    .io_outs_2(ces_19_3_io_outs_2),
    .io_outs_3(ces_19_3_io_outs_3)
  );
  Element ces_19_4 ( // @[MockArray.scala 36:52]
    .clock(ces_19_4_clock),
    .io_ins_0(ces_19_4_io_ins_0),
    .io_ins_1(ces_19_4_io_ins_1),
    .io_ins_2(ces_19_4_io_ins_2),
    .io_ins_3(ces_19_4_io_ins_3),
    .io_outs_0(ces_19_4_io_outs_0),
    .io_outs_1(ces_19_4_io_outs_1),
    .io_outs_2(ces_19_4_io_outs_2),
    .io_outs_3(ces_19_4_io_outs_3)
  );
  Element ces_19_5 ( // @[MockArray.scala 36:52]
    .clock(ces_19_5_clock),
    .io_ins_0(ces_19_5_io_ins_0),
    .io_ins_1(ces_19_5_io_ins_1),
    .io_ins_2(ces_19_5_io_ins_2),
    .io_ins_3(ces_19_5_io_ins_3),
    .io_outs_0(ces_19_5_io_outs_0),
    .io_outs_1(ces_19_5_io_outs_1),
    .io_outs_2(ces_19_5_io_outs_2),
    .io_outs_3(ces_19_5_io_outs_3)
  );
  Element ces_19_6 ( // @[MockArray.scala 36:52]
    .clock(ces_19_6_clock),
    .io_ins_0(ces_19_6_io_ins_0),
    .io_ins_1(ces_19_6_io_ins_1),
    .io_ins_2(ces_19_6_io_ins_2),
    .io_ins_3(ces_19_6_io_ins_3),
    .io_outs_0(ces_19_6_io_outs_0),
    .io_outs_1(ces_19_6_io_outs_1),
    .io_outs_2(ces_19_6_io_outs_2),
    .io_outs_3(ces_19_6_io_outs_3)
  );
  Element ces_19_7 ( // @[MockArray.scala 36:52]
    .clock(ces_19_7_clock),
    .io_ins_0(ces_19_7_io_ins_0),
    .io_ins_1(ces_19_7_io_ins_1),
    .io_ins_2(ces_19_7_io_ins_2),
    .io_ins_3(ces_19_7_io_ins_3),
    .io_outs_0(ces_19_7_io_outs_0),
    .io_outs_1(ces_19_7_io_outs_1),
    .io_outs_2(ces_19_7_io_outs_2),
    .io_outs_3(ces_19_7_io_outs_3)
  );
  Element ces_19_8 ( // @[MockArray.scala 36:52]
    .clock(ces_19_8_clock),
    .io_ins_0(ces_19_8_io_ins_0),
    .io_ins_1(ces_19_8_io_ins_1),
    .io_ins_2(ces_19_8_io_ins_2),
    .io_ins_3(ces_19_8_io_ins_3),
    .io_outs_0(ces_19_8_io_outs_0),
    .io_outs_1(ces_19_8_io_outs_1),
    .io_outs_2(ces_19_8_io_outs_2),
    .io_outs_3(ces_19_8_io_outs_3)
  );
  Element ces_19_9 ( // @[MockArray.scala 36:52]
    .clock(ces_19_9_clock),
    .io_ins_0(ces_19_9_io_ins_0),
    .io_ins_1(ces_19_9_io_ins_1),
    .io_ins_2(ces_19_9_io_ins_2),
    .io_ins_3(ces_19_9_io_ins_3),
    .io_outs_0(ces_19_9_io_outs_0),
    .io_outs_1(ces_19_9_io_outs_1),
    .io_outs_2(ces_19_9_io_outs_2),
    .io_outs_3(ces_19_9_io_outs_3)
  );
  Element ces_19_10 ( // @[MockArray.scala 36:52]
    .clock(ces_19_10_clock),
    .io_ins_0(ces_19_10_io_ins_0),
    .io_ins_1(ces_19_10_io_ins_1),
    .io_ins_2(ces_19_10_io_ins_2),
    .io_ins_3(ces_19_10_io_ins_3),
    .io_outs_0(ces_19_10_io_outs_0),
    .io_outs_1(ces_19_10_io_outs_1),
    .io_outs_2(ces_19_10_io_outs_2),
    .io_outs_3(ces_19_10_io_outs_3)
  );
  Element ces_19_11 ( // @[MockArray.scala 36:52]
    .clock(ces_19_11_clock),
    .io_ins_0(ces_19_11_io_ins_0),
    .io_ins_1(ces_19_11_io_ins_1),
    .io_ins_2(ces_19_11_io_ins_2),
    .io_ins_3(ces_19_11_io_ins_3),
    .io_outs_0(ces_19_11_io_outs_0),
    .io_outs_1(ces_19_11_io_outs_1),
    .io_outs_2(ces_19_11_io_outs_2),
    .io_outs_3(ces_19_11_io_outs_3)
  );
  Element ces_19_12 ( // @[MockArray.scala 36:52]
    .clock(ces_19_12_clock),
    .io_ins_0(ces_19_12_io_ins_0),
    .io_ins_1(ces_19_12_io_ins_1),
    .io_ins_2(ces_19_12_io_ins_2),
    .io_ins_3(ces_19_12_io_ins_3),
    .io_outs_0(ces_19_12_io_outs_0),
    .io_outs_1(ces_19_12_io_outs_1),
    .io_outs_2(ces_19_12_io_outs_2),
    .io_outs_3(ces_19_12_io_outs_3)
  );
  Element ces_19_13 ( // @[MockArray.scala 36:52]
    .clock(ces_19_13_clock),
    .io_ins_0(ces_19_13_io_ins_0),
    .io_ins_1(ces_19_13_io_ins_1),
    .io_ins_2(ces_19_13_io_ins_2),
    .io_ins_3(ces_19_13_io_ins_3),
    .io_outs_0(ces_19_13_io_outs_0),
    .io_outs_1(ces_19_13_io_outs_1),
    .io_outs_2(ces_19_13_io_outs_2),
    .io_outs_3(ces_19_13_io_outs_3)
  );
  Element ces_19_14 ( // @[MockArray.scala 36:52]
    .clock(ces_19_14_clock),
    .io_ins_0(ces_19_14_io_ins_0),
    .io_ins_1(ces_19_14_io_ins_1),
    .io_ins_2(ces_19_14_io_ins_2),
    .io_ins_3(ces_19_14_io_ins_3),
    .io_outs_0(ces_19_14_io_outs_0),
    .io_outs_1(ces_19_14_io_outs_1),
    .io_outs_2(ces_19_14_io_outs_2),
    .io_outs_3(ces_19_14_io_outs_3)
  );
  Element ces_19_15 ( // @[MockArray.scala 36:52]
    .clock(ces_19_15_clock),
    .io_ins_0(ces_19_15_io_ins_0),
    .io_ins_1(ces_19_15_io_ins_1),
    .io_ins_2(ces_19_15_io_ins_2),
    .io_ins_3(ces_19_15_io_ins_3),
    .io_outs_0(ces_19_15_io_outs_0),
    .io_outs_1(ces_19_15_io_outs_1),
    .io_outs_2(ces_19_15_io_outs_2),
    .io_outs_3(ces_19_15_io_outs_3)
  );
  Element ces_19_16 ( // @[MockArray.scala 36:52]
    .clock(ces_19_16_clock),
    .io_ins_0(ces_19_16_io_ins_0),
    .io_ins_1(ces_19_16_io_ins_1),
    .io_ins_2(ces_19_16_io_ins_2),
    .io_ins_3(ces_19_16_io_ins_3),
    .io_outs_0(ces_19_16_io_outs_0),
    .io_outs_1(ces_19_16_io_outs_1),
    .io_outs_2(ces_19_16_io_outs_2),
    .io_outs_3(ces_19_16_io_outs_3)
  );
  Element ces_19_17 ( // @[MockArray.scala 36:52]
    .clock(ces_19_17_clock),
    .io_ins_0(ces_19_17_io_ins_0),
    .io_ins_1(ces_19_17_io_ins_1),
    .io_ins_2(ces_19_17_io_ins_2),
    .io_ins_3(ces_19_17_io_ins_3),
    .io_outs_0(ces_19_17_io_outs_0),
    .io_outs_1(ces_19_17_io_outs_1),
    .io_outs_2(ces_19_17_io_outs_2),
    .io_outs_3(ces_19_17_io_outs_3)
  );
  Element ces_19_18 ( // @[MockArray.scala 36:52]
    .clock(ces_19_18_clock),
    .io_ins_0(ces_19_18_io_ins_0),
    .io_ins_1(ces_19_18_io_ins_1),
    .io_ins_2(ces_19_18_io_ins_2),
    .io_ins_3(ces_19_18_io_ins_3),
    .io_outs_0(ces_19_18_io_outs_0),
    .io_outs_1(ces_19_18_io_outs_1),
    .io_outs_2(ces_19_18_io_outs_2),
    .io_outs_3(ces_19_18_io_outs_3)
  );
  Element ces_19_19 ( // @[MockArray.scala 36:52]
    .clock(ces_19_19_clock),
    .io_ins_0(ces_19_19_io_ins_0),
    .io_ins_1(ces_19_19_io_ins_1),
    .io_ins_2(ces_19_19_io_ins_2),
    .io_ins_3(ces_19_19_io_ins_3),
    .io_outs_0(ces_19_19_io_outs_0),
    .io_outs_1(ces_19_19_io_outs_1),
    .io_outs_2(ces_19_19_io_outs_2),
    .io_outs_3(ces_19_19_io_outs_3)
  );
  Element ces_19_20 ( // @[MockArray.scala 36:52]
    .clock(ces_19_20_clock),
    .io_ins_0(ces_19_20_io_ins_0),
    .io_ins_1(ces_19_20_io_ins_1),
    .io_ins_2(ces_19_20_io_ins_2),
    .io_ins_3(ces_19_20_io_ins_3),
    .io_outs_0(ces_19_20_io_outs_0),
    .io_outs_1(ces_19_20_io_outs_1),
    .io_outs_2(ces_19_20_io_outs_2),
    .io_outs_3(ces_19_20_io_outs_3)
  );
  Element ces_19_21 ( // @[MockArray.scala 36:52]
    .clock(ces_19_21_clock),
    .io_ins_0(ces_19_21_io_ins_0),
    .io_ins_1(ces_19_21_io_ins_1),
    .io_ins_2(ces_19_21_io_ins_2),
    .io_ins_3(ces_19_21_io_ins_3),
    .io_outs_0(ces_19_21_io_outs_0),
    .io_outs_1(ces_19_21_io_outs_1),
    .io_outs_2(ces_19_21_io_outs_2),
    .io_outs_3(ces_19_21_io_outs_3)
  );
  Element ces_19_22 ( // @[MockArray.scala 36:52]
    .clock(ces_19_22_clock),
    .io_ins_0(ces_19_22_io_ins_0),
    .io_ins_1(ces_19_22_io_ins_1),
    .io_ins_2(ces_19_22_io_ins_2),
    .io_ins_3(ces_19_22_io_ins_3),
    .io_outs_0(ces_19_22_io_outs_0),
    .io_outs_1(ces_19_22_io_outs_1),
    .io_outs_2(ces_19_22_io_outs_2),
    .io_outs_3(ces_19_22_io_outs_3)
  );
  Element ces_19_23 ( // @[MockArray.scala 36:52]
    .clock(ces_19_23_clock),
    .io_ins_0(ces_19_23_io_ins_0),
    .io_ins_1(ces_19_23_io_ins_1),
    .io_ins_2(ces_19_23_io_ins_2),
    .io_ins_3(ces_19_23_io_ins_3),
    .io_outs_0(ces_19_23_io_outs_0),
    .io_outs_1(ces_19_23_io_outs_1),
    .io_outs_2(ces_19_23_io_outs_2),
    .io_outs_3(ces_19_23_io_outs_3)
  );
  Element ces_19_24 ( // @[MockArray.scala 36:52]
    .clock(ces_19_24_clock),
    .io_ins_0(ces_19_24_io_ins_0),
    .io_ins_1(ces_19_24_io_ins_1),
    .io_ins_2(ces_19_24_io_ins_2),
    .io_ins_3(ces_19_24_io_ins_3),
    .io_outs_0(ces_19_24_io_outs_0),
    .io_outs_1(ces_19_24_io_outs_1),
    .io_outs_2(ces_19_24_io_outs_2),
    .io_outs_3(ces_19_24_io_outs_3)
  );
  Element ces_19_25 ( // @[MockArray.scala 36:52]
    .clock(ces_19_25_clock),
    .io_ins_0(ces_19_25_io_ins_0),
    .io_ins_1(ces_19_25_io_ins_1),
    .io_ins_2(ces_19_25_io_ins_2),
    .io_ins_3(ces_19_25_io_ins_3),
    .io_outs_0(ces_19_25_io_outs_0),
    .io_outs_1(ces_19_25_io_outs_1),
    .io_outs_2(ces_19_25_io_outs_2),
    .io_outs_3(ces_19_25_io_outs_3)
  );
  Element ces_19_26 ( // @[MockArray.scala 36:52]
    .clock(ces_19_26_clock),
    .io_ins_0(ces_19_26_io_ins_0),
    .io_ins_1(ces_19_26_io_ins_1),
    .io_ins_2(ces_19_26_io_ins_2),
    .io_ins_3(ces_19_26_io_ins_3),
    .io_outs_0(ces_19_26_io_outs_0),
    .io_outs_1(ces_19_26_io_outs_1),
    .io_outs_2(ces_19_26_io_outs_2),
    .io_outs_3(ces_19_26_io_outs_3)
  );
  Element ces_19_27 ( // @[MockArray.scala 36:52]
    .clock(ces_19_27_clock),
    .io_ins_0(ces_19_27_io_ins_0),
    .io_ins_1(ces_19_27_io_ins_1),
    .io_ins_2(ces_19_27_io_ins_2),
    .io_ins_3(ces_19_27_io_ins_3),
    .io_outs_0(ces_19_27_io_outs_0),
    .io_outs_1(ces_19_27_io_outs_1),
    .io_outs_2(ces_19_27_io_outs_2),
    .io_outs_3(ces_19_27_io_outs_3)
  );
  Element ces_19_28 ( // @[MockArray.scala 36:52]
    .clock(ces_19_28_clock),
    .io_ins_0(ces_19_28_io_ins_0),
    .io_ins_1(ces_19_28_io_ins_1),
    .io_ins_2(ces_19_28_io_ins_2),
    .io_ins_3(ces_19_28_io_ins_3),
    .io_outs_0(ces_19_28_io_outs_0),
    .io_outs_1(ces_19_28_io_outs_1),
    .io_outs_2(ces_19_28_io_outs_2),
    .io_outs_3(ces_19_28_io_outs_3)
  );
  Element ces_19_29 ( // @[MockArray.scala 36:52]
    .clock(ces_19_29_clock),
    .io_ins_0(ces_19_29_io_ins_0),
    .io_ins_1(ces_19_29_io_ins_1),
    .io_ins_2(ces_19_29_io_ins_2),
    .io_ins_3(ces_19_29_io_ins_3),
    .io_outs_0(ces_19_29_io_outs_0),
    .io_outs_1(ces_19_29_io_outs_1),
    .io_outs_2(ces_19_29_io_outs_2),
    .io_outs_3(ces_19_29_io_outs_3)
  );
  Element ces_19_30 ( // @[MockArray.scala 36:52]
    .clock(ces_19_30_clock),
    .io_ins_0(ces_19_30_io_ins_0),
    .io_ins_1(ces_19_30_io_ins_1),
    .io_ins_2(ces_19_30_io_ins_2),
    .io_ins_3(ces_19_30_io_ins_3),
    .io_outs_0(ces_19_30_io_outs_0),
    .io_outs_1(ces_19_30_io_outs_1),
    .io_outs_2(ces_19_30_io_outs_2),
    .io_outs_3(ces_19_30_io_outs_3)
  );
  Element ces_19_31 ( // @[MockArray.scala 36:52]
    .clock(ces_19_31_clock),
    .io_ins_0(ces_19_31_io_ins_0),
    .io_ins_1(ces_19_31_io_ins_1),
    .io_ins_2(ces_19_31_io_ins_2),
    .io_ins_3(ces_19_31_io_ins_3),
    .io_outs_0(ces_19_31_io_outs_0),
    .io_outs_1(ces_19_31_io_outs_1),
    .io_outs_2(ces_19_31_io_outs_2),
    .io_outs_3(ces_19_31_io_outs_3)
  );
  Element ces_20_0 ( // @[MockArray.scala 36:52]
    .clock(ces_20_0_clock),
    .io_ins_0(ces_20_0_io_ins_0),
    .io_ins_1(ces_20_0_io_ins_1),
    .io_ins_2(ces_20_0_io_ins_2),
    .io_ins_3(ces_20_0_io_ins_3),
    .io_outs_0(ces_20_0_io_outs_0),
    .io_outs_1(ces_20_0_io_outs_1),
    .io_outs_2(ces_20_0_io_outs_2),
    .io_outs_3(ces_20_0_io_outs_3)
  );
  Element ces_20_1 ( // @[MockArray.scala 36:52]
    .clock(ces_20_1_clock),
    .io_ins_0(ces_20_1_io_ins_0),
    .io_ins_1(ces_20_1_io_ins_1),
    .io_ins_2(ces_20_1_io_ins_2),
    .io_ins_3(ces_20_1_io_ins_3),
    .io_outs_0(ces_20_1_io_outs_0),
    .io_outs_1(ces_20_1_io_outs_1),
    .io_outs_2(ces_20_1_io_outs_2),
    .io_outs_3(ces_20_1_io_outs_3)
  );
  Element ces_20_2 ( // @[MockArray.scala 36:52]
    .clock(ces_20_2_clock),
    .io_ins_0(ces_20_2_io_ins_0),
    .io_ins_1(ces_20_2_io_ins_1),
    .io_ins_2(ces_20_2_io_ins_2),
    .io_ins_3(ces_20_2_io_ins_3),
    .io_outs_0(ces_20_2_io_outs_0),
    .io_outs_1(ces_20_2_io_outs_1),
    .io_outs_2(ces_20_2_io_outs_2),
    .io_outs_3(ces_20_2_io_outs_3)
  );
  Element ces_20_3 ( // @[MockArray.scala 36:52]
    .clock(ces_20_3_clock),
    .io_ins_0(ces_20_3_io_ins_0),
    .io_ins_1(ces_20_3_io_ins_1),
    .io_ins_2(ces_20_3_io_ins_2),
    .io_ins_3(ces_20_3_io_ins_3),
    .io_outs_0(ces_20_3_io_outs_0),
    .io_outs_1(ces_20_3_io_outs_1),
    .io_outs_2(ces_20_3_io_outs_2),
    .io_outs_3(ces_20_3_io_outs_3)
  );
  Element ces_20_4 ( // @[MockArray.scala 36:52]
    .clock(ces_20_4_clock),
    .io_ins_0(ces_20_4_io_ins_0),
    .io_ins_1(ces_20_4_io_ins_1),
    .io_ins_2(ces_20_4_io_ins_2),
    .io_ins_3(ces_20_4_io_ins_3),
    .io_outs_0(ces_20_4_io_outs_0),
    .io_outs_1(ces_20_4_io_outs_1),
    .io_outs_2(ces_20_4_io_outs_2),
    .io_outs_3(ces_20_4_io_outs_3)
  );
  Element ces_20_5 ( // @[MockArray.scala 36:52]
    .clock(ces_20_5_clock),
    .io_ins_0(ces_20_5_io_ins_0),
    .io_ins_1(ces_20_5_io_ins_1),
    .io_ins_2(ces_20_5_io_ins_2),
    .io_ins_3(ces_20_5_io_ins_3),
    .io_outs_0(ces_20_5_io_outs_0),
    .io_outs_1(ces_20_5_io_outs_1),
    .io_outs_2(ces_20_5_io_outs_2),
    .io_outs_3(ces_20_5_io_outs_3)
  );
  Element ces_20_6 ( // @[MockArray.scala 36:52]
    .clock(ces_20_6_clock),
    .io_ins_0(ces_20_6_io_ins_0),
    .io_ins_1(ces_20_6_io_ins_1),
    .io_ins_2(ces_20_6_io_ins_2),
    .io_ins_3(ces_20_6_io_ins_3),
    .io_outs_0(ces_20_6_io_outs_0),
    .io_outs_1(ces_20_6_io_outs_1),
    .io_outs_2(ces_20_6_io_outs_2),
    .io_outs_3(ces_20_6_io_outs_3)
  );
  Element ces_20_7 ( // @[MockArray.scala 36:52]
    .clock(ces_20_7_clock),
    .io_ins_0(ces_20_7_io_ins_0),
    .io_ins_1(ces_20_7_io_ins_1),
    .io_ins_2(ces_20_7_io_ins_2),
    .io_ins_3(ces_20_7_io_ins_3),
    .io_outs_0(ces_20_7_io_outs_0),
    .io_outs_1(ces_20_7_io_outs_1),
    .io_outs_2(ces_20_7_io_outs_2),
    .io_outs_3(ces_20_7_io_outs_3)
  );
  Element ces_20_8 ( // @[MockArray.scala 36:52]
    .clock(ces_20_8_clock),
    .io_ins_0(ces_20_8_io_ins_0),
    .io_ins_1(ces_20_8_io_ins_1),
    .io_ins_2(ces_20_8_io_ins_2),
    .io_ins_3(ces_20_8_io_ins_3),
    .io_outs_0(ces_20_8_io_outs_0),
    .io_outs_1(ces_20_8_io_outs_1),
    .io_outs_2(ces_20_8_io_outs_2),
    .io_outs_3(ces_20_8_io_outs_3)
  );
  Element ces_20_9 ( // @[MockArray.scala 36:52]
    .clock(ces_20_9_clock),
    .io_ins_0(ces_20_9_io_ins_0),
    .io_ins_1(ces_20_9_io_ins_1),
    .io_ins_2(ces_20_9_io_ins_2),
    .io_ins_3(ces_20_9_io_ins_3),
    .io_outs_0(ces_20_9_io_outs_0),
    .io_outs_1(ces_20_9_io_outs_1),
    .io_outs_2(ces_20_9_io_outs_2),
    .io_outs_3(ces_20_9_io_outs_3)
  );
  Element ces_20_10 ( // @[MockArray.scala 36:52]
    .clock(ces_20_10_clock),
    .io_ins_0(ces_20_10_io_ins_0),
    .io_ins_1(ces_20_10_io_ins_1),
    .io_ins_2(ces_20_10_io_ins_2),
    .io_ins_3(ces_20_10_io_ins_3),
    .io_outs_0(ces_20_10_io_outs_0),
    .io_outs_1(ces_20_10_io_outs_1),
    .io_outs_2(ces_20_10_io_outs_2),
    .io_outs_3(ces_20_10_io_outs_3)
  );
  Element ces_20_11 ( // @[MockArray.scala 36:52]
    .clock(ces_20_11_clock),
    .io_ins_0(ces_20_11_io_ins_0),
    .io_ins_1(ces_20_11_io_ins_1),
    .io_ins_2(ces_20_11_io_ins_2),
    .io_ins_3(ces_20_11_io_ins_3),
    .io_outs_0(ces_20_11_io_outs_0),
    .io_outs_1(ces_20_11_io_outs_1),
    .io_outs_2(ces_20_11_io_outs_2),
    .io_outs_3(ces_20_11_io_outs_3)
  );
  Element ces_20_12 ( // @[MockArray.scala 36:52]
    .clock(ces_20_12_clock),
    .io_ins_0(ces_20_12_io_ins_0),
    .io_ins_1(ces_20_12_io_ins_1),
    .io_ins_2(ces_20_12_io_ins_2),
    .io_ins_3(ces_20_12_io_ins_3),
    .io_outs_0(ces_20_12_io_outs_0),
    .io_outs_1(ces_20_12_io_outs_1),
    .io_outs_2(ces_20_12_io_outs_2),
    .io_outs_3(ces_20_12_io_outs_3)
  );
  Element ces_20_13 ( // @[MockArray.scala 36:52]
    .clock(ces_20_13_clock),
    .io_ins_0(ces_20_13_io_ins_0),
    .io_ins_1(ces_20_13_io_ins_1),
    .io_ins_2(ces_20_13_io_ins_2),
    .io_ins_3(ces_20_13_io_ins_3),
    .io_outs_0(ces_20_13_io_outs_0),
    .io_outs_1(ces_20_13_io_outs_1),
    .io_outs_2(ces_20_13_io_outs_2),
    .io_outs_3(ces_20_13_io_outs_3)
  );
  Element ces_20_14 ( // @[MockArray.scala 36:52]
    .clock(ces_20_14_clock),
    .io_ins_0(ces_20_14_io_ins_0),
    .io_ins_1(ces_20_14_io_ins_1),
    .io_ins_2(ces_20_14_io_ins_2),
    .io_ins_3(ces_20_14_io_ins_3),
    .io_outs_0(ces_20_14_io_outs_0),
    .io_outs_1(ces_20_14_io_outs_1),
    .io_outs_2(ces_20_14_io_outs_2),
    .io_outs_3(ces_20_14_io_outs_3)
  );
  Element ces_20_15 ( // @[MockArray.scala 36:52]
    .clock(ces_20_15_clock),
    .io_ins_0(ces_20_15_io_ins_0),
    .io_ins_1(ces_20_15_io_ins_1),
    .io_ins_2(ces_20_15_io_ins_2),
    .io_ins_3(ces_20_15_io_ins_3),
    .io_outs_0(ces_20_15_io_outs_0),
    .io_outs_1(ces_20_15_io_outs_1),
    .io_outs_2(ces_20_15_io_outs_2),
    .io_outs_3(ces_20_15_io_outs_3)
  );
  Element ces_20_16 ( // @[MockArray.scala 36:52]
    .clock(ces_20_16_clock),
    .io_ins_0(ces_20_16_io_ins_0),
    .io_ins_1(ces_20_16_io_ins_1),
    .io_ins_2(ces_20_16_io_ins_2),
    .io_ins_3(ces_20_16_io_ins_3),
    .io_outs_0(ces_20_16_io_outs_0),
    .io_outs_1(ces_20_16_io_outs_1),
    .io_outs_2(ces_20_16_io_outs_2),
    .io_outs_3(ces_20_16_io_outs_3)
  );
  Element ces_20_17 ( // @[MockArray.scala 36:52]
    .clock(ces_20_17_clock),
    .io_ins_0(ces_20_17_io_ins_0),
    .io_ins_1(ces_20_17_io_ins_1),
    .io_ins_2(ces_20_17_io_ins_2),
    .io_ins_3(ces_20_17_io_ins_3),
    .io_outs_0(ces_20_17_io_outs_0),
    .io_outs_1(ces_20_17_io_outs_1),
    .io_outs_2(ces_20_17_io_outs_2),
    .io_outs_3(ces_20_17_io_outs_3)
  );
  Element ces_20_18 ( // @[MockArray.scala 36:52]
    .clock(ces_20_18_clock),
    .io_ins_0(ces_20_18_io_ins_0),
    .io_ins_1(ces_20_18_io_ins_1),
    .io_ins_2(ces_20_18_io_ins_2),
    .io_ins_3(ces_20_18_io_ins_3),
    .io_outs_0(ces_20_18_io_outs_0),
    .io_outs_1(ces_20_18_io_outs_1),
    .io_outs_2(ces_20_18_io_outs_2),
    .io_outs_3(ces_20_18_io_outs_3)
  );
  Element ces_20_19 ( // @[MockArray.scala 36:52]
    .clock(ces_20_19_clock),
    .io_ins_0(ces_20_19_io_ins_0),
    .io_ins_1(ces_20_19_io_ins_1),
    .io_ins_2(ces_20_19_io_ins_2),
    .io_ins_3(ces_20_19_io_ins_3),
    .io_outs_0(ces_20_19_io_outs_0),
    .io_outs_1(ces_20_19_io_outs_1),
    .io_outs_2(ces_20_19_io_outs_2),
    .io_outs_3(ces_20_19_io_outs_3)
  );
  Element ces_20_20 ( // @[MockArray.scala 36:52]
    .clock(ces_20_20_clock),
    .io_ins_0(ces_20_20_io_ins_0),
    .io_ins_1(ces_20_20_io_ins_1),
    .io_ins_2(ces_20_20_io_ins_2),
    .io_ins_3(ces_20_20_io_ins_3),
    .io_outs_0(ces_20_20_io_outs_0),
    .io_outs_1(ces_20_20_io_outs_1),
    .io_outs_2(ces_20_20_io_outs_2),
    .io_outs_3(ces_20_20_io_outs_3)
  );
  Element ces_20_21 ( // @[MockArray.scala 36:52]
    .clock(ces_20_21_clock),
    .io_ins_0(ces_20_21_io_ins_0),
    .io_ins_1(ces_20_21_io_ins_1),
    .io_ins_2(ces_20_21_io_ins_2),
    .io_ins_3(ces_20_21_io_ins_3),
    .io_outs_0(ces_20_21_io_outs_0),
    .io_outs_1(ces_20_21_io_outs_1),
    .io_outs_2(ces_20_21_io_outs_2),
    .io_outs_3(ces_20_21_io_outs_3)
  );
  Element ces_20_22 ( // @[MockArray.scala 36:52]
    .clock(ces_20_22_clock),
    .io_ins_0(ces_20_22_io_ins_0),
    .io_ins_1(ces_20_22_io_ins_1),
    .io_ins_2(ces_20_22_io_ins_2),
    .io_ins_3(ces_20_22_io_ins_3),
    .io_outs_0(ces_20_22_io_outs_0),
    .io_outs_1(ces_20_22_io_outs_1),
    .io_outs_2(ces_20_22_io_outs_2),
    .io_outs_3(ces_20_22_io_outs_3)
  );
  Element ces_20_23 ( // @[MockArray.scala 36:52]
    .clock(ces_20_23_clock),
    .io_ins_0(ces_20_23_io_ins_0),
    .io_ins_1(ces_20_23_io_ins_1),
    .io_ins_2(ces_20_23_io_ins_2),
    .io_ins_3(ces_20_23_io_ins_3),
    .io_outs_0(ces_20_23_io_outs_0),
    .io_outs_1(ces_20_23_io_outs_1),
    .io_outs_2(ces_20_23_io_outs_2),
    .io_outs_3(ces_20_23_io_outs_3)
  );
  Element ces_20_24 ( // @[MockArray.scala 36:52]
    .clock(ces_20_24_clock),
    .io_ins_0(ces_20_24_io_ins_0),
    .io_ins_1(ces_20_24_io_ins_1),
    .io_ins_2(ces_20_24_io_ins_2),
    .io_ins_3(ces_20_24_io_ins_3),
    .io_outs_0(ces_20_24_io_outs_0),
    .io_outs_1(ces_20_24_io_outs_1),
    .io_outs_2(ces_20_24_io_outs_2),
    .io_outs_3(ces_20_24_io_outs_3)
  );
  Element ces_20_25 ( // @[MockArray.scala 36:52]
    .clock(ces_20_25_clock),
    .io_ins_0(ces_20_25_io_ins_0),
    .io_ins_1(ces_20_25_io_ins_1),
    .io_ins_2(ces_20_25_io_ins_2),
    .io_ins_3(ces_20_25_io_ins_3),
    .io_outs_0(ces_20_25_io_outs_0),
    .io_outs_1(ces_20_25_io_outs_1),
    .io_outs_2(ces_20_25_io_outs_2),
    .io_outs_3(ces_20_25_io_outs_3)
  );
  Element ces_20_26 ( // @[MockArray.scala 36:52]
    .clock(ces_20_26_clock),
    .io_ins_0(ces_20_26_io_ins_0),
    .io_ins_1(ces_20_26_io_ins_1),
    .io_ins_2(ces_20_26_io_ins_2),
    .io_ins_3(ces_20_26_io_ins_3),
    .io_outs_0(ces_20_26_io_outs_0),
    .io_outs_1(ces_20_26_io_outs_1),
    .io_outs_2(ces_20_26_io_outs_2),
    .io_outs_3(ces_20_26_io_outs_3)
  );
  Element ces_20_27 ( // @[MockArray.scala 36:52]
    .clock(ces_20_27_clock),
    .io_ins_0(ces_20_27_io_ins_0),
    .io_ins_1(ces_20_27_io_ins_1),
    .io_ins_2(ces_20_27_io_ins_2),
    .io_ins_3(ces_20_27_io_ins_3),
    .io_outs_0(ces_20_27_io_outs_0),
    .io_outs_1(ces_20_27_io_outs_1),
    .io_outs_2(ces_20_27_io_outs_2),
    .io_outs_3(ces_20_27_io_outs_3)
  );
  Element ces_20_28 ( // @[MockArray.scala 36:52]
    .clock(ces_20_28_clock),
    .io_ins_0(ces_20_28_io_ins_0),
    .io_ins_1(ces_20_28_io_ins_1),
    .io_ins_2(ces_20_28_io_ins_2),
    .io_ins_3(ces_20_28_io_ins_3),
    .io_outs_0(ces_20_28_io_outs_0),
    .io_outs_1(ces_20_28_io_outs_1),
    .io_outs_2(ces_20_28_io_outs_2),
    .io_outs_3(ces_20_28_io_outs_3)
  );
  Element ces_20_29 ( // @[MockArray.scala 36:52]
    .clock(ces_20_29_clock),
    .io_ins_0(ces_20_29_io_ins_0),
    .io_ins_1(ces_20_29_io_ins_1),
    .io_ins_2(ces_20_29_io_ins_2),
    .io_ins_3(ces_20_29_io_ins_3),
    .io_outs_0(ces_20_29_io_outs_0),
    .io_outs_1(ces_20_29_io_outs_1),
    .io_outs_2(ces_20_29_io_outs_2),
    .io_outs_3(ces_20_29_io_outs_3)
  );
  Element ces_20_30 ( // @[MockArray.scala 36:52]
    .clock(ces_20_30_clock),
    .io_ins_0(ces_20_30_io_ins_0),
    .io_ins_1(ces_20_30_io_ins_1),
    .io_ins_2(ces_20_30_io_ins_2),
    .io_ins_3(ces_20_30_io_ins_3),
    .io_outs_0(ces_20_30_io_outs_0),
    .io_outs_1(ces_20_30_io_outs_1),
    .io_outs_2(ces_20_30_io_outs_2),
    .io_outs_3(ces_20_30_io_outs_3)
  );
  Element ces_20_31 ( // @[MockArray.scala 36:52]
    .clock(ces_20_31_clock),
    .io_ins_0(ces_20_31_io_ins_0),
    .io_ins_1(ces_20_31_io_ins_1),
    .io_ins_2(ces_20_31_io_ins_2),
    .io_ins_3(ces_20_31_io_ins_3),
    .io_outs_0(ces_20_31_io_outs_0),
    .io_outs_1(ces_20_31_io_outs_1),
    .io_outs_2(ces_20_31_io_outs_2),
    .io_outs_3(ces_20_31_io_outs_3)
  );
  Element ces_21_0 ( // @[MockArray.scala 36:52]
    .clock(ces_21_0_clock),
    .io_ins_0(ces_21_0_io_ins_0),
    .io_ins_1(ces_21_0_io_ins_1),
    .io_ins_2(ces_21_0_io_ins_2),
    .io_ins_3(ces_21_0_io_ins_3),
    .io_outs_0(ces_21_0_io_outs_0),
    .io_outs_1(ces_21_0_io_outs_1),
    .io_outs_2(ces_21_0_io_outs_2),
    .io_outs_3(ces_21_0_io_outs_3)
  );
  Element ces_21_1 ( // @[MockArray.scala 36:52]
    .clock(ces_21_1_clock),
    .io_ins_0(ces_21_1_io_ins_0),
    .io_ins_1(ces_21_1_io_ins_1),
    .io_ins_2(ces_21_1_io_ins_2),
    .io_ins_3(ces_21_1_io_ins_3),
    .io_outs_0(ces_21_1_io_outs_0),
    .io_outs_1(ces_21_1_io_outs_1),
    .io_outs_2(ces_21_1_io_outs_2),
    .io_outs_3(ces_21_1_io_outs_3)
  );
  Element ces_21_2 ( // @[MockArray.scala 36:52]
    .clock(ces_21_2_clock),
    .io_ins_0(ces_21_2_io_ins_0),
    .io_ins_1(ces_21_2_io_ins_1),
    .io_ins_2(ces_21_2_io_ins_2),
    .io_ins_3(ces_21_2_io_ins_3),
    .io_outs_0(ces_21_2_io_outs_0),
    .io_outs_1(ces_21_2_io_outs_1),
    .io_outs_2(ces_21_2_io_outs_2),
    .io_outs_3(ces_21_2_io_outs_3)
  );
  Element ces_21_3 ( // @[MockArray.scala 36:52]
    .clock(ces_21_3_clock),
    .io_ins_0(ces_21_3_io_ins_0),
    .io_ins_1(ces_21_3_io_ins_1),
    .io_ins_2(ces_21_3_io_ins_2),
    .io_ins_3(ces_21_3_io_ins_3),
    .io_outs_0(ces_21_3_io_outs_0),
    .io_outs_1(ces_21_3_io_outs_1),
    .io_outs_2(ces_21_3_io_outs_2),
    .io_outs_3(ces_21_3_io_outs_3)
  );
  Element ces_21_4 ( // @[MockArray.scala 36:52]
    .clock(ces_21_4_clock),
    .io_ins_0(ces_21_4_io_ins_0),
    .io_ins_1(ces_21_4_io_ins_1),
    .io_ins_2(ces_21_4_io_ins_2),
    .io_ins_3(ces_21_4_io_ins_3),
    .io_outs_0(ces_21_4_io_outs_0),
    .io_outs_1(ces_21_4_io_outs_1),
    .io_outs_2(ces_21_4_io_outs_2),
    .io_outs_3(ces_21_4_io_outs_3)
  );
  Element ces_21_5 ( // @[MockArray.scala 36:52]
    .clock(ces_21_5_clock),
    .io_ins_0(ces_21_5_io_ins_0),
    .io_ins_1(ces_21_5_io_ins_1),
    .io_ins_2(ces_21_5_io_ins_2),
    .io_ins_3(ces_21_5_io_ins_3),
    .io_outs_0(ces_21_5_io_outs_0),
    .io_outs_1(ces_21_5_io_outs_1),
    .io_outs_2(ces_21_5_io_outs_2),
    .io_outs_3(ces_21_5_io_outs_3)
  );
  Element ces_21_6 ( // @[MockArray.scala 36:52]
    .clock(ces_21_6_clock),
    .io_ins_0(ces_21_6_io_ins_0),
    .io_ins_1(ces_21_6_io_ins_1),
    .io_ins_2(ces_21_6_io_ins_2),
    .io_ins_3(ces_21_6_io_ins_3),
    .io_outs_0(ces_21_6_io_outs_0),
    .io_outs_1(ces_21_6_io_outs_1),
    .io_outs_2(ces_21_6_io_outs_2),
    .io_outs_3(ces_21_6_io_outs_3)
  );
  Element ces_21_7 ( // @[MockArray.scala 36:52]
    .clock(ces_21_7_clock),
    .io_ins_0(ces_21_7_io_ins_0),
    .io_ins_1(ces_21_7_io_ins_1),
    .io_ins_2(ces_21_7_io_ins_2),
    .io_ins_3(ces_21_7_io_ins_3),
    .io_outs_0(ces_21_7_io_outs_0),
    .io_outs_1(ces_21_7_io_outs_1),
    .io_outs_2(ces_21_7_io_outs_2),
    .io_outs_3(ces_21_7_io_outs_3)
  );
  Element ces_21_8 ( // @[MockArray.scala 36:52]
    .clock(ces_21_8_clock),
    .io_ins_0(ces_21_8_io_ins_0),
    .io_ins_1(ces_21_8_io_ins_1),
    .io_ins_2(ces_21_8_io_ins_2),
    .io_ins_3(ces_21_8_io_ins_3),
    .io_outs_0(ces_21_8_io_outs_0),
    .io_outs_1(ces_21_8_io_outs_1),
    .io_outs_2(ces_21_8_io_outs_2),
    .io_outs_3(ces_21_8_io_outs_3)
  );
  Element ces_21_9 ( // @[MockArray.scala 36:52]
    .clock(ces_21_9_clock),
    .io_ins_0(ces_21_9_io_ins_0),
    .io_ins_1(ces_21_9_io_ins_1),
    .io_ins_2(ces_21_9_io_ins_2),
    .io_ins_3(ces_21_9_io_ins_3),
    .io_outs_0(ces_21_9_io_outs_0),
    .io_outs_1(ces_21_9_io_outs_1),
    .io_outs_2(ces_21_9_io_outs_2),
    .io_outs_3(ces_21_9_io_outs_3)
  );
  Element ces_21_10 ( // @[MockArray.scala 36:52]
    .clock(ces_21_10_clock),
    .io_ins_0(ces_21_10_io_ins_0),
    .io_ins_1(ces_21_10_io_ins_1),
    .io_ins_2(ces_21_10_io_ins_2),
    .io_ins_3(ces_21_10_io_ins_3),
    .io_outs_0(ces_21_10_io_outs_0),
    .io_outs_1(ces_21_10_io_outs_1),
    .io_outs_2(ces_21_10_io_outs_2),
    .io_outs_3(ces_21_10_io_outs_3)
  );
  Element ces_21_11 ( // @[MockArray.scala 36:52]
    .clock(ces_21_11_clock),
    .io_ins_0(ces_21_11_io_ins_0),
    .io_ins_1(ces_21_11_io_ins_1),
    .io_ins_2(ces_21_11_io_ins_2),
    .io_ins_3(ces_21_11_io_ins_3),
    .io_outs_0(ces_21_11_io_outs_0),
    .io_outs_1(ces_21_11_io_outs_1),
    .io_outs_2(ces_21_11_io_outs_2),
    .io_outs_3(ces_21_11_io_outs_3)
  );
  Element ces_21_12 ( // @[MockArray.scala 36:52]
    .clock(ces_21_12_clock),
    .io_ins_0(ces_21_12_io_ins_0),
    .io_ins_1(ces_21_12_io_ins_1),
    .io_ins_2(ces_21_12_io_ins_2),
    .io_ins_3(ces_21_12_io_ins_3),
    .io_outs_0(ces_21_12_io_outs_0),
    .io_outs_1(ces_21_12_io_outs_1),
    .io_outs_2(ces_21_12_io_outs_2),
    .io_outs_3(ces_21_12_io_outs_3)
  );
  Element ces_21_13 ( // @[MockArray.scala 36:52]
    .clock(ces_21_13_clock),
    .io_ins_0(ces_21_13_io_ins_0),
    .io_ins_1(ces_21_13_io_ins_1),
    .io_ins_2(ces_21_13_io_ins_2),
    .io_ins_3(ces_21_13_io_ins_3),
    .io_outs_0(ces_21_13_io_outs_0),
    .io_outs_1(ces_21_13_io_outs_1),
    .io_outs_2(ces_21_13_io_outs_2),
    .io_outs_3(ces_21_13_io_outs_3)
  );
  Element ces_21_14 ( // @[MockArray.scala 36:52]
    .clock(ces_21_14_clock),
    .io_ins_0(ces_21_14_io_ins_0),
    .io_ins_1(ces_21_14_io_ins_1),
    .io_ins_2(ces_21_14_io_ins_2),
    .io_ins_3(ces_21_14_io_ins_3),
    .io_outs_0(ces_21_14_io_outs_0),
    .io_outs_1(ces_21_14_io_outs_1),
    .io_outs_2(ces_21_14_io_outs_2),
    .io_outs_3(ces_21_14_io_outs_3)
  );
  Element ces_21_15 ( // @[MockArray.scala 36:52]
    .clock(ces_21_15_clock),
    .io_ins_0(ces_21_15_io_ins_0),
    .io_ins_1(ces_21_15_io_ins_1),
    .io_ins_2(ces_21_15_io_ins_2),
    .io_ins_3(ces_21_15_io_ins_3),
    .io_outs_0(ces_21_15_io_outs_0),
    .io_outs_1(ces_21_15_io_outs_1),
    .io_outs_2(ces_21_15_io_outs_2),
    .io_outs_3(ces_21_15_io_outs_3)
  );
  Element ces_21_16 ( // @[MockArray.scala 36:52]
    .clock(ces_21_16_clock),
    .io_ins_0(ces_21_16_io_ins_0),
    .io_ins_1(ces_21_16_io_ins_1),
    .io_ins_2(ces_21_16_io_ins_2),
    .io_ins_3(ces_21_16_io_ins_3),
    .io_outs_0(ces_21_16_io_outs_0),
    .io_outs_1(ces_21_16_io_outs_1),
    .io_outs_2(ces_21_16_io_outs_2),
    .io_outs_3(ces_21_16_io_outs_3)
  );
  Element ces_21_17 ( // @[MockArray.scala 36:52]
    .clock(ces_21_17_clock),
    .io_ins_0(ces_21_17_io_ins_0),
    .io_ins_1(ces_21_17_io_ins_1),
    .io_ins_2(ces_21_17_io_ins_2),
    .io_ins_3(ces_21_17_io_ins_3),
    .io_outs_0(ces_21_17_io_outs_0),
    .io_outs_1(ces_21_17_io_outs_1),
    .io_outs_2(ces_21_17_io_outs_2),
    .io_outs_3(ces_21_17_io_outs_3)
  );
  Element ces_21_18 ( // @[MockArray.scala 36:52]
    .clock(ces_21_18_clock),
    .io_ins_0(ces_21_18_io_ins_0),
    .io_ins_1(ces_21_18_io_ins_1),
    .io_ins_2(ces_21_18_io_ins_2),
    .io_ins_3(ces_21_18_io_ins_3),
    .io_outs_0(ces_21_18_io_outs_0),
    .io_outs_1(ces_21_18_io_outs_1),
    .io_outs_2(ces_21_18_io_outs_2),
    .io_outs_3(ces_21_18_io_outs_3)
  );
  Element ces_21_19 ( // @[MockArray.scala 36:52]
    .clock(ces_21_19_clock),
    .io_ins_0(ces_21_19_io_ins_0),
    .io_ins_1(ces_21_19_io_ins_1),
    .io_ins_2(ces_21_19_io_ins_2),
    .io_ins_3(ces_21_19_io_ins_3),
    .io_outs_0(ces_21_19_io_outs_0),
    .io_outs_1(ces_21_19_io_outs_1),
    .io_outs_2(ces_21_19_io_outs_2),
    .io_outs_3(ces_21_19_io_outs_3)
  );
  Element ces_21_20 ( // @[MockArray.scala 36:52]
    .clock(ces_21_20_clock),
    .io_ins_0(ces_21_20_io_ins_0),
    .io_ins_1(ces_21_20_io_ins_1),
    .io_ins_2(ces_21_20_io_ins_2),
    .io_ins_3(ces_21_20_io_ins_3),
    .io_outs_0(ces_21_20_io_outs_0),
    .io_outs_1(ces_21_20_io_outs_1),
    .io_outs_2(ces_21_20_io_outs_2),
    .io_outs_3(ces_21_20_io_outs_3)
  );
  Element ces_21_21 ( // @[MockArray.scala 36:52]
    .clock(ces_21_21_clock),
    .io_ins_0(ces_21_21_io_ins_0),
    .io_ins_1(ces_21_21_io_ins_1),
    .io_ins_2(ces_21_21_io_ins_2),
    .io_ins_3(ces_21_21_io_ins_3),
    .io_outs_0(ces_21_21_io_outs_0),
    .io_outs_1(ces_21_21_io_outs_1),
    .io_outs_2(ces_21_21_io_outs_2),
    .io_outs_3(ces_21_21_io_outs_3)
  );
  Element ces_21_22 ( // @[MockArray.scala 36:52]
    .clock(ces_21_22_clock),
    .io_ins_0(ces_21_22_io_ins_0),
    .io_ins_1(ces_21_22_io_ins_1),
    .io_ins_2(ces_21_22_io_ins_2),
    .io_ins_3(ces_21_22_io_ins_3),
    .io_outs_0(ces_21_22_io_outs_0),
    .io_outs_1(ces_21_22_io_outs_1),
    .io_outs_2(ces_21_22_io_outs_2),
    .io_outs_3(ces_21_22_io_outs_3)
  );
  Element ces_21_23 ( // @[MockArray.scala 36:52]
    .clock(ces_21_23_clock),
    .io_ins_0(ces_21_23_io_ins_0),
    .io_ins_1(ces_21_23_io_ins_1),
    .io_ins_2(ces_21_23_io_ins_2),
    .io_ins_3(ces_21_23_io_ins_3),
    .io_outs_0(ces_21_23_io_outs_0),
    .io_outs_1(ces_21_23_io_outs_1),
    .io_outs_2(ces_21_23_io_outs_2),
    .io_outs_3(ces_21_23_io_outs_3)
  );
  Element ces_21_24 ( // @[MockArray.scala 36:52]
    .clock(ces_21_24_clock),
    .io_ins_0(ces_21_24_io_ins_0),
    .io_ins_1(ces_21_24_io_ins_1),
    .io_ins_2(ces_21_24_io_ins_2),
    .io_ins_3(ces_21_24_io_ins_3),
    .io_outs_0(ces_21_24_io_outs_0),
    .io_outs_1(ces_21_24_io_outs_1),
    .io_outs_2(ces_21_24_io_outs_2),
    .io_outs_3(ces_21_24_io_outs_3)
  );
  Element ces_21_25 ( // @[MockArray.scala 36:52]
    .clock(ces_21_25_clock),
    .io_ins_0(ces_21_25_io_ins_0),
    .io_ins_1(ces_21_25_io_ins_1),
    .io_ins_2(ces_21_25_io_ins_2),
    .io_ins_3(ces_21_25_io_ins_3),
    .io_outs_0(ces_21_25_io_outs_0),
    .io_outs_1(ces_21_25_io_outs_1),
    .io_outs_2(ces_21_25_io_outs_2),
    .io_outs_3(ces_21_25_io_outs_3)
  );
  Element ces_21_26 ( // @[MockArray.scala 36:52]
    .clock(ces_21_26_clock),
    .io_ins_0(ces_21_26_io_ins_0),
    .io_ins_1(ces_21_26_io_ins_1),
    .io_ins_2(ces_21_26_io_ins_2),
    .io_ins_3(ces_21_26_io_ins_3),
    .io_outs_0(ces_21_26_io_outs_0),
    .io_outs_1(ces_21_26_io_outs_1),
    .io_outs_2(ces_21_26_io_outs_2),
    .io_outs_3(ces_21_26_io_outs_3)
  );
  Element ces_21_27 ( // @[MockArray.scala 36:52]
    .clock(ces_21_27_clock),
    .io_ins_0(ces_21_27_io_ins_0),
    .io_ins_1(ces_21_27_io_ins_1),
    .io_ins_2(ces_21_27_io_ins_2),
    .io_ins_3(ces_21_27_io_ins_3),
    .io_outs_0(ces_21_27_io_outs_0),
    .io_outs_1(ces_21_27_io_outs_1),
    .io_outs_2(ces_21_27_io_outs_2),
    .io_outs_3(ces_21_27_io_outs_3)
  );
  Element ces_21_28 ( // @[MockArray.scala 36:52]
    .clock(ces_21_28_clock),
    .io_ins_0(ces_21_28_io_ins_0),
    .io_ins_1(ces_21_28_io_ins_1),
    .io_ins_2(ces_21_28_io_ins_2),
    .io_ins_3(ces_21_28_io_ins_3),
    .io_outs_0(ces_21_28_io_outs_0),
    .io_outs_1(ces_21_28_io_outs_1),
    .io_outs_2(ces_21_28_io_outs_2),
    .io_outs_3(ces_21_28_io_outs_3)
  );
  Element ces_21_29 ( // @[MockArray.scala 36:52]
    .clock(ces_21_29_clock),
    .io_ins_0(ces_21_29_io_ins_0),
    .io_ins_1(ces_21_29_io_ins_1),
    .io_ins_2(ces_21_29_io_ins_2),
    .io_ins_3(ces_21_29_io_ins_3),
    .io_outs_0(ces_21_29_io_outs_0),
    .io_outs_1(ces_21_29_io_outs_1),
    .io_outs_2(ces_21_29_io_outs_2),
    .io_outs_3(ces_21_29_io_outs_3)
  );
  Element ces_21_30 ( // @[MockArray.scala 36:52]
    .clock(ces_21_30_clock),
    .io_ins_0(ces_21_30_io_ins_0),
    .io_ins_1(ces_21_30_io_ins_1),
    .io_ins_2(ces_21_30_io_ins_2),
    .io_ins_3(ces_21_30_io_ins_3),
    .io_outs_0(ces_21_30_io_outs_0),
    .io_outs_1(ces_21_30_io_outs_1),
    .io_outs_2(ces_21_30_io_outs_2),
    .io_outs_3(ces_21_30_io_outs_3)
  );
  Element ces_21_31 ( // @[MockArray.scala 36:52]
    .clock(ces_21_31_clock),
    .io_ins_0(ces_21_31_io_ins_0),
    .io_ins_1(ces_21_31_io_ins_1),
    .io_ins_2(ces_21_31_io_ins_2),
    .io_ins_3(ces_21_31_io_ins_3),
    .io_outs_0(ces_21_31_io_outs_0),
    .io_outs_1(ces_21_31_io_outs_1),
    .io_outs_2(ces_21_31_io_outs_2),
    .io_outs_3(ces_21_31_io_outs_3)
  );
  Element ces_22_0 ( // @[MockArray.scala 36:52]
    .clock(ces_22_0_clock),
    .io_ins_0(ces_22_0_io_ins_0),
    .io_ins_1(ces_22_0_io_ins_1),
    .io_ins_2(ces_22_0_io_ins_2),
    .io_ins_3(ces_22_0_io_ins_3),
    .io_outs_0(ces_22_0_io_outs_0),
    .io_outs_1(ces_22_0_io_outs_1),
    .io_outs_2(ces_22_0_io_outs_2),
    .io_outs_3(ces_22_0_io_outs_3)
  );
  Element ces_22_1 ( // @[MockArray.scala 36:52]
    .clock(ces_22_1_clock),
    .io_ins_0(ces_22_1_io_ins_0),
    .io_ins_1(ces_22_1_io_ins_1),
    .io_ins_2(ces_22_1_io_ins_2),
    .io_ins_3(ces_22_1_io_ins_3),
    .io_outs_0(ces_22_1_io_outs_0),
    .io_outs_1(ces_22_1_io_outs_1),
    .io_outs_2(ces_22_1_io_outs_2),
    .io_outs_3(ces_22_1_io_outs_3)
  );
  Element ces_22_2 ( // @[MockArray.scala 36:52]
    .clock(ces_22_2_clock),
    .io_ins_0(ces_22_2_io_ins_0),
    .io_ins_1(ces_22_2_io_ins_1),
    .io_ins_2(ces_22_2_io_ins_2),
    .io_ins_3(ces_22_2_io_ins_3),
    .io_outs_0(ces_22_2_io_outs_0),
    .io_outs_1(ces_22_2_io_outs_1),
    .io_outs_2(ces_22_2_io_outs_2),
    .io_outs_3(ces_22_2_io_outs_3)
  );
  Element ces_22_3 ( // @[MockArray.scala 36:52]
    .clock(ces_22_3_clock),
    .io_ins_0(ces_22_3_io_ins_0),
    .io_ins_1(ces_22_3_io_ins_1),
    .io_ins_2(ces_22_3_io_ins_2),
    .io_ins_3(ces_22_3_io_ins_3),
    .io_outs_0(ces_22_3_io_outs_0),
    .io_outs_1(ces_22_3_io_outs_1),
    .io_outs_2(ces_22_3_io_outs_2),
    .io_outs_3(ces_22_3_io_outs_3)
  );
  Element ces_22_4 ( // @[MockArray.scala 36:52]
    .clock(ces_22_4_clock),
    .io_ins_0(ces_22_4_io_ins_0),
    .io_ins_1(ces_22_4_io_ins_1),
    .io_ins_2(ces_22_4_io_ins_2),
    .io_ins_3(ces_22_4_io_ins_3),
    .io_outs_0(ces_22_4_io_outs_0),
    .io_outs_1(ces_22_4_io_outs_1),
    .io_outs_2(ces_22_4_io_outs_2),
    .io_outs_3(ces_22_4_io_outs_3)
  );
  Element ces_22_5 ( // @[MockArray.scala 36:52]
    .clock(ces_22_5_clock),
    .io_ins_0(ces_22_5_io_ins_0),
    .io_ins_1(ces_22_5_io_ins_1),
    .io_ins_2(ces_22_5_io_ins_2),
    .io_ins_3(ces_22_5_io_ins_3),
    .io_outs_0(ces_22_5_io_outs_0),
    .io_outs_1(ces_22_5_io_outs_1),
    .io_outs_2(ces_22_5_io_outs_2),
    .io_outs_3(ces_22_5_io_outs_3)
  );
  Element ces_22_6 ( // @[MockArray.scala 36:52]
    .clock(ces_22_6_clock),
    .io_ins_0(ces_22_6_io_ins_0),
    .io_ins_1(ces_22_6_io_ins_1),
    .io_ins_2(ces_22_6_io_ins_2),
    .io_ins_3(ces_22_6_io_ins_3),
    .io_outs_0(ces_22_6_io_outs_0),
    .io_outs_1(ces_22_6_io_outs_1),
    .io_outs_2(ces_22_6_io_outs_2),
    .io_outs_3(ces_22_6_io_outs_3)
  );
  Element ces_22_7 ( // @[MockArray.scala 36:52]
    .clock(ces_22_7_clock),
    .io_ins_0(ces_22_7_io_ins_0),
    .io_ins_1(ces_22_7_io_ins_1),
    .io_ins_2(ces_22_7_io_ins_2),
    .io_ins_3(ces_22_7_io_ins_3),
    .io_outs_0(ces_22_7_io_outs_0),
    .io_outs_1(ces_22_7_io_outs_1),
    .io_outs_2(ces_22_7_io_outs_2),
    .io_outs_3(ces_22_7_io_outs_3)
  );
  Element ces_22_8 ( // @[MockArray.scala 36:52]
    .clock(ces_22_8_clock),
    .io_ins_0(ces_22_8_io_ins_0),
    .io_ins_1(ces_22_8_io_ins_1),
    .io_ins_2(ces_22_8_io_ins_2),
    .io_ins_3(ces_22_8_io_ins_3),
    .io_outs_0(ces_22_8_io_outs_0),
    .io_outs_1(ces_22_8_io_outs_1),
    .io_outs_2(ces_22_8_io_outs_2),
    .io_outs_3(ces_22_8_io_outs_3)
  );
  Element ces_22_9 ( // @[MockArray.scala 36:52]
    .clock(ces_22_9_clock),
    .io_ins_0(ces_22_9_io_ins_0),
    .io_ins_1(ces_22_9_io_ins_1),
    .io_ins_2(ces_22_9_io_ins_2),
    .io_ins_3(ces_22_9_io_ins_3),
    .io_outs_0(ces_22_9_io_outs_0),
    .io_outs_1(ces_22_9_io_outs_1),
    .io_outs_2(ces_22_9_io_outs_2),
    .io_outs_3(ces_22_9_io_outs_3)
  );
  Element ces_22_10 ( // @[MockArray.scala 36:52]
    .clock(ces_22_10_clock),
    .io_ins_0(ces_22_10_io_ins_0),
    .io_ins_1(ces_22_10_io_ins_1),
    .io_ins_2(ces_22_10_io_ins_2),
    .io_ins_3(ces_22_10_io_ins_3),
    .io_outs_0(ces_22_10_io_outs_0),
    .io_outs_1(ces_22_10_io_outs_1),
    .io_outs_2(ces_22_10_io_outs_2),
    .io_outs_3(ces_22_10_io_outs_3)
  );
  Element ces_22_11 ( // @[MockArray.scala 36:52]
    .clock(ces_22_11_clock),
    .io_ins_0(ces_22_11_io_ins_0),
    .io_ins_1(ces_22_11_io_ins_1),
    .io_ins_2(ces_22_11_io_ins_2),
    .io_ins_3(ces_22_11_io_ins_3),
    .io_outs_0(ces_22_11_io_outs_0),
    .io_outs_1(ces_22_11_io_outs_1),
    .io_outs_2(ces_22_11_io_outs_2),
    .io_outs_3(ces_22_11_io_outs_3)
  );
  Element ces_22_12 ( // @[MockArray.scala 36:52]
    .clock(ces_22_12_clock),
    .io_ins_0(ces_22_12_io_ins_0),
    .io_ins_1(ces_22_12_io_ins_1),
    .io_ins_2(ces_22_12_io_ins_2),
    .io_ins_3(ces_22_12_io_ins_3),
    .io_outs_0(ces_22_12_io_outs_0),
    .io_outs_1(ces_22_12_io_outs_1),
    .io_outs_2(ces_22_12_io_outs_2),
    .io_outs_3(ces_22_12_io_outs_3)
  );
  Element ces_22_13 ( // @[MockArray.scala 36:52]
    .clock(ces_22_13_clock),
    .io_ins_0(ces_22_13_io_ins_0),
    .io_ins_1(ces_22_13_io_ins_1),
    .io_ins_2(ces_22_13_io_ins_2),
    .io_ins_3(ces_22_13_io_ins_3),
    .io_outs_0(ces_22_13_io_outs_0),
    .io_outs_1(ces_22_13_io_outs_1),
    .io_outs_2(ces_22_13_io_outs_2),
    .io_outs_3(ces_22_13_io_outs_3)
  );
  Element ces_22_14 ( // @[MockArray.scala 36:52]
    .clock(ces_22_14_clock),
    .io_ins_0(ces_22_14_io_ins_0),
    .io_ins_1(ces_22_14_io_ins_1),
    .io_ins_2(ces_22_14_io_ins_2),
    .io_ins_3(ces_22_14_io_ins_3),
    .io_outs_0(ces_22_14_io_outs_0),
    .io_outs_1(ces_22_14_io_outs_1),
    .io_outs_2(ces_22_14_io_outs_2),
    .io_outs_3(ces_22_14_io_outs_3)
  );
  Element ces_22_15 ( // @[MockArray.scala 36:52]
    .clock(ces_22_15_clock),
    .io_ins_0(ces_22_15_io_ins_0),
    .io_ins_1(ces_22_15_io_ins_1),
    .io_ins_2(ces_22_15_io_ins_2),
    .io_ins_3(ces_22_15_io_ins_3),
    .io_outs_0(ces_22_15_io_outs_0),
    .io_outs_1(ces_22_15_io_outs_1),
    .io_outs_2(ces_22_15_io_outs_2),
    .io_outs_3(ces_22_15_io_outs_3)
  );
  Element ces_22_16 ( // @[MockArray.scala 36:52]
    .clock(ces_22_16_clock),
    .io_ins_0(ces_22_16_io_ins_0),
    .io_ins_1(ces_22_16_io_ins_1),
    .io_ins_2(ces_22_16_io_ins_2),
    .io_ins_3(ces_22_16_io_ins_3),
    .io_outs_0(ces_22_16_io_outs_0),
    .io_outs_1(ces_22_16_io_outs_1),
    .io_outs_2(ces_22_16_io_outs_2),
    .io_outs_3(ces_22_16_io_outs_3)
  );
  Element ces_22_17 ( // @[MockArray.scala 36:52]
    .clock(ces_22_17_clock),
    .io_ins_0(ces_22_17_io_ins_0),
    .io_ins_1(ces_22_17_io_ins_1),
    .io_ins_2(ces_22_17_io_ins_2),
    .io_ins_3(ces_22_17_io_ins_3),
    .io_outs_0(ces_22_17_io_outs_0),
    .io_outs_1(ces_22_17_io_outs_1),
    .io_outs_2(ces_22_17_io_outs_2),
    .io_outs_3(ces_22_17_io_outs_3)
  );
  Element ces_22_18 ( // @[MockArray.scala 36:52]
    .clock(ces_22_18_clock),
    .io_ins_0(ces_22_18_io_ins_0),
    .io_ins_1(ces_22_18_io_ins_1),
    .io_ins_2(ces_22_18_io_ins_2),
    .io_ins_3(ces_22_18_io_ins_3),
    .io_outs_0(ces_22_18_io_outs_0),
    .io_outs_1(ces_22_18_io_outs_1),
    .io_outs_2(ces_22_18_io_outs_2),
    .io_outs_3(ces_22_18_io_outs_3)
  );
  Element ces_22_19 ( // @[MockArray.scala 36:52]
    .clock(ces_22_19_clock),
    .io_ins_0(ces_22_19_io_ins_0),
    .io_ins_1(ces_22_19_io_ins_1),
    .io_ins_2(ces_22_19_io_ins_2),
    .io_ins_3(ces_22_19_io_ins_3),
    .io_outs_0(ces_22_19_io_outs_0),
    .io_outs_1(ces_22_19_io_outs_1),
    .io_outs_2(ces_22_19_io_outs_2),
    .io_outs_3(ces_22_19_io_outs_3)
  );
  Element ces_22_20 ( // @[MockArray.scala 36:52]
    .clock(ces_22_20_clock),
    .io_ins_0(ces_22_20_io_ins_0),
    .io_ins_1(ces_22_20_io_ins_1),
    .io_ins_2(ces_22_20_io_ins_2),
    .io_ins_3(ces_22_20_io_ins_3),
    .io_outs_0(ces_22_20_io_outs_0),
    .io_outs_1(ces_22_20_io_outs_1),
    .io_outs_2(ces_22_20_io_outs_2),
    .io_outs_3(ces_22_20_io_outs_3)
  );
  Element ces_22_21 ( // @[MockArray.scala 36:52]
    .clock(ces_22_21_clock),
    .io_ins_0(ces_22_21_io_ins_0),
    .io_ins_1(ces_22_21_io_ins_1),
    .io_ins_2(ces_22_21_io_ins_2),
    .io_ins_3(ces_22_21_io_ins_3),
    .io_outs_0(ces_22_21_io_outs_0),
    .io_outs_1(ces_22_21_io_outs_1),
    .io_outs_2(ces_22_21_io_outs_2),
    .io_outs_3(ces_22_21_io_outs_3)
  );
  Element ces_22_22 ( // @[MockArray.scala 36:52]
    .clock(ces_22_22_clock),
    .io_ins_0(ces_22_22_io_ins_0),
    .io_ins_1(ces_22_22_io_ins_1),
    .io_ins_2(ces_22_22_io_ins_2),
    .io_ins_3(ces_22_22_io_ins_3),
    .io_outs_0(ces_22_22_io_outs_0),
    .io_outs_1(ces_22_22_io_outs_1),
    .io_outs_2(ces_22_22_io_outs_2),
    .io_outs_3(ces_22_22_io_outs_3)
  );
  Element ces_22_23 ( // @[MockArray.scala 36:52]
    .clock(ces_22_23_clock),
    .io_ins_0(ces_22_23_io_ins_0),
    .io_ins_1(ces_22_23_io_ins_1),
    .io_ins_2(ces_22_23_io_ins_2),
    .io_ins_3(ces_22_23_io_ins_3),
    .io_outs_0(ces_22_23_io_outs_0),
    .io_outs_1(ces_22_23_io_outs_1),
    .io_outs_2(ces_22_23_io_outs_2),
    .io_outs_3(ces_22_23_io_outs_3)
  );
  Element ces_22_24 ( // @[MockArray.scala 36:52]
    .clock(ces_22_24_clock),
    .io_ins_0(ces_22_24_io_ins_0),
    .io_ins_1(ces_22_24_io_ins_1),
    .io_ins_2(ces_22_24_io_ins_2),
    .io_ins_3(ces_22_24_io_ins_3),
    .io_outs_0(ces_22_24_io_outs_0),
    .io_outs_1(ces_22_24_io_outs_1),
    .io_outs_2(ces_22_24_io_outs_2),
    .io_outs_3(ces_22_24_io_outs_3)
  );
  Element ces_22_25 ( // @[MockArray.scala 36:52]
    .clock(ces_22_25_clock),
    .io_ins_0(ces_22_25_io_ins_0),
    .io_ins_1(ces_22_25_io_ins_1),
    .io_ins_2(ces_22_25_io_ins_2),
    .io_ins_3(ces_22_25_io_ins_3),
    .io_outs_0(ces_22_25_io_outs_0),
    .io_outs_1(ces_22_25_io_outs_1),
    .io_outs_2(ces_22_25_io_outs_2),
    .io_outs_3(ces_22_25_io_outs_3)
  );
  Element ces_22_26 ( // @[MockArray.scala 36:52]
    .clock(ces_22_26_clock),
    .io_ins_0(ces_22_26_io_ins_0),
    .io_ins_1(ces_22_26_io_ins_1),
    .io_ins_2(ces_22_26_io_ins_2),
    .io_ins_3(ces_22_26_io_ins_3),
    .io_outs_0(ces_22_26_io_outs_0),
    .io_outs_1(ces_22_26_io_outs_1),
    .io_outs_2(ces_22_26_io_outs_2),
    .io_outs_3(ces_22_26_io_outs_3)
  );
  Element ces_22_27 ( // @[MockArray.scala 36:52]
    .clock(ces_22_27_clock),
    .io_ins_0(ces_22_27_io_ins_0),
    .io_ins_1(ces_22_27_io_ins_1),
    .io_ins_2(ces_22_27_io_ins_2),
    .io_ins_3(ces_22_27_io_ins_3),
    .io_outs_0(ces_22_27_io_outs_0),
    .io_outs_1(ces_22_27_io_outs_1),
    .io_outs_2(ces_22_27_io_outs_2),
    .io_outs_3(ces_22_27_io_outs_3)
  );
  Element ces_22_28 ( // @[MockArray.scala 36:52]
    .clock(ces_22_28_clock),
    .io_ins_0(ces_22_28_io_ins_0),
    .io_ins_1(ces_22_28_io_ins_1),
    .io_ins_2(ces_22_28_io_ins_2),
    .io_ins_3(ces_22_28_io_ins_3),
    .io_outs_0(ces_22_28_io_outs_0),
    .io_outs_1(ces_22_28_io_outs_1),
    .io_outs_2(ces_22_28_io_outs_2),
    .io_outs_3(ces_22_28_io_outs_3)
  );
  Element ces_22_29 ( // @[MockArray.scala 36:52]
    .clock(ces_22_29_clock),
    .io_ins_0(ces_22_29_io_ins_0),
    .io_ins_1(ces_22_29_io_ins_1),
    .io_ins_2(ces_22_29_io_ins_2),
    .io_ins_3(ces_22_29_io_ins_3),
    .io_outs_0(ces_22_29_io_outs_0),
    .io_outs_1(ces_22_29_io_outs_1),
    .io_outs_2(ces_22_29_io_outs_2),
    .io_outs_3(ces_22_29_io_outs_3)
  );
  Element ces_22_30 ( // @[MockArray.scala 36:52]
    .clock(ces_22_30_clock),
    .io_ins_0(ces_22_30_io_ins_0),
    .io_ins_1(ces_22_30_io_ins_1),
    .io_ins_2(ces_22_30_io_ins_2),
    .io_ins_3(ces_22_30_io_ins_3),
    .io_outs_0(ces_22_30_io_outs_0),
    .io_outs_1(ces_22_30_io_outs_1),
    .io_outs_2(ces_22_30_io_outs_2),
    .io_outs_3(ces_22_30_io_outs_3)
  );
  Element ces_22_31 ( // @[MockArray.scala 36:52]
    .clock(ces_22_31_clock),
    .io_ins_0(ces_22_31_io_ins_0),
    .io_ins_1(ces_22_31_io_ins_1),
    .io_ins_2(ces_22_31_io_ins_2),
    .io_ins_3(ces_22_31_io_ins_3),
    .io_outs_0(ces_22_31_io_outs_0),
    .io_outs_1(ces_22_31_io_outs_1),
    .io_outs_2(ces_22_31_io_outs_2),
    .io_outs_3(ces_22_31_io_outs_3)
  );
  Element ces_23_0 ( // @[MockArray.scala 36:52]
    .clock(ces_23_0_clock),
    .io_ins_0(ces_23_0_io_ins_0),
    .io_ins_1(ces_23_0_io_ins_1),
    .io_ins_2(ces_23_0_io_ins_2),
    .io_ins_3(ces_23_0_io_ins_3),
    .io_outs_0(ces_23_0_io_outs_0),
    .io_outs_1(ces_23_0_io_outs_1),
    .io_outs_2(ces_23_0_io_outs_2),
    .io_outs_3(ces_23_0_io_outs_3)
  );
  Element ces_23_1 ( // @[MockArray.scala 36:52]
    .clock(ces_23_1_clock),
    .io_ins_0(ces_23_1_io_ins_0),
    .io_ins_1(ces_23_1_io_ins_1),
    .io_ins_2(ces_23_1_io_ins_2),
    .io_ins_3(ces_23_1_io_ins_3),
    .io_outs_0(ces_23_1_io_outs_0),
    .io_outs_1(ces_23_1_io_outs_1),
    .io_outs_2(ces_23_1_io_outs_2),
    .io_outs_3(ces_23_1_io_outs_3)
  );
  Element ces_23_2 ( // @[MockArray.scala 36:52]
    .clock(ces_23_2_clock),
    .io_ins_0(ces_23_2_io_ins_0),
    .io_ins_1(ces_23_2_io_ins_1),
    .io_ins_2(ces_23_2_io_ins_2),
    .io_ins_3(ces_23_2_io_ins_3),
    .io_outs_0(ces_23_2_io_outs_0),
    .io_outs_1(ces_23_2_io_outs_1),
    .io_outs_2(ces_23_2_io_outs_2),
    .io_outs_3(ces_23_2_io_outs_3)
  );
  Element ces_23_3 ( // @[MockArray.scala 36:52]
    .clock(ces_23_3_clock),
    .io_ins_0(ces_23_3_io_ins_0),
    .io_ins_1(ces_23_3_io_ins_1),
    .io_ins_2(ces_23_3_io_ins_2),
    .io_ins_3(ces_23_3_io_ins_3),
    .io_outs_0(ces_23_3_io_outs_0),
    .io_outs_1(ces_23_3_io_outs_1),
    .io_outs_2(ces_23_3_io_outs_2),
    .io_outs_3(ces_23_3_io_outs_3)
  );
  Element ces_23_4 ( // @[MockArray.scala 36:52]
    .clock(ces_23_4_clock),
    .io_ins_0(ces_23_4_io_ins_0),
    .io_ins_1(ces_23_4_io_ins_1),
    .io_ins_2(ces_23_4_io_ins_2),
    .io_ins_3(ces_23_4_io_ins_3),
    .io_outs_0(ces_23_4_io_outs_0),
    .io_outs_1(ces_23_4_io_outs_1),
    .io_outs_2(ces_23_4_io_outs_2),
    .io_outs_3(ces_23_4_io_outs_3)
  );
  Element ces_23_5 ( // @[MockArray.scala 36:52]
    .clock(ces_23_5_clock),
    .io_ins_0(ces_23_5_io_ins_0),
    .io_ins_1(ces_23_5_io_ins_1),
    .io_ins_2(ces_23_5_io_ins_2),
    .io_ins_3(ces_23_5_io_ins_3),
    .io_outs_0(ces_23_5_io_outs_0),
    .io_outs_1(ces_23_5_io_outs_1),
    .io_outs_2(ces_23_5_io_outs_2),
    .io_outs_3(ces_23_5_io_outs_3)
  );
  Element ces_23_6 ( // @[MockArray.scala 36:52]
    .clock(ces_23_6_clock),
    .io_ins_0(ces_23_6_io_ins_0),
    .io_ins_1(ces_23_6_io_ins_1),
    .io_ins_2(ces_23_6_io_ins_2),
    .io_ins_3(ces_23_6_io_ins_3),
    .io_outs_0(ces_23_6_io_outs_0),
    .io_outs_1(ces_23_6_io_outs_1),
    .io_outs_2(ces_23_6_io_outs_2),
    .io_outs_3(ces_23_6_io_outs_3)
  );
  Element ces_23_7 ( // @[MockArray.scala 36:52]
    .clock(ces_23_7_clock),
    .io_ins_0(ces_23_7_io_ins_0),
    .io_ins_1(ces_23_7_io_ins_1),
    .io_ins_2(ces_23_7_io_ins_2),
    .io_ins_3(ces_23_7_io_ins_3),
    .io_outs_0(ces_23_7_io_outs_0),
    .io_outs_1(ces_23_7_io_outs_1),
    .io_outs_2(ces_23_7_io_outs_2),
    .io_outs_3(ces_23_7_io_outs_3)
  );
  Element ces_23_8 ( // @[MockArray.scala 36:52]
    .clock(ces_23_8_clock),
    .io_ins_0(ces_23_8_io_ins_0),
    .io_ins_1(ces_23_8_io_ins_1),
    .io_ins_2(ces_23_8_io_ins_2),
    .io_ins_3(ces_23_8_io_ins_3),
    .io_outs_0(ces_23_8_io_outs_0),
    .io_outs_1(ces_23_8_io_outs_1),
    .io_outs_2(ces_23_8_io_outs_2),
    .io_outs_3(ces_23_8_io_outs_3)
  );
  Element ces_23_9 ( // @[MockArray.scala 36:52]
    .clock(ces_23_9_clock),
    .io_ins_0(ces_23_9_io_ins_0),
    .io_ins_1(ces_23_9_io_ins_1),
    .io_ins_2(ces_23_9_io_ins_2),
    .io_ins_3(ces_23_9_io_ins_3),
    .io_outs_0(ces_23_9_io_outs_0),
    .io_outs_1(ces_23_9_io_outs_1),
    .io_outs_2(ces_23_9_io_outs_2),
    .io_outs_3(ces_23_9_io_outs_3)
  );
  Element ces_23_10 ( // @[MockArray.scala 36:52]
    .clock(ces_23_10_clock),
    .io_ins_0(ces_23_10_io_ins_0),
    .io_ins_1(ces_23_10_io_ins_1),
    .io_ins_2(ces_23_10_io_ins_2),
    .io_ins_3(ces_23_10_io_ins_3),
    .io_outs_0(ces_23_10_io_outs_0),
    .io_outs_1(ces_23_10_io_outs_1),
    .io_outs_2(ces_23_10_io_outs_2),
    .io_outs_3(ces_23_10_io_outs_3)
  );
  Element ces_23_11 ( // @[MockArray.scala 36:52]
    .clock(ces_23_11_clock),
    .io_ins_0(ces_23_11_io_ins_0),
    .io_ins_1(ces_23_11_io_ins_1),
    .io_ins_2(ces_23_11_io_ins_2),
    .io_ins_3(ces_23_11_io_ins_3),
    .io_outs_0(ces_23_11_io_outs_0),
    .io_outs_1(ces_23_11_io_outs_1),
    .io_outs_2(ces_23_11_io_outs_2),
    .io_outs_3(ces_23_11_io_outs_3)
  );
  Element ces_23_12 ( // @[MockArray.scala 36:52]
    .clock(ces_23_12_clock),
    .io_ins_0(ces_23_12_io_ins_0),
    .io_ins_1(ces_23_12_io_ins_1),
    .io_ins_2(ces_23_12_io_ins_2),
    .io_ins_3(ces_23_12_io_ins_3),
    .io_outs_0(ces_23_12_io_outs_0),
    .io_outs_1(ces_23_12_io_outs_1),
    .io_outs_2(ces_23_12_io_outs_2),
    .io_outs_3(ces_23_12_io_outs_3)
  );
  Element ces_23_13 ( // @[MockArray.scala 36:52]
    .clock(ces_23_13_clock),
    .io_ins_0(ces_23_13_io_ins_0),
    .io_ins_1(ces_23_13_io_ins_1),
    .io_ins_2(ces_23_13_io_ins_2),
    .io_ins_3(ces_23_13_io_ins_3),
    .io_outs_0(ces_23_13_io_outs_0),
    .io_outs_1(ces_23_13_io_outs_1),
    .io_outs_2(ces_23_13_io_outs_2),
    .io_outs_3(ces_23_13_io_outs_3)
  );
  Element ces_23_14 ( // @[MockArray.scala 36:52]
    .clock(ces_23_14_clock),
    .io_ins_0(ces_23_14_io_ins_0),
    .io_ins_1(ces_23_14_io_ins_1),
    .io_ins_2(ces_23_14_io_ins_2),
    .io_ins_3(ces_23_14_io_ins_3),
    .io_outs_0(ces_23_14_io_outs_0),
    .io_outs_1(ces_23_14_io_outs_1),
    .io_outs_2(ces_23_14_io_outs_2),
    .io_outs_3(ces_23_14_io_outs_3)
  );
  Element ces_23_15 ( // @[MockArray.scala 36:52]
    .clock(ces_23_15_clock),
    .io_ins_0(ces_23_15_io_ins_0),
    .io_ins_1(ces_23_15_io_ins_1),
    .io_ins_2(ces_23_15_io_ins_2),
    .io_ins_3(ces_23_15_io_ins_3),
    .io_outs_0(ces_23_15_io_outs_0),
    .io_outs_1(ces_23_15_io_outs_1),
    .io_outs_2(ces_23_15_io_outs_2),
    .io_outs_3(ces_23_15_io_outs_3)
  );
  Element ces_23_16 ( // @[MockArray.scala 36:52]
    .clock(ces_23_16_clock),
    .io_ins_0(ces_23_16_io_ins_0),
    .io_ins_1(ces_23_16_io_ins_1),
    .io_ins_2(ces_23_16_io_ins_2),
    .io_ins_3(ces_23_16_io_ins_3),
    .io_outs_0(ces_23_16_io_outs_0),
    .io_outs_1(ces_23_16_io_outs_1),
    .io_outs_2(ces_23_16_io_outs_2),
    .io_outs_3(ces_23_16_io_outs_3)
  );
  Element ces_23_17 ( // @[MockArray.scala 36:52]
    .clock(ces_23_17_clock),
    .io_ins_0(ces_23_17_io_ins_0),
    .io_ins_1(ces_23_17_io_ins_1),
    .io_ins_2(ces_23_17_io_ins_2),
    .io_ins_3(ces_23_17_io_ins_3),
    .io_outs_0(ces_23_17_io_outs_0),
    .io_outs_1(ces_23_17_io_outs_1),
    .io_outs_2(ces_23_17_io_outs_2),
    .io_outs_3(ces_23_17_io_outs_3)
  );
  Element ces_23_18 ( // @[MockArray.scala 36:52]
    .clock(ces_23_18_clock),
    .io_ins_0(ces_23_18_io_ins_0),
    .io_ins_1(ces_23_18_io_ins_1),
    .io_ins_2(ces_23_18_io_ins_2),
    .io_ins_3(ces_23_18_io_ins_3),
    .io_outs_0(ces_23_18_io_outs_0),
    .io_outs_1(ces_23_18_io_outs_1),
    .io_outs_2(ces_23_18_io_outs_2),
    .io_outs_3(ces_23_18_io_outs_3)
  );
  Element ces_23_19 ( // @[MockArray.scala 36:52]
    .clock(ces_23_19_clock),
    .io_ins_0(ces_23_19_io_ins_0),
    .io_ins_1(ces_23_19_io_ins_1),
    .io_ins_2(ces_23_19_io_ins_2),
    .io_ins_3(ces_23_19_io_ins_3),
    .io_outs_0(ces_23_19_io_outs_0),
    .io_outs_1(ces_23_19_io_outs_1),
    .io_outs_2(ces_23_19_io_outs_2),
    .io_outs_3(ces_23_19_io_outs_3)
  );
  Element ces_23_20 ( // @[MockArray.scala 36:52]
    .clock(ces_23_20_clock),
    .io_ins_0(ces_23_20_io_ins_0),
    .io_ins_1(ces_23_20_io_ins_1),
    .io_ins_2(ces_23_20_io_ins_2),
    .io_ins_3(ces_23_20_io_ins_3),
    .io_outs_0(ces_23_20_io_outs_0),
    .io_outs_1(ces_23_20_io_outs_1),
    .io_outs_2(ces_23_20_io_outs_2),
    .io_outs_3(ces_23_20_io_outs_3)
  );
  Element ces_23_21 ( // @[MockArray.scala 36:52]
    .clock(ces_23_21_clock),
    .io_ins_0(ces_23_21_io_ins_0),
    .io_ins_1(ces_23_21_io_ins_1),
    .io_ins_2(ces_23_21_io_ins_2),
    .io_ins_3(ces_23_21_io_ins_3),
    .io_outs_0(ces_23_21_io_outs_0),
    .io_outs_1(ces_23_21_io_outs_1),
    .io_outs_2(ces_23_21_io_outs_2),
    .io_outs_3(ces_23_21_io_outs_3)
  );
  Element ces_23_22 ( // @[MockArray.scala 36:52]
    .clock(ces_23_22_clock),
    .io_ins_0(ces_23_22_io_ins_0),
    .io_ins_1(ces_23_22_io_ins_1),
    .io_ins_2(ces_23_22_io_ins_2),
    .io_ins_3(ces_23_22_io_ins_3),
    .io_outs_0(ces_23_22_io_outs_0),
    .io_outs_1(ces_23_22_io_outs_1),
    .io_outs_2(ces_23_22_io_outs_2),
    .io_outs_3(ces_23_22_io_outs_3)
  );
  Element ces_23_23 ( // @[MockArray.scala 36:52]
    .clock(ces_23_23_clock),
    .io_ins_0(ces_23_23_io_ins_0),
    .io_ins_1(ces_23_23_io_ins_1),
    .io_ins_2(ces_23_23_io_ins_2),
    .io_ins_3(ces_23_23_io_ins_3),
    .io_outs_0(ces_23_23_io_outs_0),
    .io_outs_1(ces_23_23_io_outs_1),
    .io_outs_2(ces_23_23_io_outs_2),
    .io_outs_3(ces_23_23_io_outs_3)
  );
  Element ces_23_24 ( // @[MockArray.scala 36:52]
    .clock(ces_23_24_clock),
    .io_ins_0(ces_23_24_io_ins_0),
    .io_ins_1(ces_23_24_io_ins_1),
    .io_ins_2(ces_23_24_io_ins_2),
    .io_ins_3(ces_23_24_io_ins_3),
    .io_outs_0(ces_23_24_io_outs_0),
    .io_outs_1(ces_23_24_io_outs_1),
    .io_outs_2(ces_23_24_io_outs_2),
    .io_outs_3(ces_23_24_io_outs_3)
  );
  Element ces_23_25 ( // @[MockArray.scala 36:52]
    .clock(ces_23_25_clock),
    .io_ins_0(ces_23_25_io_ins_0),
    .io_ins_1(ces_23_25_io_ins_1),
    .io_ins_2(ces_23_25_io_ins_2),
    .io_ins_3(ces_23_25_io_ins_3),
    .io_outs_0(ces_23_25_io_outs_0),
    .io_outs_1(ces_23_25_io_outs_1),
    .io_outs_2(ces_23_25_io_outs_2),
    .io_outs_3(ces_23_25_io_outs_3)
  );
  Element ces_23_26 ( // @[MockArray.scala 36:52]
    .clock(ces_23_26_clock),
    .io_ins_0(ces_23_26_io_ins_0),
    .io_ins_1(ces_23_26_io_ins_1),
    .io_ins_2(ces_23_26_io_ins_2),
    .io_ins_3(ces_23_26_io_ins_3),
    .io_outs_0(ces_23_26_io_outs_0),
    .io_outs_1(ces_23_26_io_outs_1),
    .io_outs_2(ces_23_26_io_outs_2),
    .io_outs_3(ces_23_26_io_outs_3)
  );
  Element ces_23_27 ( // @[MockArray.scala 36:52]
    .clock(ces_23_27_clock),
    .io_ins_0(ces_23_27_io_ins_0),
    .io_ins_1(ces_23_27_io_ins_1),
    .io_ins_2(ces_23_27_io_ins_2),
    .io_ins_3(ces_23_27_io_ins_3),
    .io_outs_0(ces_23_27_io_outs_0),
    .io_outs_1(ces_23_27_io_outs_1),
    .io_outs_2(ces_23_27_io_outs_2),
    .io_outs_3(ces_23_27_io_outs_3)
  );
  Element ces_23_28 ( // @[MockArray.scala 36:52]
    .clock(ces_23_28_clock),
    .io_ins_0(ces_23_28_io_ins_0),
    .io_ins_1(ces_23_28_io_ins_1),
    .io_ins_2(ces_23_28_io_ins_2),
    .io_ins_3(ces_23_28_io_ins_3),
    .io_outs_0(ces_23_28_io_outs_0),
    .io_outs_1(ces_23_28_io_outs_1),
    .io_outs_2(ces_23_28_io_outs_2),
    .io_outs_3(ces_23_28_io_outs_3)
  );
  Element ces_23_29 ( // @[MockArray.scala 36:52]
    .clock(ces_23_29_clock),
    .io_ins_0(ces_23_29_io_ins_0),
    .io_ins_1(ces_23_29_io_ins_1),
    .io_ins_2(ces_23_29_io_ins_2),
    .io_ins_3(ces_23_29_io_ins_3),
    .io_outs_0(ces_23_29_io_outs_0),
    .io_outs_1(ces_23_29_io_outs_1),
    .io_outs_2(ces_23_29_io_outs_2),
    .io_outs_3(ces_23_29_io_outs_3)
  );
  Element ces_23_30 ( // @[MockArray.scala 36:52]
    .clock(ces_23_30_clock),
    .io_ins_0(ces_23_30_io_ins_0),
    .io_ins_1(ces_23_30_io_ins_1),
    .io_ins_2(ces_23_30_io_ins_2),
    .io_ins_3(ces_23_30_io_ins_3),
    .io_outs_0(ces_23_30_io_outs_0),
    .io_outs_1(ces_23_30_io_outs_1),
    .io_outs_2(ces_23_30_io_outs_2),
    .io_outs_3(ces_23_30_io_outs_3)
  );
  Element ces_23_31 ( // @[MockArray.scala 36:52]
    .clock(ces_23_31_clock),
    .io_ins_0(ces_23_31_io_ins_0),
    .io_ins_1(ces_23_31_io_ins_1),
    .io_ins_2(ces_23_31_io_ins_2),
    .io_ins_3(ces_23_31_io_ins_3),
    .io_outs_0(ces_23_31_io_outs_0),
    .io_outs_1(ces_23_31_io_outs_1),
    .io_outs_2(ces_23_31_io_outs_2),
    .io_outs_3(ces_23_31_io_outs_3)
  );
  Element ces_24_0 ( // @[MockArray.scala 36:52]
    .clock(ces_24_0_clock),
    .io_ins_0(ces_24_0_io_ins_0),
    .io_ins_1(ces_24_0_io_ins_1),
    .io_ins_2(ces_24_0_io_ins_2),
    .io_ins_3(ces_24_0_io_ins_3),
    .io_outs_0(ces_24_0_io_outs_0),
    .io_outs_1(ces_24_0_io_outs_1),
    .io_outs_2(ces_24_0_io_outs_2),
    .io_outs_3(ces_24_0_io_outs_3)
  );
  Element ces_24_1 ( // @[MockArray.scala 36:52]
    .clock(ces_24_1_clock),
    .io_ins_0(ces_24_1_io_ins_0),
    .io_ins_1(ces_24_1_io_ins_1),
    .io_ins_2(ces_24_1_io_ins_2),
    .io_ins_3(ces_24_1_io_ins_3),
    .io_outs_0(ces_24_1_io_outs_0),
    .io_outs_1(ces_24_1_io_outs_1),
    .io_outs_2(ces_24_1_io_outs_2),
    .io_outs_3(ces_24_1_io_outs_3)
  );
  Element ces_24_2 ( // @[MockArray.scala 36:52]
    .clock(ces_24_2_clock),
    .io_ins_0(ces_24_2_io_ins_0),
    .io_ins_1(ces_24_2_io_ins_1),
    .io_ins_2(ces_24_2_io_ins_2),
    .io_ins_3(ces_24_2_io_ins_3),
    .io_outs_0(ces_24_2_io_outs_0),
    .io_outs_1(ces_24_2_io_outs_1),
    .io_outs_2(ces_24_2_io_outs_2),
    .io_outs_3(ces_24_2_io_outs_3)
  );
  Element ces_24_3 ( // @[MockArray.scala 36:52]
    .clock(ces_24_3_clock),
    .io_ins_0(ces_24_3_io_ins_0),
    .io_ins_1(ces_24_3_io_ins_1),
    .io_ins_2(ces_24_3_io_ins_2),
    .io_ins_3(ces_24_3_io_ins_3),
    .io_outs_0(ces_24_3_io_outs_0),
    .io_outs_1(ces_24_3_io_outs_1),
    .io_outs_2(ces_24_3_io_outs_2),
    .io_outs_3(ces_24_3_io_outs_3)
  );
  Element ces_24_4 ( // @[MockArray.scala 36:52]
    .clock(ces_24_4_clock),
    .io_ins_0(ces_24_4_io_ins_0),
    .io_ins_1(ces_24_4_io_ins_1),
    .io_ins_2(ces_24_4_io_ins_2),
    .io_ins_3(ces_24_4_io_ins_3),
    .io_outs_0(ces_24_4_io_outs_0),
    .io_outs_1(ces_24_4_io_outs_1),
    .io_outs_2(ces_24_4_io_outs_2),
    .io_outs_3(ces_24_4_io_outs_3)
  );
  Element ces_24_5 ( // @[MockArray.scala 36:52]
    .clock(ces_24_5_clock),
    .io_ins_0(ces_24_5_io_ins_0),
    .io_ins_1(ces_24_5_io_ins_1),
    .io_ins_2(ces_24_5_io_ins_2),
    .io_ins_3(ces_24_5_io_ins_3),
    .io_outs_0(ces_24_5_io_outs_0),
    .io_outs_1(ces_24_5_io_outs_1),
    .io_outs_2(ces_24_5_io_outs_2),
    .io_outs_3(ces_24_5_io_outs_3)
  );
  Element ces_24_6 ( // @[MockArray.scala 36:52]
    .clock(ces_24_6_clock),
    .io_ins_0(ces_24_6_io_ins_0),
    .io_ins_1(ces_24_6_io_ins_1),
    .io_ins_2(ces_24_6_io_ins_2),
    .io_ins_3(ces_24_6_io_ins_3),
    .io_outs_0(ces_24_6_io_outs_0),
    .io_outs_1(ces_24_6_io_outs_1),
    .io_outs_2(ces_24_6_io_outs_2),
    .io_outs_3(ces_24_6_io_outs_3)
  );
  Element ces_24_7 ( // @[MockArray.scala 36:52]
    .clock(ces_24_7_clock),
    .io_ins_0(ces_24_7_io_ins_0),
    .io_ins_1(ces_24_7_io_ins_1),
    .io_ins_2(ces_24_7_io_ins_2),
    .io_ins_3(ces_24_7_io_ins_3),
    .io_outs_0(ces_24_7_io_outs_0),
    .io_outs_1(ces_24_7_io_outs_1),
    .io_outs_2(ces_24_7_io_outs_2),
    .io_outs_3(ces_24_7_io_outs_3)
  );
  Element ces_24_8 ( // @[MockArray.scala 36:52]
    .clock(ces_24_8_clock),
    .io_ins_0(ces_24_8_io_ins_0),
    .io_ins_1(ces_24_8_io_ins_1),
    .io_ins_2(ces_24_8_io_ins_2),
    .io_ins_3(ces_24_8_io_ins_3),
    .io_outs_0(ces_24_8_io_outs_0),
    .io_outs_1(ces_24_8_io_outs_1),
    .io_outs_2(ces_24_8_io_outs_2),
    .io_outs_3(ces_24_8_io_outs_3)
  );
  Element ces_24_9 ( // @[MockArray.scala 36:52]
    .clock(ces_24_9_clock),
    .io_ins_0(ces_24_9_io_ins_0),
    .io_ins_1(ces_24_9_io_ins_1),
    .io_ins_2(ces_24_9_io_ins_2),
    .io_ins_3(ces_24_9_io_ins_3),
    .io_outs_0(ces_24_9_io_outs_0),
    .io_outs_1(ces_24_9_io_outs_1),
    .io_outs_2(ces_24_9_io_outs_2),
    .io_outs_3(ces_24_9_io_outs_3)
  );
  Element ces_24_10 ( // @[MockArray.scala 36:52]
    .clock(ces_24_10_clock),
    .io_ins_0(ces_24_10_io_ins_0),
    .io_ins_1(ces_24_10_io_ins_1),
    .io_ins_2(ces_24_10_io_ins_2),
    .io_ins_3(ces_24_10_io_ins_3),
    .io_outs_0(ces_24_10_io_outs_0),
    .io_outs_1(ces_24_10_io_outs_1),
    .io_outs_2(ces_24_10_io_outs_2),
    .io_outs_3(ces_24_10_io_outs_3)
  );
  Element ces_24_11 ( // @[MockArray.scala 36:52]
    .clock(ces_24_11_clock),
    .io_ins_0(ces_24_11_io_ins_0),
    .io_ins_1(ces_24_11_io_ins_1),
    .io_ins_2(ces_24_11_io_ins_2),
    .io_ins_3(ces_24_11_io_ins_3),
    .io_outs_0(ces_24_11_io_outs_0),
    .io_outs_1(ces_24_11_io_outs_1),
    .io_outs_2(ces_24_11_io_outs_2),
    .io_outs_3(ces_24_11_io_outs_3)
  );
  Element ces_24_12 ( // @[MockArray.scala 36:52]
    .clock(ces_24_12_clock),
    .io_ins_0(ces_24_12_io_ins_0),
    .io_ins_1(ces_24_12_io_ins_1),
    .io_ins_2(ces_24_12_io_ins_2),
    .io_ins_3(ces_24_12_io_ins_3),
    .io_outs_0(ces_24_12_io_outs_0),
    .io_outs_1(ces_24_12_io_outs_1),
    .io_outs_2(ces_24_12_io_outs_2),
    .io_outs_3(ces_24_12_io_outs_3)
  );
  Element ces_24_13 ( // @[MockArray.scala 36:52]
    .clock(ces_24_13_clock),
    .io_ins_0(ces_24_13_io_ins_0),
    .io_ins_1(ces_24_13_io_ins_1),
    .io_ins_2(ces_24_13_io_ins_2),
    .io_ins_3(ces_24_13_io_ins_3),
    .io_outs_0(ces_24_13_io_outs_0),
    .io_outs_1(ces_24_13_io_outs_1),
    .io_outs_2(ces_24_13_io_outs_2),
    .io_outs_3(ces_24_13_io_outs_3)
  );
  Element ces_24_14 ( // @[MockArray.scala 36:52]
    .clock(ces_24_14_clock),
    .io_ins_0(ces_24_14_io_ins_0),
    .io_ins_1(ces_24_14_io_ins_1),
    .io_ins_2(ces_24_14_io_ins_2),
    .io_ins_3(ces_24_14_io_ins_3),
    .io_outs_0(ces_24_14_io_outs_0),
    .io_outs_1(ces_24_14_io_outs_1),
    .io_outs_2(ces_24_14_io_outs_2),
    .io_outs_3(ces_24_14_io_outs_3)
  );
  Element ces_24_15 ( // @[MockArray.scala 36:52]
    .clock(ces_24_15_clock),
    .io_ins_0(ces_24_15_io_ins_0),
    .io_ins_1(ces_24_15_io_ins_1),
    .io_ins_2(ces_24_15_io_ins_2),
    .io_ins_3(ces_24_15_io_ins_3),
    .io_outs_0(ces_24_15_io_outs_0),
    .io_outs_1(ces_24_15_io_outs_1),
    .io_outs_2(ces_24_15_io_outs_2),
    .io_outs_3(ces_24_15_io_outs_3)
  );
  Element ces_24_16 ( // @[MockArray.scala 36:52]
    .clock(ces_24_16_clock),
    .io_ins_0(ces_24_16_io_ins_0),
    .io_ins_1(ces_24_16_io_ins_1),
    .io_ins_2(ces_24_16_io_ins_2),
    .io_ins_3(ces_24_16_io_ins_3),
    .io_outs_0(ces_24_16_io_outs_0),
    .io_outs_1(ces_24_16_io_outs_1),
    .io_outs_2(ces_24_16_io_outs_2),
    .io_outs_3(ces_24_16_io_outs_3)
  );
  Element ces_24_17 ( // @[MockArray.scala 36:52]
    .clock(ces_24_17_clock),
    .io_ins_0(ces_24_17_io_ins_0),
    .io_ins_1(ces_24_17_io_ins_1),
    .io_ins_2(ces_24_17_io_ins_2),
    .io_ins_3(ces_24_17_io_ins_3),
    .io_outs_0(ces_24_17_io_outs_0),
    .io_outs_1(ces_24_17_io_outs_1),
    .io_outs_2(ces_24_17_io_outs_2),
    .io_outs_3(ces_24_17_io_outs_3)
  );
  Element ces_24_18 ( // @[MockArray.scala 36:52]
    .clock(ces_24_18_clock),
    .io_ins_0(ces_24_18_io_ins_0),
    .io_ins_1(ces_24_18_io_ins_1),
    .io_ins_2(ces_24_18_io_ins_2),
    .io_ins_3(ces_24_18_io_ins_3),
    .io_outs_0(ces_24_18_io_outs_0),
    .io_outs_1(ces_24_18_io_outs_1),
    .io_outs_2(ces_24_18_io_outs_2),
    .io_outs_3(ces_24_18_io_outs_3)
  );
  Element ces_24_19 ( // @[MockArray.scala 36:52]
    .clock(ces_24_19_clock),
    .io_ins_0(ces_24_19_io_ins_0),
    .io_ins_1(ces_24_19_io_ins_1),
    .io_ins_2(ces_24_19_io_ins_2),
    .io_ins_3(ces_24_19_io_ins_3),
    .io_outs_0(ces_24_19_io_outs_0),
    .io_outs_1(ces_24_19_io_outs_1),
    .io_outs_2(ces_24_19_io_outs_2),
    .io_outs_3(ces_24_19_io_outs_3)
  );
  Element ces_24_20 ( // @[MockArray.scala 36:52]
    .clock(ces_24_20_clock),
    .io_ins_0(ces_24_20_io_ins_0),
    .io_ins_1(ces_24_20_io_ins_1),
    .io_ins_2(ces_24_20_io_ins_2),
    .io_ins_3(ces_24_20_io_ins_3),
    .io_outs_0(ces_24_20_io_outs_0),
    .io_outs_1(ces_24_20_io_outs_1),
    .io_outs_2(ces_24_20_io_outs_2),
    .io_outs_3(ces_24_20_io_outs_3)
  );
  Element ces_24_21 ( // @[MockArray.scala 36:52]
    .clock(ces_24_21_clock),
    .io_ins_0(ces_24_21_io_ins_0),
    .io_ins_1(ces_24_21_io_ins_1),
    .io_ins_2(ces_24_21_io_ins_2),
    .io_ins_3(ces_24_21_io_ins_3),
    .io_outs_0(ces_24_21_io_outs_0),
    .io_outs_1(ces_24_21_io_outs_1),
    .io_outs_2(ces_24_21_io_outs_2),
    .io_outs_3(ces_24_21_io_outs_3)
  );
  Element ces_24_22 ( // @[MockArray.scala 36:52]
    .clock(ces_24_22_clock),
    .io_ins_0(ces_24_22_io_ins_0),
    .io_ins_1(ces_24_22_io_ins_1),
    .io_ins_2(ces_24_22_io_ins_2),
    .io_ins_3(ces_24_22_io_ins_3),
    .io_outs_0(ces_24_22_io_outs_0),
    .io_outs_1(ces_24_22_io_outs_1),
    .io_outs_2(ces_24_22_io_outs_2),
    .io_outs_3(ces_24_22_io_outs_3)
  );
  Element ces_24_23 ( // @[MockArray.scala 36:52]
    .clock(ces_24_23_clock),
    .io_ins_0(ces_24_23_io_ins_0),
    .io_ins_1(ces_24_23_io_ins_1),
    .io_ins_2(ces_24_23_io_ins_2),
    .io_ins_3(ces_24_23_io_ins_3),
    .io_outs_0(ces_24_23_io_outs_0),
    .io_outs_1(ces_24_23_io_outs_1),
    .io_outs_2(ces_24_23_io_outs_2),
    .io_outs_3(ces_24_23_io_outs_3)
  );
  Element ces_24_24 ( // @[MockArray.scala 36:52]
    .clock(ces_24_24_clock),
    .io_ins_0(ces_24_24_io_ins_0),
    .io_ins_1(ces_24_24_io_ins_1),
    .io_ins_2(ces_24_24_io_ins_2),
    .io_ins_3(ces_24_24_io_ins_3),
    .io_outs_0(ces_24_24_io_outs_0),
    .io_outs_1(ces_24_24_io_outs_1),
    .io_outs_2(ces_24_24_io_outs_2),
    .io_outs_3(ces_24_24_io_outs_3)
  );
  Element ces_24_25 ( // @[MockArray.scala 36:52]
    .clock(ces_24_25_clock),
    .io_ins_0(ces_24_25_io_ins_0),
    .io_ins_1(ces_24_25_io_ins_1),
    .io_ins_2(ces_24_25_io_ins_2),
    .io_ins_3(ces_24_25_io_ins_3),
    .io_outs_0(ces_24_25_io_outs_0),
    .io_outs_1(ces_24_25_io_outs_1),
    .io_outs_2(ces_24_25_io_outs_2),
    .io_outs_3(ces_24_25_io_outs_3)
  );
  Element ces_24_26 ( // @[MockArray.scala 36:52]
    .clock(ces_24_26_clock),
    .io_ins_0(ces_24_26_io_ins_0),
    .io_ins_1(ces_24_26_io_ins_1),
    .io_ins_2(ces_24_26_io_ins_2),
    .io_ins_3(ces_24_26_io_ins_3),
    .io_outs_0(ces_24_26_io_outs_0),
    .io_outs_1(ces_24_26_io_outs_1),
    .io_outs_2(ces_24_26_io_outs_2),
    .io_outs_3(ces_24_26_io_outs_3)
  );
  Element ces_24_27 ( // @[MockArray.scala 36:52]
    .clock(ces_24_27_clock),
    .io_ins_0(ces_24_27_io_ins_0),
    .io_ins_1(ces_24_27_io_ins_1),
    .io_ins_2(ces_24_27_io_ins_2),
    .io_ins_3(ces_24_27_io_ins_3),
    .io_outs_0(ces_24_27_io_outs_0),
    .io_outs_1(ces_24_27_io_outs_1),
    .io_outs_2(ces_24_27_io_outs_2),
    .io_outs_3(ces_24_27_io_outs_3)
  );
  Element ces_24_28 ( // @[MockArray.scala 36:52]
    .clock(ces_24_28_clock),
    .io_ins_0(ces_24_28_io_ins_0),
    .io_ins_1(ces_24_28_io_ins_1),
    .io_ins_2(ces_24_28_io_ins_2),
    .io_ins_3(ces_24_28_io_ins_3),
    .io_outs_0(ces_24_28_io_outs_0),
    .io_outs_1(ces_24_28_io_outs_1),
    .io_outs_2(ces_24_28_io_outs_2),
    .io_outs_3(ces_24_28_io_outs_3)
  );
  Element ces_24_29 ( // @[MockArray.scala 36:52]
    .clock(ces_24_29_clock),
    .io_ins_0(ces_24_29_io_ins_0),
    .io_ins_1(ces_24_29_io_ins_1),
    .io_ins_2(ces_24_29_io_ins_2),
    .io_ins_3(ces_24_29_io_ins_3),
    .io_outs_0(ces_24_29_io_outs_0),
    .io_outs_1(ces_24_29_io_outs_1),
    .io_outs_2(ces_24_29_io_outs_2),
    .io_outs_3(ces_24_29_io_outs_3)
  );
  Element ces_24_30 ( // @[MockArray.scala 36:52]
    .clock(ces_24_30_clock),
    .io_ins_0(ces_24_30_io_ins_0),
    .io_ins_1(ces_24_30_io_ins_1),
    .io_ins_2(ces_24_30_io_ins_2),
    .io_ins_3(ces_24_30_io_ins_3),
    .io_outs_0(ces_24_30_io_outs_0),
    .io_outs_1(ces_24_30_io_outs_1),
    .io_outs_2(ces_24_30_io_outs_2),
    .io_outs_3(ces_24_30_io_outs_3)
  );
  Element ces_24_31 ( // @[MockArray.scala 36:52]
    .clock(ces_24_31_clock),
    .io_ins_0(ces_24_31_io_ins_0),
    .io_ins_1(ces_24_31_io_ins_1),
    .io_ins_2(ces_24_31_io_ins_2),
    .io_ins_3(ces_24_31_io_ins_3),
    .io_outs_0(ces_24_31_io_outs_0),
    .io_outs_1(ces_24_31_io_outs_1),
    .io_outs_2(ces_24_31_io_outs_2),
    .io_outs_3(ces_24_31_io_outs_3)
  );
  Element ces_25_0 ( // @[MockArray.scala 36:52]
    .clock(ces_25_0_clock),
    .io_ins_0(ces_25_0_io_ins_0),
    .io_ins_1(ces_25_0_io_ins_1),
    .io_ins_2(ces_25_0_io_ins_2),
    .io_ins_3(ces_25_0_io_ins_3),
    .io_outs_0(ces_25_0_io_outs_0),
    .io_outs_1(ces_25_0_io_outs_1),
    .io_outs_2(ces_25_0_io_outs_2),
    .io_outs_3(ces_25_0_io_outs_3)
  );
  Element ces_25_1 ( // @[MockArray.scala 36:52]
    .clock(ces_25_1_clock),
    .io_ins_0(ces_25_1_io_ins_0),
    .io_ins_1(ces_25_1_io_ins_1),
    .io_ins_2(ces_25_1_io_ins_2),
    .io_ins_3(ces_25_1_io_ins_3),
    .io_outs_0(ces_25_1_io_outs_0),
    .io_outs_1(ces_25_1_io_outs_1),
    .io_outs_2(ces_25_1_io_outs_2),
    .io_outs_3(ces_25_1_io_outs_3)
  );
  Element ces_25_2 ( // @[MockArray.scala 36:52]
    .clock(ces_25_2_clock),
    .io_ins_0(ces_25_2_io_ins_0),
    .io_ins_1(ces_25_2_io_ins_1),
    .io_ins_2(ces_25_2_io_ins_2),
    .io_ins_3(ces_25_2_io_ins_3),
    .io_outs_0(ces_25_2_io_outs_0),
    .io_outs_1(ces_25_2_io_outs_1),
    .io_outs_2(ces_25_2_io_outs_2),
    .io_outs_3(ces_25_2_io_outs_3)
  );
  Element ces_25_3 ( // @[MockArray.scala 36:52]
    .clock(ces_25_3_clock),
    .io_ins_0(ces_25_3_io_ins_0),
    .io_ins_1(ces_25_3_io_ins_1),
    .io_ins_2(ces_25_3_io_ins_2),
    .io_ins_3(ces_25_3_io_ins_3),
    .io_outs_0(ces_25_3_io_outs_0),
    .io_outs_1(ces_25_3_io_outs_1),
    .io_outs_2(ces_25_3_io_outs_2),
    .io_outs_3(ces_25_3_io_outs_3)
  );
  Element ces_25_4 ( // @[MockArray.scala 36:52]
    .clock(ces_25_4_clock),
    .io_ins_0(ces_25_4_io_ins_0),
    .io_ins_1(ces_25_4_io_ins_1),
    .io_ins_2(ces_25_4_io_ins_2),
    .io_ins_3(ces_25_4_io_ins_3),
    .io_outs_0(ces_25_4_io_outs_0),
    .io_outs_1(ces_25_4_io_outs_1),
    .io_outs_2(ces_25_4_io_outs_2),
    .io_outs_3(ces_25_4_io_outs_3)
  );
  Element ces_25_5 ( // @[MockArray.scala 36:52]
    .clock(ces_25_5_clock),
    .io_ins_0(ces_25_5_io_ins_0),
    .io_ins_1(ces_25_5_io_ins_1),
    .io_ins_2(ces_25_5_io_ins_2),
    .io_ins_3(ces_25_5_io_ins_3),
    .io_outs_0(ces_25_5_io_outs_0),
    .io_outs_1(ces_25_5_io_outs_1),
    .io_outs_2(ces_25_5_io_outs_2),
    .io_outs_3(ces_25_5_io_outs_3)
  );
  Element ces_25_6 ( // @[MockArray.scala 36:52]
    .clock(ces_25_6_clock),
    .io_ins_0(ces_25_6_io_ins_0),
    .io_ins_1(ces_25_6_io_ins_1),
    .io_ins_2(ces_25_6_io_ins_2),
    .io_ins_3(ces_25_6_io_ins_3),
    .io_outs_0(ces_25_6_io_outs_0),
    .io_outs_1(ces_25_6_io_outs_1),
    .io_outs_2(ces_25_6_io_outs_2),
    .io_outs_3(ces_25_6_io_outs_3)
  );
  Element ces_25_7 ( // @[MockArray.scala 36:52]
    .clock(ces_25_7_clock),
    .io_ins_0(ces_25_7_io_ins_0),
    .io_ins_1(ces_25_7_io_ins_1),
    .io_ins_2(ces_25_7_io_ins_2),
    .io_ins_3(ces_25_7_io_ins_3),
    .io_outs_0(ces_25_7_io_outs_0),
    .io_outs_1(ces_25_7_io_outs_1),
    .io_outs_2(ces_25_7_io_outs_2),
    .io_outs_3(ces_25_7_io_outs_3)
  );
  Element ces_25_8 ( // @[MockArray.scala 36:52]
    .clock(ces_25_8_clock),
    .io_ins_0(ces_25_8_io_ins_0),
    .io_ins_1(ces_25_8_io_ins_1),
    .io_ins_2(ces_25_8_io_ins_2),
    .io_ins_3(ces_25_8_io_ins_3),
    .io_outs_0(ces_25_8_io_outs_0),
    .io_outs_1(ces_25_8_io_outs_1),
    .io_outs_2(ces_25_8_io_outs_2),
    .io_outs_3(ces_25_8_io_outs_3)
  );
  Element ces_25_9 ( // @[MockArray.scala 36:52]
    .clock(ces_25_9_clock),
    .io_ins_0(ces_25_9_io_ins_0),
    .io_ins_1(ces_25_9_io_ins_1),
    .io_ins_2(ces_25_9_io_ins_2),
    .io_ins_3(ces_25_9_io_ins_3),
    .io_outs_0(ces_25_9_io_outs_0),
    .io_outs_1(ces_25_9_io_outs_1),
    .io_outs_2(ces_25_9_io_outs_2),
    .io_outs_3(ces_25_9_io_outs_3)
  );
  Element ces_25_10 ( // @[MockArray.scala 36:52]
    .clock(ces_25_10_clock),
    .io_ins_0(ces_25_10_io_ins_0),
    .io_ins_1(ces_25_10_io_ins_1),
    .io_ins_2(ces_25_10_io_ins_2),
    .io_ins_3(ces_25_10_io_ins_3),
    .io_outs_0(ces_25_10_io_outs_0),
    .io_outs_1(ces_25_10_io_outs_1),
    .io_outs_2(ces_25_10_io_outs_2),
    .io_outs_3(ces_25_10_io_outs_3)
  );
  Element ces_25_11 ( // @[MockArray.scala 36:52]
    .clock(ces_25_11_clock),
    .io_ins_0(ces_25_11_io_ins_0),
    .io_ins_1(ces_25_11_io_ins_1),
    .io_ins_2(ces_25_11_io_ins_2),
    .io_ins_3(ces_25_11_io_ins_3),
    .io_outs_0(ces_25_11_io_outs_0),
    .io_outs_1(ces_25_11_io_outs_1),
    .io_outs_2(ces_25_11_io_outs_2),
    .io_outs_3(ces_25_11_io_outs_3)
  );
  Element ces_25_12 ( // @[MockArray.scala 36:52]
    .clock(ces_25_12_clock),
    .io_ins_0(ces_25_12_io_ins_0),
    .io_ins_1(ces_25_12_io_ins_1),
    .io_ins_2(ces_25_12_io_ins_2),
    .io_ins_3(ces_25_12_io_ins_3),
    .io_outs_0(ces_25_12_io_outs_0),
    .io_outs_1(ces_25_12_io_outs_1),
    .io_outs_2(ces_25_12_io_outs_2),
    .io_outs_3(ces_25_12_io_outs_3)
  );
  Element ces_25_13 ( // @[MockArray.scala 36:52]
    .clock(ces_25_13_clock),
    .io_ins_0(ces_25_13_io_ins_0),
    .io_ins_1(ces_25_13_io_ins_1),
    .io_ins_2(ces_25_13_io_ins_2),
    .io_ins_3(ces_25_13_io_ins_3),
    .io_outs_0(ces_25_13_io_outs_0),
    .io_outs_1(ces_25_13_io_outs_1),
    .io_outs_2(ces_25_13_io_outs_2),
    .io_outs_3(ces_25_13_io_outs_3)
  );
  Element ces_25_14 ( // @[MockArray.scala 36:52]
    .clock(ces_25_14_clock),
    .io_ins_0(ces_25_14_io_ins_0),
    .io_ins_1(ces_25_14_io_ins_1),
    .io_ins_2(ces_25_14_io_ins_2),
    .io_ins_3(ces_25_14_io_ins_3),
    .io_outs_0(ces_25_14_io_outs_0),
    .io_outs_1(ces_25_14_io_outs_1),
    .io_outs_2(ces_25_14_io_outs_2),
    .io_outs_3(ces_25_14_io_outs_3)
  );
  Element ces_25_15 ( // @[MockArray.scala 36:52]
    .clock(ces_25_15_clock),
    .io_ins_0(ces_25_15_io_ins_0),
    .io_ins_1(ces_25_15_io_ins_1),
    .io_ins_2(ces_25_15_io_ins_2),
    .io_ins_3(ces_25_15_io_ins_3),
    .io_outs_0(ces_25_15_io_outs_0),
    .io_outs_1(ces_25_15_io_outs_1),
    .io_outs_2(ces_25_15_io_outs_2),
    .io_outs_3(ces_25_15_io_outs_3)
  );
  Element ces_25_16 ( // @[MockArray.scala 36:52]
    .clock(ces_25_16_clock),
    .io_ins_0(ces_25_16_io_ins_0),
    .io_ins_1(ces_25_16_io_ins_1),
    .io_ins_2(ces_25_16_io_ins_2),
    .io_ins_3(ces_25_16_io_ins_3),
    .io_outs_0(ces_25_16_io_outs_0),
    .io_outs_1(ces_25_16_io_outs_1),
    .io_outs_2(ces_25_16_io_outs_2),
    .io_outs_3(ces_25_16_io_outs_3)
  );
  Element ces_25_17 ( // @[MockArray.scala 36:52]
    .clock(ces_25_17_clock),
    .io_ins_0(ces_25_17_io_ins_0),
    .io_ins_1(ces_25_17_io_ins_1),
    .io_ins_2(ces_25_17_io_ins_2),
    .io_ins_3(ces_25_17_io_ins_3),
    .io_outs_0(ces_25_17_io_outs_0),
    .io_outs_1(ces_25_17_io_outs_1),
    .io_outs_2(ces_25_17_io_outs_2),
    .io_outs_3(ces_25_17_io_outs_3)
  );
  Element ces_25_18 ( // @[MockArray.scala 36:52]
    .clock(ces_25_18_clock),
    .io_ins_0(ces_25_18_io_ins_0),
    .io_ins_1(ces_25_18_io_ins_1),
    .io_ins_2(ces_25_18_io_ins_2),
    .io_ins_3(ces_25_18_io_ins_3),
    .io_outs_0(ces_25_18_io_outs_0),
    .io_outs_1(ces_25_18_io_outs_1),
    .io_outs_2(ces_25_18_io_outs_2),
    .io_outs_3(ces_25_18_io_outs_3)
  );
  Element ces_25_19 ( // @[MockArray.scala 36:52]
    .clock(ces_25_19_clock),
    .io_ins_0(ces_25_19_io_ins_0),
    .io_ins_1(ces_25_19_io_ins_1),
    .io_ins_2(ces_25_19_io_ins_2),
    .io_ins_3(ces_25_19_io_ins_3),
    .io_outs_0(ces_25_19_io_outs_0),
    .io_outs_1(ces_25_19_io_outs_1),
    .io_outs_2(ces_25_19_io_outs_2),
    .io_outs_3(ces_25_19_io_outs_3)
  );
  Element ces_25_20 ( // @[MockArray.scala 36:52]
    .clock(ces_25_20_clock),
    .io_ins_0(ces_25_20_io_ins_0),
    .io_ins_1(ces_25_20_io_ins_1),
    .io_ins_2(ces_25_20_io_ins_2),
    .io_ins_3(ces_25_20_io_ins_3),
    .io_outs_0(ces_25_20_io_outs_0),
    .io_outs_1(ces_25_20_io_outs_1),
    .io_outs_2(ces_25_20_io_outs_2),
    .io_outs_3(ces_25_20_io_outs_3)
  );
  Element ces_25_21 ( // @[MockArray.scala 36:52]
    .clock(ces_25_21_clock),
    .io_ins_0(ces_25_21_io_ins_0),
    .io_ins_1(ces_25_21_io_ins_1),
    .io_ins_2(ces_25_21_io_ins_2),
    .io_ins_3(ces_25_21_io_ins_3),
    .io_outs_0(ces_25_21_io_outs_0),
    .io_outs_1(ces_25_21_io_outs_1),
    .io_outs_2(ces_25_21_io_outs_2),
    .io_outs_3(ces_25_21_io_outs_3)
  );
  Element ces_25_22 ( // @[MockArray.scala 36:52]
    .clock(ces_25_22_clock),
    .io_ins_0(ces_25_22_io_ins_0),
    .io_ins_1(ces_25_22_io_ins_1),
    .io_ins_2(ces_25_22_io_ins_2),
    .io_ins_3(ces_25_22_io_ins_3),
    .io_outs_0(ces_25_22_io_outs_0),
    .io_outs_1(ces_25_22_io_outs_1),
    .io_outs_2(ces_25_22_io_outs_2),
    .io_outs_3(ces_25_22_io_outs_3)
  );
  Element ces_25_23 ( // @[MockArray.scala 36:52]
    .clock(ces_25_23_clock),
    .io_ins_0(ces_25_23_io_ins_0),
    .io_ins_1(ces_25_23_io_ins_1),
    .io_ins_2(ces_25_23_io_ins_2),
    .io_ins_3(ces_25_23_io_ins_3),
    .io_outs_0(ces_25_23_io_outs_0),
    .io_outs_1(ces_25_23_io_outs_1),
    .io_outs_2(ces_25_23_io_outs_2),
    .io_outs_3(ces_25_23_io_outs_3)
  );
  Element ces_25_24 ( // @[MockArray.scala 36:52]
    .clock(ces_25_24_clock),
    .io_ins_0(ces_25_24_io_ins_0),
    .io_ins_1(ces_25_24_io_ins_1),
    .io_ins_2(ces_25_24_io_ins_2),
    .io_ins_3(ces_25_24_io_ins_3),
    .io_outs_0(ces_25_24_io_outs_0),
    .io_outs_1(ces_25_24_io_outs_1),
    .io_outs_2(ces_25_24_io_outs_2),
    .io_outs_3(ces_25_24_io_outs_3)
  );
  Element ces_25_25 ( // @[MockArray.scala 36:52]
    .clock(ces_25_25_clock),
    .io_ins_0(ces_25_25_io_ins_0),
    .io_ins_1(ces_25_25_io_ins_1),
    .io_ins_2(ces_25_25_io_ins_2),
    .io_ins_3(ces_25_25_io_ins_3),
    .io_outs_0(ces_25_25_io_outs_0),
    .io_outs_1(ces_25_25_io_outs_1),
    .io_outs_2(ces_25_25_io_outs_2),
    .io_outs_3(ces_25_25_io_outs_3)
  );
  Element ces_25_26 ( // @[MockArray.scala 36:52]
    .clock(ces_25_26_clock),
    .io_ins_0(ces_25_26_io_ins_0),
    .io_ins_1(ces_25_26_io_ins_1),
    .io_ins_2(ces_25_26_io_ins_2),
    .io_ins_3(ces_25_26_io_ins_3),
    .io_outs_0(ces_25_26_io_outs_0),
    .io_outs_1(ces_25_26_io_outs_1),
    .io_outs_2(ces_25_26_io_outs_2),
    .io_outs_3(ces_25_26_io_outs_3)
  );
  Element ces_25_27 ( // @[MockArray.scala 36:52]
    .clock(ces_25_27_clock),
    .io_ins_0(ces_25_27_io_ins_0),
    .io_ins_1(ces_25_27_io_ins_1),
    .io_ins_2(ces_25_27_io_ins_2),
    .io_ins_3(ces_25_27_io_ins_3),
    .io_outs_0(ces_25_27_io_outs_0),
    .io_outs_1(ces_25_27_io_outs_1),
    .io_outs_2(ces_25_27_io_outs_2),
    .io_outs_3(ces_25_27_io_outs_3)
  );
  Element ces_25_28 ( // @[MockArray.scala 36:52]
    .clock(ces_25_28_clock),
    .io_ins_0(ces_25_28_io_ins_0),
    .io_ins_1(ces_25_28_io_ins_1),
    .io_ins_2(ces_25_28_io_ins_2),
    .io_ins_3(ces_25_28_io_ins_3),
    .io_outs_0(ces_25_28_io_outs_0),
    .io_outs_1(ces_25_28_io_outs_1),
    .io_outs_2(ces_25_28_io_outs_2),
    .io_outs_3(ces_25_28_io_outs_3)
  );
  Element ces_25_29 ( // @[MockArray.scala 36:52]
    .clock(ces_25_29_clock),
    .io_ins_0(ces_25_29_io_ins_0),
    .io_ins_1(ces_25_29_io_ins_1),
    .io_ins_2(ces_25_29_io_ins_2),
    .io_ins_3(ces_25_29_io_ins_3),
    .io_outs_0(ces_25_29_io_outs_0),
    .io_outs_1(ces_25_29_io_outs_1),
    .io_outs_2(ces_25_29_io_outs_2),
    .io_outs_3(ces_25_29_io_outs_3)
  );
  Element ces_25_30 ( // @[MockArray.scala 36:52]
    .clock(ces_25_30_clock),
    .io_ins_0(ces_25_30_io_ins_0),
    .io_ins_1(ces_25_30_io_ins_1),
    .io_ins_2(ces_25_30_io_ins_2),
    .io_ins_3(ces_25_30_io_ins_3),
    .io_outs_0(ces_25_30_io_outs_0),
    .io_outs_1(ces_25_30_io_outs_1),
    .io_outs_2(ces_25_30_io_outs_2),
    .io_outs_3(ces_25_30_io_outs_3)
  );
  Element ces_25_31 ( // @[MockArray.scala 36:52]
    .clock(ces_25_31_clock),
    .io_ins_0(ces_25_31_io_ins_0),
    .io_ins_1(ces_25_31_io_ins_1),
    .io_ins_2(ces_25_31_io_ins_2),
    .io_ins_3(ces_25_31_io_ins_3),
    .io_outs_0(ces_25_31_io_outs_0),
    .io_outs_1(ces_25_31_io_outs_1),
    .io_outs_2(ces_25_31_io_outs_2),
    .io_outs_3(ces_25_31_io_outs_3)
  );
  Element ces_26_0 ( // @[MockArray.scala 36:52]
    .clock(ces_26_0_clock),
    .io_ins_0(ces_26_0_io_ins_0),
    .io_ins_1(ces_26_0_io_ins_1),
    .io_ins_2(ces_26_0_io_ins_2),
    .io_ins_3(ces_26_0_io_ins_3),
    .io_outs_0(ces_26_0_io_outs_0),
    .io_outs_1(ces_26_0_io_outs_1),
    .io_outs_2(ces_26_0_io_outs_2),
    .io_outs_3(ces_26_0_io_outs_3)
  );
  Element ces_26_1 ( // @[MockArray.scala 36:52]
    .clock(ces_26_1_clock),
    .io_ins_0(ces_26_1_io_ins_0),
    .io_ins_1(ces_26_1_io_ins_1),
    .io_ins_2(ces_26_1_io_ins_2),
    .io_ins_3(ces_26_1_io_ins_3),
    .io_outs_0(ces_26_1_io_outs_0),
    .io_outs_1(ces_26_1_io_outs_1),
    .io_outs_2(ces_26_1_io_outs_2),
    .io_outs_3(ces_26_1_io_outs_3)
  );
  Element ces_26_2 ( // @[MockArray.scala 36:52]
    .clock(ces_26_2_clock),
    .io_ins_0(ces_26_2_io_ins_0),
    .io_ins_1(ces_26_2_io_ins_1),
    .io_ins_2(ces_26_2_io_ins_2),
    .io_ins_3(ces_26_2_io_ins_3),
    .io_outs_0(ces_26_2_io_outs_0),
    .io_outs_1(ces_26_2_io_outs_1),
    .io_outs_2(ces_26_2_io_outs_2),
    .io_outs_3(ces_26_2_io_outs_3)
  );
  Element ces_26_3 ( // @[MockArray.scala 36:52]
    .clock(ces_26_3_clock),
    .io_ins_0(ces_26_3_io_ins_0),
    .io_ins_1(ces_26_3_io_ins_1),
    .io_ins_2(ces_26_3_io_ins_2),
    .io_ins_3(ces_26_3_io_ins_3),
    .io_outs_0(ces_26_3_io_outs_0),
    .io_outs_1(ces_26_3_io_outs_1),
    .io_outs_2(ces_26_3_io_outs_2),
    .io_outs_3(ces_26_3_io_outs_3)
  );
  Element ces_26_4 ( // @[MockArray.scala 36:52]
    .clock(ces_26_4_clock),
    .io_ins_0(ces_26_4_io_ins_0),
    .io_ins_1(ces_26_4_io_ins_1),
    .io_ins_2(ces_26_4_io_ins_2),
    .io_ins_3(ces_26_4_io_ins_3),
    .io_outs_0(ces_26_4_io_outs_0),
    .io_outs_1(ces_26_4_io_outs_1),
    .io_outs_2(ces_26_4_io_outs_2),
    .io_outs_3(ces_26_4_io_outs_3)
  );
  Element ces_26_5 ( // @[MockArray.scala 36:52]
    .clock(ces_26_5_clock),
    .io_ins_0(ces_26_5_io_ins_0),
    .io_ins_1(ces_26_5_io_ins_1),
    .io_ins_2(ces_26_5_io_ins_2),
    .io_ins_3(ces_26_5_io_ins_3),
    .io_outs_0(ces_26_5_io_outs_0),
    .io_outs_1(ces_26_5_io_outs_1),
    .io_outs_2(ces_26_5_io_outs_2),
    .io_outs_3(ces_26_5_io_outs_3)
  );
  Element ces_26_6 ( // @[MockArray.scala 36:52]
    .clock(ces_26_6_clock),
    .io_ins_0(ces_26_6_io_ins_0),
    .io_ins_1(ces_26_6_io_ins_1),
    .io_ins_2(ces_26_6_io_ins_2),
    .io_ins_3(ces_26_6_io_ins_3),
    .io_outs_0(ces_26_6_io_outs_0),
    .io_outs_1(ces_26_6_io_outs_1),
    .io_outs_2(ces_26_6_io_outs_2),
    .io_outs_3(ces_26_6_io_outs_3)
  );
  Element ces_26_7 ( // @[MockArray.scala 36:52]
    .clock(ces_26_7_clock),
    .io_ins_0(ces_26_7_io_ins_0),
    .io_ins_1(ces_26_7_io_ins_1),
    .io_ins_2(ces_26_7_io_ins_2),
    .io_ins_3(ces_26_7_io_ins_3),
    .io_outs_0(ces_26_7_io_outs_0),
    .io_outs_1(ces_26_7_io_outs_1),
    .io_outs_2(ces_26_7_io_outs_2),
    .io_outs_3(ces_26_7_io_outs_3)
  );
  Element ces_26_8 ( // @[MockArray.scala 36:52]
    .clock(ces_26_8_clock),
    .io_ins_0(ces_26_8_io_ins_0),
    .io_ins_1(ces_26_8_io_ins_1),
    .io_ins_2(ces_26_8_io_ins_2),
    .io_ins_3(ces_26_8_io_ins_3),
    .io_outs_0(ces_26_8_io_outs_0),
    .io_outs_1(ces_26_8_io_outs_1),
    .io_outs_2(ces_26_8_io_outs_2),
    .io_outs_3(ces_26_8_io_outs_3)
  );
  Element ces_26_9 ( // @[MockArray.scala 36:52]
    .clock(ces_26_9_clock),
    .io_ins_0(ces_26_9_io_ins_0),
    .io_ins_1(ces_26_9_io_ins_1),
    .io_ins_2(ces_26_9_io_ins_2),
    .io_ins_3(ces_26_9_io_ins_3),
    .io_outs_0(ces_26_9_io_outs_0),
    .io_outs_1(ces_26_9_io_outs_1),
    .io_outs_2(ces_26_9_io_outs_2),
    .io_outs_3(ces_26_9_io_outs_3)
  );
  Element ces_26_10 ( // @[MockArray.scala 36:52]
    .clock(ces_26_10_clock),
    .io_ins_0(ces_26_10_io_ins_0),
    .io_ins_1(ces_26_10_io_ins_1),
    .io_ins_2(ces_26_10_io_ins_2),
    .io_ins_3(ces_26_10_io_ins_3),
    .io_outs_0(ces_26_10_io_outs_0),
    .io_outs_1(ces_26_10_io_outs_1),
    .io_outs_2(ces_26_10_io_outs_2),
    .io_outs_3(ces_26_10_io_outs_3)
  );
  Element ces_26_11 ( // @[MockArray.scala 36:52]
    .clock(ces_26_11_clock),
    .io_ins_0(ces_26_11_io_ins_0),
    .io_ins_1(ces_26_11_io_ins_1),
    .io_ins_2(ces_26_11_io_ins_2),
    .io_ins_3(ces_26_11_io_ins_3),
    .io_outs_0(ces_26_11_io_outs_0),
    .io_outs_1(ces_26_11_io_outs_1),
    .io_outs_2(ces_26_11_io_outs_2),
    .io_outs_3(ces_26_11_io_outs_3)
  );
  Element ces_26_12 ( // @[MockArray.scala 36:52]
    .clock(ces_26_12_clock),
    .io_ins_0(ces_26_12_io_ins_0),
    .io_ins_1(ces_26_12_io_ins_1),
    .io_ins_2(ces_26_12_io_ins_2),
    .io_ins_3(ces_26_12_io_ins_3),
    .io_outs_0(ces_26_12_io_outs_0),
    .io_outs_1(ces_26_12_io_outs_1),
    .io_outs_2(ces_26_12_io_outs_2),
    .io_outs_3(ces_26_12_io_outs_3)
  );
  Element ces_26_13 ( // @[MockArray.scala 36:52]
    .clock(ces_26_13_clock),
    .io_ins_0(ces_26_13_io_ins_0),
    .io_ins_1(ces_26_13_io_ins_1),
    .io_ins_2(ces_26_13_io_ins_2),
    .io_ins_3(ces_26_13_io_ins_3),
    .io_outs_0(ces_26_13_io_outs_0),
    .io_outs_1(ces_26_13_io_outs_1),
    .io_outs_2(ces_26_13_io_outs_2),
    .io_outs_3(ces_26_13_io_outs_3)
  );
  Element ces_26_14 ( // @[MockArray.scala 36:52]
    .clock(ces_26_14_clock),
    .io_ins_0(ces_26_14_io_ins_0),
    .io_ins_1(ces_26_14_io_ins_1),
    .io_ins_2(ces_26_14_io_ins_2),
    .io_ins_3(ces_26_14_io_ins_3),
    .io_outs_0(ces_26_14_io_outs_0),
    .io_outs_1(ces_26_14_io_outs_1),
    .io_outs_2(ces_26_14_io_outs_2),
    .io_outs_3(ces_26_14_io_outs_3)
  );
  Element ces_26_15 ( // @[MockArray.scala 36:52]
    .clock(ces_26_15_clock),
    .io_ins_0(ces_26_15_io_ins_0),
    .io_ins_1(ces_26_15_io_ins_1),
    .io_ins_2(ces_26_15_io_ins_2),
    .io_ins_3(ces_26_15_io_ins_3),
    .io_outs_0(ces_26_15_io_outs_0),
    .io_outs_1(ces_26_15_io_outs_1),
    .io_outs_2(ces_26_15_io_outs_2),
    .io_outs_3(ces_26_15_io_outs_3)
  );
  Element ces_26_16 ( // @[MockArray.scala 36:52]
    .clock(ces_26_16_clock),
    .io_ins_0(ces_26_16_io_ins_0),
    .io_ins_1(ces_26_16_io_ins_1),
    .io_ins_2(ces_26_16_io_ins_2),
    .io_ins_3(ces_26_16_io_ins_3),
    .io_outs_0(ces_26_16_io_outs_0),
    .io_outs_1(ces_26_16_io_outs_1),
    .io_outs_2(ces_26_16_io_outs_2),
    .io_outs_3(ces_26_16_io_outs_3)
  );
  Element ces_26_17 ( // @[MockArray.scala 36:52]
    .clock(ces_26_17_clock),
    .io_ins_0(ces_26_17_io_ins_0),
    .io_ins_1(ces_26_17_io_ins_1),
    .io_ins_2(ces_26_17_io_ins_2),
    .io_ins_3(ces_26_17_io_ins_3),
    .io_outs_0(ces_26_17_io_outs_0),
    .io_outs_1(ces_26_17_io_outs_1),
    .io_outs_2(ces_26_17_io_outs_2),
    .io_outs_3(ces_26_17_io_outs_3)
  );
  Element ces_26_18 ( // @[MockArray.scala 36:52]
    .clock(ces_26_18_clock),
    .io_ins_0(ces_26_18_io_ins_0),
    .io_ins_1(ces_26_18_io_ins_1),
    .io_ins_2(ces_26_18_io_ins_2),
    .io_ins_3(ces_26_18_io_ins_3),
    .io_outs_0(ces_26_18_io_outs_0),
    .io_outs_1(ces_26_18_io_outs_1),
    .io_outs_2(ces_26_18_io_outs_2),
    .io_outs_3(ces_26_18_io_outs_3)
  );
  Element ces_26_19 ( // @[MockArray.scala 36:52]
    .clock(ces_26_19_clock),
    .io_ins_0(ces_26_19_io_ins_0),
    .io_ins_1(ces_26_19_io_ins_1),
    .io_ins_2(ces_26_19_io_ins_2),
    .io_ins_3(ces_26_19_io_ins_3),
    .io_outs_0(ces_26_19_io_outs_0),
    .io_outs_1(ces_26_19_io_outs_1),
    .io_outs_2(ces_26_19_io_outs_2),
    .io_outs_3(ces_26_19_io_outs_3)
  );
  Element ces_26_20 ( // @[MockArray.scala 36:52]
    .clock(ces_26_20_clock),
    .io_ins_0(ces_26_20_io_ins_0),
    .io_ins_1(ces_26_20_io_ins_1),
    .io_ins_2(ces_26_20_io_ins_2),
    .io_ins_3(ces_26_20_io_ins_3),
    .io_outs_0(ces_26_20_io_outs_0),
    .io_outs_1(ces_26_20_io_outs_1),
    .io_outs_2(ces_26_20_io_outs_2),
    .io_outs_3(ces_26_20_io_outs_3)
  );
  Element ces_26_21 ( // @[MockArray.scala 36:52]
    .clock(ces_26_21_clock),
    .io_ins_0(ces_26_21_io_ins_0),
    .io_ins_1(ces_26_21_io_ins_1),
    .io_ins_2(ces_26_21_io_ins_2),
    .io_ins_3(ces_26_21_io_ins_3),
    .io_outs_0(ces_26_21_io_outs_0),
    .io_outs_1(ces_26_21_io_outs_1),
    .io_outs_2(ces_26_21_io_outs_2),
    .io_outs_3(ces_26_21_io_outs_3)
  );
  Element ces_26_22 ( // @[MockArray.scala 36:52]
    .clock(ces_26_22_clock),
    .io_ins_0(ces_26_22_io_ins_0),
    .io_ins_1(ces_26_22_io_ins_1),
    .io_ins_2(ces_26_22_io_ins_2),
    .io_ins_3(ces_26_22_io_ins_3),
    .io_outs_0(ces_26_22_io_outs_0),
    .io_outs_1(ces_26_22_io_outs_1),
    .io_outs_2(ces_26_22_io_outs_2),
    .io_outs_3(ces_26_22_io_outs_3)
  );
  Element ces_26_23 ( // @[MockArray.scala 36:52]
    .clock(ces_26_23_clock),
    .io_ins_0(ces_26_23_io_ins_0),
    .io_ins_1(ces_26_23_io_ins_1),
    .io_ins_2(ces_26_23_io_ins_2),
    .io_ins_3(ces_26_23_io_ins_3),
    .io_outs_0(ces_26_23_io_outs_0),
    .io_outs_1(ces_26_23_io_outs_1),
    .io_outs_2(ces_26_23_io_outs_2),
    .io_outs_3(ces_26_23_io_outs_3)
  );
  Element ces_26_24 ( // @[MockArray.scala 36:52]
    .clock(ces_26_24_clock),
    .io_ins_0(ces_26_24_io_ins_0),
    .io_ins_1(ces_26_24_io_ins_1),
    .io_ins_2(ces_26_24_io_ins_2),
    .io_ins_3(ces_26_24_io_ins_3),
    .io_outs_0(ces_26_24_io_outs_0),
    .io_outs_1(ces_26_24_io_outs_1),
    .io_outs_2(ces_26_24_io_outs_2),
    .io_outs_3(ces_26_24_io_outs_3)
  );
  Element ces_26_25 ( // @[MockArray.scala 36:52]
    .clock(ces_26_25_clock),
    .io_ins_0(ces_26_25_io_ins_0),
    .io_ins_1(ces_26_25_io_ins_1),
    .io_ins_2(ces_26_25_io_ins_2),
    .io_ins_3(ces_26_25_io_ins_3),
    .io_outs_0(ces_26_25_io_outs_0),
    .io_outs_1(ces_26_25_io_outs_1),
    .io_outs_2(ces_26_25_io_outs_2),
    .io_outs_3(ces_26_25_io_outs_3)
  );
  Element ces_26_26 ( // @[MockArray.scala 36:52]
    .clock(ces_26_26_clock),
    .io_ins_0(ces_26_26_io_ins_0),
    .io_ins_1(ces_26_26_io_ins_1),
    .io_ins_2(ces_26_26_io_ins_2),
    .io_ins_3(ces_26_26_io_ins_3),
    .io_outs_0(ces_26_26_io_outs_0),
    .io_outs_1(ces_26_26_io_outs_1),
    .io_outs_2(ces_26_26_io_outs_2),
    .io_outs_3(ces_26_26_io_outs_3)
  );
  Element ces_26_27 ( // @[MockArray.scala 36:52]
    .clock(ces_26_27_clock),
    .io_ins_0(ces_26_27_io_ins_0),
    .io_ins_1(ces_26_27_io_ins_1),
    .io_ins_2(ces_26_27_io_ins_2),
    .io_ins_3(ces_26_27_io_ins_3),
    .io_outs_0(ces_26_27_io_outs_0),
    .io_outs_1(ces_26_27_io_outs_1),
    .io_outs_2(ces_26_27_io_outs_2),
    .io_outs_3(ces_26_27_io_outs_3)
  );
  Element ces_26_28 ( // @[MockArray.scala 36:52]
    .clock(ces_26_28_clock),
    .io_ins_0(ces_26_28_io_ins_0),
    .io_ins_1(ces_26_28_io_ins_1),
    .io_ins_2(ces_26_28_io_ins_2),
    .io_ins_3(ces_26_28_io_ins_3),
    .io_outs_0(ces_26_28_io_outs_0),
    .io_outs_1(ces_26_28_io_outs_1),
    .io_outs_2(ces_26_28_io_outs_2),
    .io_outs_3(ces_26_28_io_outs_3)
  );
  Element ces_26_29 ( // @[MockArray.scala 36:52]
    .clock(ces_26_29_clock),
    .io_ins_0(ces_26_29_io_ins_0),
    .io_ins_1(ces_26_29_io_ins_1),
    .io_ins_2(ces_26_29_io_ins_2),
    .io_ins_3(ces_26_29_io_ins_3),
    .io_outs_0(ces_26_29_io_outs_0),
    .io_outs_1(ces_26_29_io_outs_1),
    .io_outs_2(ces_26_29_io_outs_2),
    .io_outs_3(ces_26_29_io_outs_3)
  );
  Element ces_26_30 ( // @[MockArray.scala 36:52]
    .clock(ces_26_30_clock),
    .io_ins_0(ces_26_30_io_ins_0),
    .io_ins_1(ces_26_30_io_ins_1),
    .io_ins_2(ces_26_30_io_ins_2),
    .io_ins_3(ces_26_30_io_ins_3),
    .io_outs_0(ces_26_30_io_outs_0),
    .io_outs_1(ces_26_30_io_outs_1),
    .io_outs_2(ces_26_30_io_outs_2),
    .io_outs_3(ces_26_30_io_outs_3)
  );
  Element ces_26_31 ( // @[MockArray.scala 36:52]
    .clock(ces_26_31_clock),
    .io_ins_0(ces_26_31_io_ins_0),
    .io_ins_1(ces_26_31_io_ins_1),
    .io_ins_2(ces_26_31_io_ins_2),
    .io_ins_3(ces_26_31_io_ins_3),
    .io_outs_0(ces_26_31_io_outs_0),
    .io_outs_1(ces_26_31_io_outs_1),
    .io_outs_2(ces_26_31_io_outs_2),
    .io_outs_3(ces_26_31_io_outs_3)
  );
  Element ces_27_0 ( // @[MockArray.scala 36:52]
    .clock(ces_27_0_clock),
    .io_ins_0(ces_27_0_io_ins_0),
    .io_ins_1(ces_27_0_io_ins_1),
    .io_ins_2(ces_27_0_io_ins_2),
    .io_ins_3(ces_27_0_io_ins_3),
    .io_outs_0(ces_27_0_io_outs_0),
    .io_outs_1(ces_27_0_io_outs_1),
    .io_outs_2(ces_27_0_io_outs_2),
    .io_outs_3(ces_27_0_io_outs_3)
  );
  Element ces_27_1 ( // @[MockArray.scala 36:52]
    .clock(ces_27_1_clock),
    .io_ins_0(ces_27_1_io_ins_0),
    .io_ins_1(ces_27_1_io_ins_1),
    .io_ins_2(ces_27_1_io_ins_2),
    .io_ins_3(ces_27_1_io_ins_3),
    .io_outs_0(ces_27_1_io_outs_0),
    .io_outs_1(ces_27_1_io_outs_1),
    .io_outs_2(ces_27_1_io_outs_2),
    .io_outs_3(ces_27_1_io_outs_3)
  );
  Element ces_27_2 ( // @[MockArray.scala 36:52]
    .clock(ces_27_2_clock),
    .io_ins_0(ces_27_2_io_ins_0),
    .io_ins_1(ces_27_2_io_ins_1),
    .io_ins_2(ces_27_2_io_ins_2),
    .io_ins_3(ces_27_2_io_ins_3),
    .io_outs_0(ces_27_2_io_outs_0),
    .io_outs_1(ces_27_2_io_outs_1),
    .io_outs_2(ces_27_2_io_outs_2),
    .io_outs_3(ces_27_2_io_outs_3)
  );
  Element ces_27_3 ( // @[MockArray.scala 36:52]
    .clock(ces_27_3_clock),
    .io_ins_0(ces_27_3_io_ins_0),
    .io_ins_1(ces_27_3_io_ins_1),
    .io_ins_2(ces_27_3_io_ins_2),
    .io_ins_3(ces_27_3_io_ins_3),
    .io_outs_0(ces_27_3_io_outs_0),
    .io_outs_1(ces_27_3_io_outs_1),
    .io_outs_2(ces_27_3_io_outs_2),
    .io_outs_3(ces_27_3_io_outs_3)
  );
  Element ces_27_4 ( // @[MockArray.scala 36:52]
    .clock(ces_27_4_clock),
    .io_ins_0(ces_27_4_io_ins_0),
    .io_ins_1(ces_27_4_io_ins_1),
    .io_ins_2(ces_27_4_io_ins_2),
    .io_ins_3(ces_27_4_io_ins_3),
    .io_outs_0(ces_27_4_io_outs_0),
    .io_outs_1(ces_27_4_io_outs_1),
    .io_outs_2(ces_27_4_io_outs_2),
    .io_outs_3(ces_27_4_io_outs_3)
  );
  Element ces_27_5 ( // @[MockArray.scala 36:52]
    .clock(ces_27_5_clock),
    .io_ins_0(ces_27_5_io_ins_0),
    .io_ins_1(ces_27_5_io_ins_1),
    .io_ins_2(ces_27_5_io_ins_2),
    .io_ins_3(ces_27_5_io_ins_3),
    .io_outs_0(ces_27_5_io_outs_0),
    .io_outs_1(ces_27_5_io_outs_1),
    .io_outs_2(ces_27_5_io_outs_2),
    .io_outs_3(ces_27_5_io_outs_3)
  );
  Element ces_27_6 ( // @[MockArray.scala 36:52]
    .clock(ces_27_6_clock),
    .io_ins_0(ces_27_6_io_ins_0),
    .io_ins_1(ces_27_6_io_ins_1),
    .io_ins_2(ces_27_6_io_ins_2),
    .io_ins_3(ces_27_6_io_ins_3),
    .io_outs_0(ces_27_6_io_outs_0),
    .io_outs_1(ces_27_6_io_outs_1),
    .io_outs_2(ces_27_6_io_outs_2),
    .io_outs_3(ces_27_6_io_outs_3)
  );
  Element ces_27_7 ( // @[MockArray.scala 36:52]
    .clock(ces_27_7_clock),
    .io_ins_0(ces_27_7_io_ins_0),
    .io_ins_1(ces_27_7_io_ins_1),
    .io_ins_2(ces_27_7_io_ins_2),
    .io_ins_3(ces_27_7_io_ins_3),
    .io_outs_0(ces_27_7_io_outs_0),
    .io_outs_1(ces_27_7_io_outs_1),
    .io_outs_2(ces_27_7_io_outs_2),
    .io_outs_3(ces_27_7_io_outs_3)
  );
  Element ces_27_8 ( // @[MockArray.scala 36:52]
    .clock(ces_27_8_clock),
    .io_ins_0(ces_27_8_io_ins_0),
    .io_ins_1(ces_27_8_io_ins_1),
    .io_ins_2(ces_27_8_io_ins_2),
    .io_ins_3(ces_27_8_io_ins_3),
    .io_outs_0(ces_27_8_io_outs_0),
    .io_outs_1(ces_27_8_io_outs_1),
    .io_outs_2(ces_27_8_io_outs_2),
    .io_outs_3(ces_27_8_io_outs_3)
  );
  Element ces_27_9 ( // @[MockArray.scala 36:52]
    .clock(ces_27_9_clock),
    .io_ins_0(ces_27_9_io_ins_0),
    .io_ins_1(ces_27_9_io_ins_1),
    .io_ins_2(ces_27_9_io_ins_2),
    .io_ins_3(ces_27_9_io_ins_3),
    .io_outs_0(ces_27_9_io_outs_0),
    .io_outs_1(ces_27_9_io_outs_1),
    .io_outs_2(ces_27_9_io_outs_2),
    .io_outs_3(ces_27_9_io_outs_3)
  );
  Element ces_27_10 ( // @[MockArray.scala 36:52]
    .clock(ces_27_10_clock),
    .io_ins_0(ces_27_10_io_ins_0),
    .io_ins_1(ces_27_10_io_ins_1),
    .io_ins_2(ces_27_10_io_ins_2),
    .io_ins_3(ces_27_10_io_ins_3),
    .io_outs_0(ces_27_10_io_outs_0),
    .io_outs_1(ces_27_10_io_outs_1),
    .io_outs_2(ces_27_10_io_outs_2),
    .io_outs_3(ces_27_10_io_outs_3)
  );
  Element ces_27_11 ( // @[MockArray.scala 36:52]
    .clock(ces_27_11_clock),
    .io_ins_0(ces_27_11_io_ins_0),
    .io_ins_1(ces_27_11_io_ins_1),
    .io_ins_2(ces_27_11_io_ins_2),
    .io_ins_3(ces_27_11_io_ins_3),
    .io_outs_0(ces_27_11_io_outs_0),
    .io_outs_1(ces_27_11_io_outs_1),
    .io_outs_2(ces_27_11_io_outs_2),
    .io_outs_3(ces_27_11_io_outs_3)
  );
  Element ces_27_12 ( // @[MockArray.scala 36:52]
    .clock(ces_27_12_clock),
    .io_ins_0(ces_27_12_io_ins_0),
    .io_ins_1(ces_27_12_io_ins_1),
    .io_ins_2(ces_27_12_io_ins_2),
    .io_ins_3(ces_27_12_io_ins_3),
    .io_outs_0(ces_27_12_io_outs_0),
    .io_outs_1(ces_27_12_io_outs_1),
    .io_outs_2(ces_27_12_io_outs_2),
    .io_outs_3(ces_27_12_io_outs_3)
  );
  Element ces_27_13 ( // @[MockArray.scala 36:52]
    .clock(ces_27_13_clock),
    .io_ins_0(ces_27_13_io_ins_0),
    .io_ins_1(ces_27_13_io_ins_1),
    .io_ins_2(ces_27_13_io_ins_2),
    .io_ins_3(ces_27_13_io_ins_3),
    .io_outs_0(ces_27_13_io_outs_0),
    .io_outs_1(ces_27_13_io_outs_1),
    .io_outs_2(ces_27_13_io_outs_2),
    .io_outs_3(ces_27_13_io_outs_3)
  );
  Element ces_27_14 ( // @[MockArray.scala 36:52]
    .clock(ces_27_14_clock),
    .io_ins_0(ces_27_14_io_ins_0),
    .io_ins_1(ces_27_14_io_ins_1),
    .io_ins_2(ces_27_14_io_ins_2),
    .io_ins_3(ces_27_14_io_ins_3),
    .io_outs_0(ces_27_14_io_outs_0),
    .io_outs_1(ces_27_14_io_outs_1),
    .io_outs_2(ces_27_14_io_outs_2),
    .io_outs_3(ces_27_14_io_outs_3)
  );
  Element ces_27_15 ( // @[MockArray.scala 36:52]
    .clock(ces_27_15_clock),
    .io_ins_0(ces_27_15_io_ins_0),
    .io_ins_1(ces_27_15_io_ins_1),
    .io_ins_2(ces_27_15_io_ins_2),
    .io_ins_3(ces_27_15_io_ins_3),
    .io_outs_0(ces_27_15_io_outs_0),
    .io_outs_1(ces_27_15_io_outs_1),
    .io_outs_2(ces_27_15_io_outs_2),
    .io_outs_3(ces_27_15_io_outs_3)
  );
  Element ces_27_16 ( // @[MockArray.scala 36:52]
    .clock(ces_27_16_clock),
    .io_ins_0(ces_27_16_io_ins_0),
    .io_ins_1(ces_27_16_io_ins_1),
    .io_ins_2(ces_27_16_io_ins_2),
    .io_ins_3(ces_27_16_io_ins_3),
    .io_outs_0(ces_27_16_io_outs_0),
    .io_outs_1(ces_27_16_io_outs_1),
    .io_outs_2(ces_27_16_io_outs_2),
    .io_outs_3(ces_27_16_io_outs_3)
  );
  Element ces_27_17 ( // @[MockArray.scala 36:52]
    .clock(ces_27_17_clock),
    .io_ins_0(ces_27_17_io_ins_0),
    .io_ins_1(ces_27_17_io_ins_1),
    .io_ins_2(ces_27_17_io_ins_2),
    .io_ins_3(ces_27_17_io_ins_3),
    .io_outs_0(ces_27_17_io_outs_0),
    .io_outs_1(ces_27_17_io_outs_1),
    .io_outs_2(ces_27_17_io_outs_2),
    .io_outs_3(ces_27_17_io_outs_3)
  );
  Element ces_27_18 ( // @[MockArray.scala 36:52]
    .clock(ces_27_18_clock),
    .io_ins_0(ces_27_18_io_ins_0),
    .io_ins_1(ces_27_18_io_ins_1),
    .io_ins_2(ces_27_18_io_ins_2),
    .io_ins_3(ces_27_18_io_ins_3),
    .io_outs_0(ces_27_18_io_outs_0),
    .io_outs_1(ces_27_18_io_outs_1),
    .io_outs_2(ces_27_18_io_outs_2),
    .io_outs_3(ces_27_18_io_outs_3)
  );
  Element ces_27_19 ( // @[MockArray.scala 36:52]
    .clock(ces_27_19_clock),
    .io_ins_0(ces_27_19_io_ins_0),
    .io_ins_1(ces_27_19_io_ins_1),
    .io_ins_2(ces_27_19_io_ins_2),
    .io_ins_3(ces_27_19_io_ins_3),
    .io_outs_0(ces_27_19_io_outs_0),
    .io_outs_1(ces_27_19_io_outs_1),
    .io_outs_2(ces_27_19_io_outs_2),
    .io_outs_3(ces_27_19_io_outs_3)
  );
  Element ces_27_20 ( // @[MockArray.scala 36:52]
    .clock(ces_27_20_clock),
    .io_ins_0(ces_27_20_io_ins_0),
    .io_ins_1(ces_27_20_io_ins_1),
    .io_ins_2(ces_27_20_io_ins_2),
    .io_ins_3(ces_27_20_io_ins_3),
    .io_outs_0(ces_27_20_io_outs_0),
    .io_outs_1(ces_27_20_io_outs_1),
    .io_outs_2(ces_27_20_io_outs_2),
    .io_outs_3(ces_27_20_io_outs_3)
  );
  Element ces_27_21 ( // @[MockArray.scala 36:52]
    .clock(ces_27_21_clock),
    .io_ins_0(ces_27_21_io_ins_0),
    .io_ins_1(ces_27_21_io_ins_1),
    .io_ins_2(ces_27_21_io_ins_2),
    .io_ins_3(ces_27_21_io_ins_3),
    .io_outs_0(ces_27_21_io_outs_0),
    .io_outs_1(ces_27_21_io_outs_1),
    .io_outs_2(ces_27_21_io_outs_2),
    .io_outs_3(ces_27_21_io_outs_3)
  );
  Element ces_27_22 ( // @[MockArray.scala 36:52]
    .clock(ces_27_22_clock),
    .io_ins_0(ces_27_22_io_ins_0),
    .io_ins_1(ces_27_22_io_ins_1),
    .io_ins_2(ces_27_22_io_ins_2),
    .io_ins_3(ces_27_22_io_ins_3),
    .io_outs_0(ces_27_22_io_outs_0),
    .io_outs_1(ces_27_22_io_outs_1),
    .io_outs_2(ces_27_22_io_outs_2),
    .io_outs_3(ces_27_22_io_outs_3)
  );
  Element ces_27_23 ( // @[MockArray.scala 36:52]
    .clock(ces_27_23_clock),
    .io_ins_0(ces_27_23_io_ins_0),
    .io_ins_1(ces_27_23_io_ins_1),
    .io_ins_2(ces_27_23_io_ins_2),
    .io_ins_3(ces_27_23_io_ins_3),
    .io_outs_0(ces_27_23_io_outs_0),
    .io_outs_1(ces_27_23_io_outs_1),
    .io_outs_2(ces_27_23_io_outs_2),
    .io_outs_3(ces_27_23_io_outs_3)
  );
  Element ces_27_24 ( // @[MockArray.scala 36:52]
    .clock(ces_27_24_clock),
    .io_ins_0(ces_27_24_io_ins_0),
    .io_ins_1(ces_27_24_io_ins_1),
    .io_ins_2(ces_27_24_io_ins_2),
    .io_ins_3(ces_27_24_io_ins_3),
    .io_outs_0(ces_27_24_io_outs_0),
    .io_outs_1(ces_27_24_io_outs_1),
    .io_outs_2(ces_27_24_io_outs_2),
    .io_outs_3(ces_27_24_io_outs_3)
  );
  Element ces_27_25 ( // @[MockArray.scala 36:52]
    .clock(ces_27_25_clock),
    .io_ins_0(ces_27_25_io_ins_0),
    .io_ins_1(ces_27_25_io_ins_1),
    .io_ins_2(ces_27_25_io_ins_2),
    .io_ins_3(ces_27_25_io_ins_3),
    .io_outs_0(ces_27_25_io_outs_0),
    .io_outs_1(ces_27_25_io_outs_1),
    .io_outs_2(ces_27_25_io_outs_2),
    .io_outs_3(ces_27_25_io_outs_3)
  );
  Element ces_27_26 ( // @[MockArray.scala 36:52]
    .clock(ces_27_26_clock),
    .io_ins_0(ces_27_26_io_ins_0),
    .io_ins_1(ces_27_26_io_ins_1),
    .io_ins_2(ces_27_26_io_ins_2),
    .io_ins_3(ces_27_26_io_ins_3),
    .io_outs_0(ces_27_26_io_outs_0),
    .io_outs_1(ces_27_26_io_outs_1),
    .io_outs_2(ces_27_26_io_outs_2),
    .io_outs_3(ces_27_26_io_outs_3)
  );
  Element ces_27_27 ( // @[MockArray.scala 36:52]
    .clock(ces_27_27_clock),
    .io_ins_0(ces_27_27_io_ins_0),
    .io_ins_1(ces_27_27_io_ins_1),
    .io_ins_2(ces_27_27_io_ins_2),
    .io_ins_3(ces_27_27_io_ins_3),
    .io_outs_0(ces_27_27_io_outs_0),
    .io_outs_1(ces_27_27_io_outs_1),
    .io_outs_2(ces_27_27_io_outs_2),
    .io_outs_3(ces_27_27_io_outs_3)
  );
  Element ces_27_28 ( // @[MockArray.scala 36:52]
    .clock(ces_27_28_clock),
    .io_ins_0(ces_27_28_io_ins_0),
    .io_ins_1(ces_27_28_io_ins_1),
    .io_ins_2(ces_27_28_io_ins_2),
    .io_ins_3(ces_27_28_io_ins_3),
    .io_outs_0(ces_27_28_io_outs_0),
    .io_outs_1(ces_27_28_io_outs_1),
    .io_outs_2(ces_27_28_io_outs_2),
    .io_outs_3(ces_27_28_io_outs_3)
  );
  Element ces_27_29 ( // @[MockArray.scala 36:52]
    .clock(ces_27_29_clock),
    .io_ins_0(ces_27_29_io_ins_0),
    .io_ins_1(ces_27_29_io_ins_1),
    .io_ins_2(ces_27_29_io_ins_2),
    .io_ins_3(ces_27_29_io_ins_3),
    .io_outs_0(ces_27_29_io_outs_0),
    .io_outs_1(ces_27_29_io_outs_1),
    .io_outs_2(ces_27_29_io_outs_2),
    .io_outs_3(ces_27_29_io_outs_3)
  );
  Element ces_27_30 ( // @[MockArray.scala 36:52]
    .clock(ces_27_30_clock),
    .io_ins_0(ces_27_30_io_ins_0),
    .io_ins_1(ces_27_30_io_ins_1),
    .io_ins_2(ces_27_30_io_ins_2),
    .io_ins_3(ces_27_30_io_ins_3),
    .io_outs_0(ces_27_30_io_outs_0),
    .io_outs_1(ces_27_30_io_outs_1),
    .io_outs_2(ces_27_30_io_outs_2),
    .io_outs_3(ces_27_30_io_outs_3)
  );
  Element ces_27_31 ( // @[MockArray.scala 36:52]
    .clock(ces_27_31_clock),
    .io_ins_0(ces_27_31_io_ins_0),
    .io_ins_1(ces_27_31_io_ins_1),
    .io_ins_2(ces_27_31_io_ins_2),
    .io_ins_3(ces_27_31_io_ins_3),
    .io_outs_0(ces_27_31_io_outs_0),
    .io_outs_1(ces_27_31_io_outs_1),
    .io_outs_2(ces_27_31_io_outs_2),
    .io_outs_3(ces_27_31_io_outs_3)
  );
  Element ces_28_0 ( // @[MockArray.scala 36:52]
    .clock(ces_28_0_clock),
    .io_ins_0(ces_28_0_io_ins_0),
    .io_ins_1(ces_28_0_io_ins_1),
    .io_ins_2(ces_28_0_io_ins_2),
    .io_ins_3(ces_28_0_io_ins_3),
    .io_outs_0(ces_28_0_io_outs_0),
    .io_outs_1(ces_28_0_io_outs_1),
    .io_outs_2(ces_28_0_io_outs_2),
    .io_outs_3(ces_28_0_io_outs_3)
  );
  Element ces_28_1 ( // @[MockArray.scala 36:52]
    .clock(ces_28_1_clock),
    .io_ins_0(ces_28_1_io_ins_0),
    .io_ins_1(ces_28_1_io_ins_1),
    .io_ins_2(ces_28_1_io_ins_2),
    .io_ins_3(ces_28_1_io_ins_3),
    .io_outs_0(ces_28_1_io_outs_0),
    .io_outs_1(ces_28_1_io_outs_1),
    .io_outs_2(ces_28_1_io_outs_2),
    .io_outs_3(ces_28_1_io_outs_3)
  );
  Element ces_28_2 ( // @[MockArray.scala 36:52]
    .clock(ces_28_2_clock),
    .io_ins_0(ces_28_2_io_ins_0),
    .io_ins_1(ces_28_2_io_ins_1),
    .io_ins_2(ces_28_2_io_ins_2),
    .io_ins_3(ces_28_2_io_ins_3),
    .io_outs_0(ces_28_2_io_outs_0),
    .io_outs_1(ces_28_2_io_outs_1),
    .io_outs_2(ces_28_2_io_outs_2),
    .io_outs_3(ces_28_2_io_outs_3)
  );
  Element ces_28_3 ( // @[MockArray.scala 36:52]
    .clock(ces_28_3_clock),
    .io_ins_0(ces_28_3_io_ins_0),
    .io_ins_1(ces_28_3_io_ins_1),
    .io_ins_2(ces_28_3_io_ins_2),
    .io_ins_3(ces_28_3_io_ins_3),
    .io_outs_0(ces_28_3_io_outs_0),
    .io_outs_1(ces_28_3_io_outs_1),
    .io_outs_2(ces_28_3_io_outs_2),
    .io_outs_3(ces_28_3_io_outs_3)
  );
  Element ces_28_4 ( // @[MockArray.scala 36:52]
    .clock(ces_28_4_clock),
    .io_ins_0(ces_28_4_io_ins_0),
    .io_ins_1(ces_28_4_io_ins_1),
    .io_ins_2(ces_28_4_io_ins_2),
    .io_ins_3(ces_28_4_io_ins_3),
    .io_outs_0(ces_28_4_io_outs_0),
    .io_outs_1(ces_28_4_io_outs_1),
    .io_outs_2(ces_28_4_io_outs_2),
    .io_outs_3(ces_28_4_io_outs_3)
  );
  Element ces_28_5 ( // @[MockArray.scala 36:52]
    .clock(ces_28_5_clock),
    .io_ins_0(ces_28_5_io_ins_0),
    .io_ins_1(ces_28_5_io_ins_1),
    .io_ins_2(ces_28_5_io_ins_2),
    .io_ins_3(ces_28_5_io_ins_3),
    .io_outs_0(ces_28_5_io_outs_0),
    .io_outs_1(ces_28_5_io_outs_1),
    .io_outs_2(ces_28_5_io_outs_2),
    .io_outs_3(ces_28_5_io_outs_3)
  );
  Element ces_28_6 ( // @[MockArray.scala 36:52]
    .clock(ces_28_6_clock),
    .io_ins_0(ces_28_6_io_ins_0),
    .io_ins_1(ces_28_6_io_ins_1),
    .io_ins_2(ces_28_6_io_ins_2),
    .io_ins_3(ces_28_6_io_ins_3),
    .io_outs_0(ces_28_6_io_outs_0),
    .io_outs_1(ces_28_6_io_outs_1),
    .io_outs_2(ces_28_6_io_outs_2),
    .io_outs_3(ces_28_6_io_outs_3)
  );
  Element ces_28_7 ( // @[MockArray.scala 36:52]
    .clock(ces_28_7_clock),
    .io_ins_0(ces_28_7_io_ins_0),
    .io_ins_1(ces_28_7_io_ins_1),
    .io_ins_2(ces_28_7_io_ins_2),
    .io_ins_3(ces_28_7_io_ins_3),
    .io_outs_0(ces_28_7_io_outs_0),
    .io_outs_1(ces_28_7_io_outs_1),
    .io_outs_2(ces_28_7_io_outs_2),
    .io_outs_3(ces_28_7_io_outs_3)
  );
  Element ces_28_8 ( // @[MockArray.scala 36:52]
    .clock(ces_28_8_clock),
    .io_ins_0(ces_28_8_io_ins_0),
    .io_ins_1(ces_28_8_io_ins_1),
    .io_ins_2(ces_28_8_io_ins_2),
    .io_ins_3(ces_28_8_io_ins_3),
    .io_outs_0(ces_28_8_io_outs_0),
    .io_outs_1(ces_28_8_io_outs_1),
    .io_outs_2(ces_28_8_io_outs_2),
    .io_outs_3(ces_28_8_io_outs_3)
  );
  Element ces_28_9 ( // @[MockArray.scala 36:52]
    .clock(ces_28_9_clock),
    .io_ins_0(ces_28_9_io_ins_0),
    .io_ins_1(ces_28_9_io_ins_1),
    .io_ins_2(ces_28_9_io_ins_2),
    .io_ins_3(ces_28_9_io_ins_3),
    .io_outs_0(ces_28_9_io_outs_0),
    .io_outs_1(ces_28_9_io_outs_1),
    .io_outs_2(ces_28_9_io_outs_2),
    .io_outs_3(ces_28_9_io_outs_3)
  );
  Element ces_28_10 ( // @[MockArray.scala 36:52]
    .clock(ces_28_10_clock),
    .io_ins_0(ces_28_10_io_ins_0),
    .io_ins_1(ces_28_10_io_ins_1),
    .io_ins_2(ces_28_10_io_ins_2),
    .io_ins_3(ces_28_10_io_ins_3),
    .io_outs_0(ces_28_10_io_outs_0),
    .io_outs_1(ces_28_10_io_outs_1),
    .io_outs_2(ces_28_10_io_outs_2),
    .io_outs_3(ces_28_10_io_outs_3)
  );
  Element ces_28_11 ( // @[MockArray.scala 36:52]
    .clock(ces_28_11_clock),
    .io_ins_0(ces_28_11_io_ins_0),
    .io_ins_1(ces_28_11_io_ins_1),
    .io_ins_2(ces_28_11_io_ins_2),
    .io_ins_3(ces_28_11_io_ins_3),
    .io_outs_0(ces_28_11_io_outs_0),
    .io_outs_1(ces_28_11_io_outs_1),
    .io_outs_2(ces_28_11_io_outs_2),
    .io_outs_3(ces_28_11_io_outs_3)
  );
  Element ces_28_12 ( // @[MockArray.scala 36:52]
    .clock(ces_28_12_clock),
    .io_ins_0(ces_28_12_io_ins_0),
    .io_ins_1(ces_28_12_io_ins_1),
    .io_ins_2(ces_28_12_io_ins_2),
    .io_ins_3(ces_28_12_io_ins_3),
    .io_outs_0(ces_28_12_io_outs_0),
    .io_outs_1(ces_28_12_io_outs_1),
    .io_outs_2(ces_28_12_io_outs_2),
    .io_outs_3(ces_28_12_io_outs_3)
  );
  Element ces_28_13 ( // @[MockArray.scala 36:52]
    .clock(ces_28_13_clock),
    .io_ins_0(ces_28_13_io_ins_0),
    .io_ins_1(ces_28_13_io_ins_1),
    .io_ins_2(ces_28_13_io_ins_2),
    .io_ins_3(ces_28_13_io_ins_3),
    .io_outs_0(ces_28_13_io_outs_0),
    .io_outs_1(ces_28_13_io_outs_1),
    .io_outs_2(ces_28_13_io_outs_2),
    .io_outs_3(ces_28_13_io_outs_3)
  );
  Element ces_28_14 ( // @[MockArray.scala 36:52]
    .clock(ces_28_14_clock),
    .io_ins_0(ces_28_14_io_ins_0),
    .io_ins_1(ces_28_14_io_ins_1),
    .io_ins_2(ces_28_14_io_ins_2),
    .io_ins_3(ces_28_14_io_ins_3),
    .io_outs_0(ces_28_14_io_outs_0),
    .io_outs_1(ces_28_14_io_outs_1),
    .io_outs_2(ces_28_14_io_outs_2),
    .io_outs_3(ces_28_14_io_outs_3)
  );
  Element ces_28_15 ( // @[MockArray.scala 36:52]
    .clock(ces_28_15_clock),
    .io_ins_0(ces_28_15_io_ins_0),
    .io_ins_1(ces_28_15_io_ins_1),
    .io_ins_2(ces_28_15_io_ins_2),
    .io_ins_3(ces_28_15_io_ins_3),
    .io_outs_0(ces_28_15_io_outs_0),
    .io_outs_1(ces_28_15_io_outs_1),
    .io_outs_2(ces_28_15_io_outs_2),
    .io_outs_3(ces_28_15_io_outs_3)
  );
  Element ces_28_16 ( // @[MockArray.scala 36:52]
    .clock(ces_28_16_clock),
    .io_ins_0(ces_28_16_io_ins_0),
    .io_ins_1(ces_28_16_io_ins_1),
    .io_ins_2(ces_28_16_io_ins_2),
    .io_ins_3(ces_28_16_io_ins_3),
    .io_outs_0(ces_28_16_io_outs_0),
    .io_outs_1(ces_28_16_io_outs_1),
    .io_outs_2(ces_28_16_io_outs_2),
    .io_outs_3(ces_28_16_io_outs_3)
  );
  Element ces_28_17 ( // @[MockArray.scala 36:52]
    .clock(ces_28_17_clock),
    .io_ins_0(ces_28_17_io_ins_0),
    .io_ins_1(ces_28_17_io_ins_1),
    .io_ins_2(ces_28_17_io_ins_2),
    .io_ins_3(ces_28_17_io_ins_3),
    .io_outs_0(ces_28_17_io_outs_0),
    .io_outs_1(ces_28_17_io_outs_1),
    .io_outs_2(ces_28_17_io_outs_2),
    .io_outs_3(ces_28_17_io_outs_3)
  );
  Element ces_28_18 ( // @[MockArray.scala 36:52]
    .clock(ces_28_18_clock),
    .io_ins_0(ces_28_18_io_ins_0),
    .io_ins_1(ces_28_18_io_ins_1),
    .io_ins_2(ces_28_18_io_ins_2),
    .io_ins_3(ces_28_18_io_ins_3),
    .io_outs_0(ces_28_18_io_outs_0),
    .io_outs_1(ces_28_18_io_outs_1),
    .io_outs_2(ces_28_18_io_outs_2),
    .io_outs_3(ces_28_18_io_outs_3)
  );
  Element ces_28_19 ( // @[MockArray.scala 36:52]
    .clock(ces_28_19_clock),
    .io_ins_0(ces_28_19_io_ins_0),
    .io_ins_1(ces_28_19_io_ins_1),
    .io_ins_2(ces_28_19_io_ins_2),
    .io_ins_3(ces_28_19_io_ins_3),
    .io_outs_0(ces_28_19_io_outs_0),
    .io_outs_1(ces_28_19_io_outs_1),
    .io_outs_2(ces_28_19_io_outs_2),
    .io_outs_3(ces_28_19_io_outs_3)
  );
  Element ces_28_20 ( // @[MockArray.scala 36:52]
    .clock(ces_28_20_clock),
    .io_ins_0(ces_28_20_io_ins_0),
    .io_ins_1(ces_28_20_io_ins_1),
    .io_ins_2(ces_28_20_io_ins_2),
    .io_ins_3(ces_28_20_io_ins_3),
    .io_outs_0(ces_28_20_io_outs_0),
    .io_outs_1(ces_28_20_io_outs_1),
    .io_outs_2(ces_28_20_io_outs_2),
    .io_outs_3(ces_28_20_io_outs_3)
  );
  Element ces_28_21 ( // @[MockArray.scala 36:52]
    .clock(ces_28_21_clock),
    .io_ins_0(ces_28_21_io_ins_0),
    .io_ins_1(ces_28_21_io_ins_1),
    .io_ins_2(ces_28_21_io_ins_2),
    .io_ins_3(ces_28_21_io_ins_3),
    .io_outs_0(ces_28_21_io_outs_0),
    .io_outs_1(ces_28_21_io_outs_1),
    .io_outs_2(ces_28_21_io_outs_2),
    .io_outs_3(ces_28_21_io_outs_3)
  );
  Element ces_28_22 ( // @[MockArray.scala 36:52]
    .clock(ces_28_22_clock),
    .io_ins_0(ces_28_22_io_ins_0),
    .io_ins_1(ces_28_22_io_ins_1),
    .io_ins_2(ces_28_22_io_ins_2),
    .io_ins_3(ces_28_22_io_ins_3),
    .io_outs_0(ces_28_22_io_outs_0),
    .io_outs_1(ces_28_22_io_outs_1),
    .io_outs_2(ces_28_22_io_outs_2),
    .io_outs_3(ces_28_22_io_outs_3)
  );
  Element ces_28_23 ( // @[MockArray.scala 36:52]
    .clock(ces_28_23_clock),
    .io_ins_0(ces_28_23_io_ins_0),
    .io_ins_1(ces_28_23_io_ins_1),
    .io_ins_2(ces_28_23_io_ins_2),
    .io_ins_3(ces_28_23_io_ins_3),
    .io_outs_0(ces_28_23_io_outs_0),
    .io_outs_1(ces_28_23_io_outs_1),
    .io_outs_2(ces_28_23_io_outs_2),
    .io_outs_3(ces_28_23_io_outs_3)
  );
  Element ces_28_24 ( // @[MockArray.scala 36:52]
    .clock(ces_28_24_clock),
    .io_ins_0(ces_28_24_io_ins_0),
    .io_ins_1(ces_28_24_io_ins_1),
    .io_ins_2(ces_28_24_io_ins_2),
    .io_ins_3(ces_28_24_io_ins_3),
    .io_outs_0(ces_28_24_io_outs_0),
    .io_outs_1(ces_28_24_io_outs_1),
    .io_outs_2(ces_28_24_io_outs_2),
    .io_outs_3(ces_28_24_io_outs_3)
  );
  Element ces_28_25 ( // @[MockArray.scala 36:52]
    .clock(ces_28_25_clock),
    .io_ins_0(ces_28_25_io_ins_0),
    .io_ins_1(ces_28_25_io_ins_1),
    .io_ins_2(ces_28_25_io_ins_2),
    .io_ins_3(ces_28_25_io_ins_3),
    .io_outs_0(ces_28_25_io_outs_0),
    .io_outs_1(ces_28_25_io_outs_1),
    .io_outs_2(ces_28_25_io_outs_2),
    .io_outs_3(ces_28_25_io_outs_3)
  );
  Element ces_28_26 ( // @[MockArray.scala 36:52]
    .clock(ces_28_26_clock),
    .io_ins_0(ces_28_26_io_ins_0),
    .io_ins_1(ces_28_26_io_ins_1),
    .io_ins_2(ces_28_26_io_ins_2),
    .io_ins_3(ces_28_26_io_ins_3),
    .io_outs_0(ces_28_26_io_outs_0),
    .io_outs_1(ces_28_26_io_outs_1),
    .io_outs_2(ces_28_26_io_outs_2),
    .io_outs_3(ces_28_26_io_outs_3)
  );
  Element ces_28_27 ( // @[MockArray.scala 36:52]
    .clock(ces_28_27_clock),
    .io_ins_0(ces_28_27_io_ins_0),
    .io_ins_1(ces_28_27_io_ins_1),
    .io_ins_2(ces_28_27_io_ins_2),
    .io_ins_3(ces_28_27_io_ins_3),
    .io_outs_0(ces_28_27_io_outs_0),
    .io_outs_1(ces_28_27_io_outs_1),
    .io_outs_2(ces_28_27_io_outs_2),
    .io_outs_3(ces_28_27_io_outs_3)
  );
  Element ces_28_28 ( // @[MockArray.scala 36:52]
    .clock(ces_28_28_clock),
    .io_ins_0(ces_28_28_io_ins_0),
    .io_ins_1(ces_28_28_io_ins_1),
    .io_ins_2(ces_28_28_io_ins_2),
    .io_ins_3(ces_28_28_io_ins_3),
    .io_outs_0(ces_28_28_io_outs_0),
    .io_outs_1(ces_28_28_io_outs_1),
    .io_outs_2(ces_28_28_io_outs_2),
    .io_outs_3(ces_28_28_io_outs_3)
  );
  Element ces_28_29 ( // @[MockArray.scala 36:52]
    .clock(ces_28_29_clock),
    .io_ins_0(ces_28_29_io_ins_0),
    .io_ins_1(ces_28_29_io_ins_1),
    .io_ins_2(ces_28_29_io_ins_2),
    .io_ins_3(ces_28_29_io_ins_3),
    .io_outs_0(ces_28_29_io_outs_0),
    .io_outs_1(ces_28_29_io_outs_1),
    .io_outs_2(ces_28_29_io_outs_2),
    .io_outs_3(ces_28_29_io_outs_3)
  );
  Element ces_28_30 ( // @[MockArray.scala 36:52]
    .clock(ces_28_30_clock),
    .io_ins_0(ces_28_30_io_ins_0),
    .io_ins_1(ces_28_30_io_ins_1),
    .io_ins_2(ces_28_30_io_ins_2),
    .io_ins_3(ces_28_30_io_ins_3),
    .io_outs_0(ces_28_30_io_outs_0),
    .io_outs_1(ces_28_30_io_outs_1),
    .io_outs_2(ces_28_30_io_outs_2),
    .io_outs_3(ces_28_30_io_outs_3)
  );
  Element ces_28_31 ( // @[MockArray.scala 36:52]
    .clock(ces_28_31_clock),
    .io_ins_0(ces_28_31_io_ins_0),
    .io_ins_1(ces_28_31_io_ins_1),
    .io_ins_2(ces_28_31_io_ins_2),
    .io_ins_3(ces_28_31_io_ins_3),
    .io_outs_0(ces_28_31_io_outs_0),
    .io_outs_1(ces_28_31_io_outs_1),
    .io_outs_2(ces_28_31_io_outs_2),
    .io_outs_3(ces_28_31_io_outs_3)
  );
  Element ces_29_0 ( // @[MockArray.scala 36:52]
    .clock(ces_29_0_clock),
    .io_ins_0(ces_29_0_io_ins_0),
    .io_ins_1(ces_29_0_io_ins_1),
    .io_ins_2(ces_29_0_io_ins_2),
    .io_ins_3(ces_29_0_io_ins_3),
    .io_outs_0(ces_29_0_io_outs_0),
    .io_outs_1(ces_29_0_io_outs_1),
    .io_outs_2(ces_29_0_io_outs_2),
    .io_outs_3(ces_29_0_io_outs_3)
  );
  Element ces_29_1 ( // @[MockArray.scala 36:52]
    .clock(ces_29_1_clock),
    .io_ins_0(ces_29_1_io_ins_0),
    .io_ins_1(ces_29_1_io_ins_1),
    .io_ins_2(ces_29_1_io_ins_2),
    .io_ins_3(ces_29_1_io_ins_3),
    .io_outs_0(ces_29_1_io_outs_0),
    .io_outs_1(ces_29_1_io_outs_1),
    .io_outs_2(ces_29_1_io_outs_2),
    .io_outs_3(ces_29_1_io_outs_3)
  );
  Element ces_29_2 ( // @[MockArray.scala 36:52]
    .clock(ces_29_2_clock),
    .io_ins_0(ces_29_2_io_ins_0),
    .io_ins_1(ces_29_2_io_ins_1),
    .io_ins_2(ces_29_2_io_ins_2),
    .io_ins_3(ces_29_2_io_ins_3),
    .io_outs_0(ces_29_2_io_outs_0),
    .io_outs_1(ces_29_2_io_outs_1),
    .io_outs_2(ces_29_2_io_outs_2),
    .io_outs_3(ces_29_2_io_outs_3)
  );
  Element ces_29_3 ( // @[MockArray.scala 36:52]
    .clock(ces_29_3_clock),
    .io_ins_0(ces_29_3_io_ins_0),
    .io_ins_1(ces_29_3_io_ins_1),
    .io_ins_2(ces_29_3_io_ins_2),
    .io_ins_3(ces_29_3_io_ins_3),
    .io_outs_0(ces_29_3_io_outs_0),
    .io_outs_1(ces_29_3_io_outs_1),
    .io_outs_2(ces_29_3_io_outs_2),
    .io_outs_3(ces_29_3_io_outs_3)
  );
  Element ces_29_4 ( // @[MockArray.scala 36:52]
    .clock(ces_29_4_clock),
    .io_ins_0(ces_29_4_io_ins_0),
    .io_ins_1(ces_29_4_io_ins_1),
    .io_ins_2(ces_29_4_io_ins_2),
    .io_ins_3(ces_29_4_io_ins_3),
    .io_outs_0(ces_29_4_io_outs_0),
    .io_outs_1(ces_29_4_io_outs_1),
    .io_outs_2(ces_29_4_io_outs_2),
    .io_outs_3(ces_29_4_io_outs_3)
  );
  Element ces_29_5 ( // @[MockArray.scala 36:52]
    .clock(ces_29_5_clock),
    .io_ins_0(ces_29_5_io_ins_0),
    .io_ins_1(ces_29_5_io_ins_1),
    .io_ins_2(ces_29_5_io_ins_2),
    .io_ins_3(ces_29_5_io_ins_3),
    .io_outs_0(ces_29_5_io_outs_0),
    .io_outs_1(ces_29_5_io_outs_1),
    .io_outs_2(ces_29_5_io_outs_2),
    .io_outs_3(ces_29_5_io_outs_3)
  );
  Element ces_29_6 ( // @[MockArray.scala 36:52]
    .clock(ces_29_6_clock),
    .io_ins_0(ces_29_6_io_ins_0),
    .io_ins_1(ces_29_6_io_ins_1),
    .io_ins_2(ces_29_6_io_ins_2),
    .io_ins_3(ces_29_6_io_ins_3),
    .io_outs_0(ces_29_6_io_outs_0),
    .io_outs_1(ces_29_6_io_outs_1),
    .io_outs_2(ces_29_6_io_outs_2),
    .io_outs_3(ces_29_6_io_outs_3)
  );
  Element ces_29_7 ( // @[MockArray.scala 36:52]
    .clock(ces_29_7_clock),
    .io_ins_0(ces_29_7_io_ins_0),
    .io_ins_1(ces_29_7_io_ins_1),
    .io_ins_2(ces_29_7_io_ins_2),
    .io_ins_3(ces_29_7_io_ins_3),
    .io_outs_0(ces_29_7_io_outs_0),
    .io_outs_1(ces_29_7_io_outs_1),
    .io_outs_2(ces_29_7_io_outs_2),
    .io_outs_3(ces_29_7_io_outs_3)
  );
  Element ces_29_8 ( // @[MockArray.scala 36:52]
    .clock(ces_29_8_clock),
    .io_ins_0(ces_29_8_io_ins_0),
    .io_ins_1(ces_29_8_io_ins_1),
    .io_ins_2(ces_29_8_io_ins_2),
    .io_ins_3(ces_29_8_io_ins_3),
    .io_outs_0(ces_29_8_io_outs_0),
    .io_outs_1(ces_29_8_io_outs_1),
    .io_outs_2(ces_29_8_io_outs_2),
    .io_outs_3(ces_29_8_io_outs_3)
  );
  Element ces_29_9 ( // @[MockArray.scala 36:52]
    .clock(ces_29_9_clock),
    .io_ins_0(ces_29_9_io_ins_0),
    .io_ins_1(ces_29_9_io_ins_1),
    .io_ins_2(ces_29_9_io_ins_2),
    .io_ins_3(ces_29_9_io_ins_3),
    .io_outs_0(ces_29_9_io_outs_0),
    .io_outs_1(ces_29_9_io_outs_1),
    .io_outs_2(ces_29_9_io_outs_2),
    .io_outs_3(ces_29_9_io_outs_3)
  );
  Element ces_29_10 ( // @[MockArray.scala 36:52]
    .clock(ces_29_10_clock),
    .io_ins_0(ces_29_10_io_ins_0),
    .io_ins_1(ces_29_10_io_ins_1),
    .io_ins_2(ces_29_10_io_ins_2),
    .io_ins_3(ces_29_10_io_ins_3),
    .io_outs_0(ces_29_10_io_outs_0),
    .io_outs_1(ces_29_10_io_outs_1),
    .io_outs_2(ces_29_10_io_outs_2),
    .io_outs_3(ces_29_10_io_outs_3)
  );
  Element ces_29_11 ( // @[MockArray.scala 36:52]
    .clock(ces_29_11_clock),
    .io_ins_0(ces_29_11_io_ins_0),
    .io_ins_1(ces_29_11_io_ins_1),
    .io_ins_2(ces_29_11_io_ins_2),
    .io_ins_3(ces_29_11_io_ins_3),
    .io_outs_0(ces_29_11_io_outs_0),
    .io_outs_1(ces_29_11_io_outs_1),
    .io_outs_2(ces_29_11_io_outs_2),
    .io_outs_3(ces_29_11_io_outs_3)
  );
  Element ces_29_12 ( // @[MockArray.scala 36:52]
    .clock(ces_29_12_clock),
    .io_ins_0(ces_29_12_io_ins_0),
    .io_ins_1(ces_29_12_io_ins_1),
    .io_ins_2(ces_29_12_io_ins_2),
    .io_ins_3(ces_29_12_io_ins_3),
    .io_outs_0(ces_29_12_io_outs_0),
    .io_outs_1(ces_29_12_io_outs_1),
    .io_outs_2(ces_29_12_io_outs_2),
    .io_outs_3(ces_29_12_io_outs_3)
  );
  Element ces_29_13 ( // @[MockArray.scala 36:52]
    .clock(ces_29_13_clock),
    .io_ins_0(ces_29_13_io_ins_0),
    .io_ins_1(ces_29_13_io_ins_1),
    .io_ins_2(ces_29_13_io_ins_2),
    .io_ins_3(ces_29_13_io_ins_3),
    .io_outs_0(ces_29_13_io_outs_0),
    .io_outs_1(ces_29_13_io_outs_1),
    .io_outs_2(ces_29_13_io_outs_2),
    .io_outs_3(ces_29_13_io_outs_3)
  );
  Element ces_29_14 ( // @[MockArray.scala 36:52]
    .clock(ces_29_14_clock),
    .io_ins_0(ces_29_14_io_ins_0),
    .io_ins_1(ces_29_14_io_ins_1),
    .io_ins_2(ces_29_14_io_ins_2),
    .io_ins_3(ces_29_14_io_ins_3),
    .io_outs_0(ces_29_14_io_outs_0),
    .io_outs_1(ces_29_14_io_outs_1),
    .io_outs_2(ces_29_14_io_outs_2),
    .io_outs_3(ces_29_14_io_outs_3)
  );
  Element ces_29_15 ( // @[MockArray.scala 36:52]
    .clock(ces_29_15_clock),
    .io_ins_0(ces_29_15_io_ins_0),
    .io_ins_1(ces_29_15_io_ins_1),
    .io_ins_2(ces_29_15_io_ins_2),
    .io_ins_3(ces_29_15_io_ins_3),
    .io_outs_0(ces_29_15_io_outs_0),
    .io_outs_1(ces_29_15_io_outs_1),
    .io_outs_2(ces_29_15_io_outs_2),
    .io_outs_3(ces_29_15_io_outs_3)
  );
  Element ces_29_16 ( // @[MockArray.scala 36:52]
    .clock(ces_29_16_clock),
    .io_ins_0(ces_29_16_io_ins_0),
    .io_ins_1(ces_29_16_io_ins_1),
    .io_ins_2(ces_29_16_io_ins_2),
    .io_ins_3(ces_29_16_io_ins_3),
    .io_outs_0(ces_29_16_io_outs_0),
    .io_outs_1(ces_29_16_io_outs_1),
    .io_outs_2(ces_29_16_io_outs_2),
    .io_outs_3(ces_29_16_io_outs_3)
  );
  Element ces_29_17 ( // @[MockArray.scala 36:52]
    .clock(ces_29_17_clock),
    .io_ins_0(ces_29_17_io_ins_0),
    .io_ins_1(ces_29_17_io_ins_1),
    .io_ins_2(ces_29_17_io_ins_2),
    .io_ins_3(ces_29_17_io_ins_3),
    .io_outs_0(ces_29_17_io_outs_0),
    .io_outs_1(ces_29_17_io_outs_1),
    .io_outs_2(ces_29_17_io_outs_2),
    .io_outs_3(ces_29_17_io_outs_3)
  );
  Element ces_29_18 ( // @[MockArray.scala 36:52]
    .clock(ces_29_18_clock),
    .io_ins_0(ces_29_18_io_ins_0),
    .io_ins_1(ces_29_18_io_ins_1),
    .io_ins_2(ces_29_18_io_ins_2),
    .io_ins_3(ces_29_18_io_ins_3),
    .io_outs_0(ces_29_18_io_outs_0),
    .io_outs_1(ces_29_18_io_outs_1),
    .io_outs_2(ces_29_18_io_outs_2),
    .io_outs_3(ces_29_18_io_outs_3)
  );
  Element ces_29_19 ( // @[MockArray.scala 36:52]
    .clock(ces_29_19_clock),
    .io_ins_0(ces_29_19_io_ins_0),
    .io_ins_1(ces_29_19_io_ins_1),
    .io_ins_2(ces_29_19_io_ins_2),
    .io_ins_3(ces_29_19_io_ins_3),
    .io_outs_0(ces_29_19_io_outs_0),
    .io_outs_1(ces_29_19_io_outs_1),
    .io_outs_2(ces_29_19_io_outs_2),
    .io_outs_3(ces_29_19_io_outs_3)
  );
  Element ces_29_20 ( // @[MockArray.scala 36:52]
    .clock(ces_29_20_clock),
    .io_ins_0(ces_29_20_io_ins_0),
    .io_ins_1(ces_29_20_io_ins_1),
    .io_ins_2(ces_29_20_io_ins_2),
    .io_ins_3(ces_29_20_io_ins_3),
    .io_outs_0(ces_29_20_io_outs_0),
    .io_outs_1(ces_29_20_io_outs_1),
    .io_outs_2(ces_29_20_io_outs_2),
    .io_outs_3(ces_29_20_io_outs_3)
  );
  Element ces_29_21 ( // @[MockArray.scala 36:52]
    .clock(ces_29_21_clock),
    .io_ins_0(ces_29_21_io_ins_0),
    .io_ins_1(ces_29_21_io_ins_1),
    .io_ins_2(ces_29_21_io_ins_2),
    .io_ins_3(ces_29_21_io_ins_3),
    .io_outs_0(ces_29_21_io_outs_0),
    .io_outs_1(ces_29_21_io_outs_1),
    .io_outs_2(ces_29_21_io_outs_2),
    .io_outs_3(ces_29_21_io_outs_3)
  );
  Element ces_29_22 ( // @[MockArray.scala 36:52]
    .clock(ces_29_22_clock),
    .io_ins_0(ces_29_22_io_ins_0),
    .io_ins_1(ces_29_22_io_ins_1),
    .io_ins_2(ces_29_22_io_ins_2),
    .io_ins_3(ces_29_22_io_ins_3),
    .io_outs_0(ces_29_22_io_outs_0),
    .io_outs_1(ces_29_22_io_outs_1),
    .io_outs_2(ces_29_22_io_outs_2),
    .io_outs_3(ces_29_22_io_outs_3)
  );
  Element ces_29_23 ( // @[MockArray.scala 36:52]
    .clock(ces_29_23_clock),
    .io_ins_0(ces_29_23_io_ins_0),
    .io_ins_1(ces_29_23_io_ins_1),
    .io_ins_2(ces_29_23_io_ins_2),
    .io_ins_3(ces_29_23_io_ins_3),
    .io_outs_0(ces_29_23_io_outs_0),
    .io_outs_1(ces_29_23_io_outs_1),
    .io_outs_2(ces_29_23_io_outs_2),
    .io_outs_3(ces_29_23_io_outs_3)
  );
  Element ces_29_24 ( // @[MockArray.scala 36:52]
    .clock(ces_29_24_clock),
    .io_ins_0(ces_29_24_io_ins_0),
    .io_ins_1(ces_29_24_io_ins_1),
    .io_ins_2(ces_29_24_io_ins_2),
    .io_ins_3(ces_29_24_io_ins_3),
    .io_outs_0(ces_29_24_io_outs_0),
    .io_outs_1(ces_29_24_io_outs_1),
    .io_outs_2(ces_29_24_io_outs_2),
    .io_outs_3(ces_29_24_io_outs_3)
  );
  Element ces_29_25 ( // @[MockArray.scala 36:52]
    .clock(ces_29_25_clock),
    .io_ins_0(ces_29_25_io_ins_0),
    .io_ins_1(ces_29_25_io_ins_1),
    .io_ins_2(ces_29_25_io_ins_2),
    .io_ins_3(ces_29_25_io_ins_3),
    .io_outs_0(ces_29_25_io_outs_0),
    .io_outs_1(ces_29_25_io_outs_1),
    .io_outs_2(ces_29_25_io_outs_2),
    .io_outs_3(ces_29_25_io_outs_3)
  );
  Element ces_29_26 ( // @[MockArray.scala 36:52]
    .clock(ces_29_26_clock),
    .io_ins_0(ces_29_26_io_ins_0),
    .io_ins_1(ces_29_26_io_ins_1),
    .io_ins_2(ces_29_26_io_ins_2),
    .io_ins_3(ces_29_26_io_ins_3),
    .io_outs_0(ces_29_26_io_outs_0),
    .io_outs_1(ces_29_26_io_outs_1),
    .io_outs_2(ces_29_26_io_outs_2),
    .io_outs_3(ces_29_26_io_outs_3)
  );
  Element ces_29_27 ( // @[MockArray.scala 36:52]
    .clock(ces_29_27_clock),
    .io_ins_0(ces_29_27_io_ins_0),
    .io_ins_1(ces_29_27_io_ins_1),
    .io_ins_2(ces_29_27_io_ins_2),
    .io_ins_3(ces_29_27_io_ins_3),
    .io_outs_0(ces_29_27_io_outs_0),
    .io_outs_1(ces_29_27_io_outs_1),
    .io_outs_2(ces_29_27_io_outs_2),
    .io_outs_3(ces_29_27_io_outs_3)
  );
  Element ces_29_28 ( // @[MockArray.scala 36:52]
    .clock(ces_29_28_clock),
    .io_ins_0(ces_29_28_io_ins_0),
    .io_ins_1(ces_29_28_io_ins_1),
    .io_ins_2(ces_29_28_io_ins_2),
    .io_ins_3(ces_29_28_io_ins_3),
    .io_outs_0(ces_29_28_io_outs_0),
    .io_outs_1(ces_29_28_io_outs_1),
    .io_outs_2(ces_29_28_io_outs_2),
    .io_outs_3(ces_29_28_io_outs_3)
  );
  Element ces_29_29 ( // @[MockArray.scala 36:52]
    .clock(ces_29_29_clock),
    .io_ins_0(ces_29_29_io_ins_0),
    .io_ins_1(ces_29_29_io_ins_1),
    .io_ins_2(ces_29_29_io_ins_2),
    .io_ins_3(ces_29_29_io_ins_3),
    .io_outs_0(ces_29_29_io_outs_0),
    .io_outs_1(ces_29_29_io_outs_1),
    .io_outs_2(ces_29_29_io_outs_2),
    .io_outs_3(ces_29_29_io_outs_3)
  );
  Element ces_29_30 ( // @[MockArray.scala 36:52]
    .clock(ces_29_30_clock),
    .io_ins_0(ces_29_30_io_ins_0),
    .io_ins_1(ces_29_30_io_ins_1),
    .io_ins_2(ces_29_30_io_ins_2),
    .io_ins_3(ces_29_30_io_ins_3),
    .io_outs_0(ces_29_30_io_outs_0),
    .io_outs_1(ces_29_30_io_outs_1),
    .io_outs_2(ces_29_30_io_outs_2),
    .io_outs_3(ces_29_30_io_outs_3)
  );
  Element ces_29_31 ( // @[MockArray.scala 36:52]
    .clock(ces_29_31_clock),
    .io_ins_0(ces_29_31_io_ins_0),
    .io_ins_1(ces_29_31_io_ins_1),
    .io_ins_2(ces_29_31_io_ins_2),
    .io_ins_3(ces_29_31_io_ins_3),
    .io_outs_0(ces_29_31_io_outs_0),
    .io_outs_1(ces_29_31_io_outs_1),
    .io_outs_2(ces_29_31_io_outs_2),
    .io_outs_3(ces_29_31_io_outs_3)
  );
  Element ces_30_0 ( // @[MockArray.scala 36:52]
    .clock(ces_30_0_clock),
    .io_ins_0(ces_30_0_io_ins_0),
    .io_ins_1(ces_30_0_io_ins_1),
    .io_ins_2(ces_30_0_io_ins_2),
    .io_ins_3(ces_30_0_io_ins_3),
    .io_outs_0(ces_30_0_io_outs_0),
    .io_outs_1(ces_30_0_io_outs_1),
    .io_outs_2(ces_30_0_io_outs_2),
    .io_outs_3(ces_30_0_io_outs_3)
  );
  Element ces_30_1 ( // @[MockArray.scala 36:52]
    .clock(ces_30_1_clock),
    .io_ins_0(ces_30_1_io_ins_0),
    .io_ins_1(ces_30_1_io_ins_1),
    .io_ins_2(ces_30_1_io_ins_2),
    .io_ins_3(ces_30_1_io_ins_3),
    .io_outs_0(ces_30_1_io_outs_0),
    .io_outs_1(ces_30_1_io_outs_1),
    .io_outs_2(ces_30_1_io_outs_2),
    .io_outs_3(ces_30_1_io_outs_3)
  );
  Element ces_30_2 ( // @[MockArray.scala 36:52]
    .clock(ces_30_2_clock),
    .io_ins_0(ces_30_2_io_ins_0),
    .io_ins_1(ces_30_2_io_ins_1),
    .io_ins_2(ces_30_2_io_ins_2),
    .io_ins_3(ces_30_2_io_ins_3),
    .io_outs_0(ces_30_2_io_outs_0),
    .io_outs_1(ces_30_2_io_outs_1),
    .io_outs_2(ces_30_2_io_outs_2),
    .io_outs_3(ces_30_2_io_outs_3)
  );
  Element ces_30_3 ( // @[MockArray.scala 36:52]
    .clock(ces_30_3_clock),
    .io_ins_0(ces_30_3_io_ins_0),
    .io_ins_1(ces_30_3_io_ins_1),
    .io_ins_2(ces_30_3_io_ins_2),
    .io_ins_3(ces_30_3_io_ins_3),
    .io_outs_0(ces_30_3_io_outs_0),
    .io_outs_1(ces_30_3_io_outs_1),
    .io_outs_2(ces_30_3_io_outs_2),
    .io_outs_3(ces_30_3_io_outs_3)
  );
  Element ces_30_4 ( // @[MockArray.scala 36:52]
    .clock(ces_30_4_clock),
    .io_ins_0(ces_30_4_io_ins_0),
    .io_ins_1(ces_30_4_io_ins_1),
    .io_ins_2(ces_30_4_io_ins_2),
    .io_ins_3(ces_30_4_io_ins_3),
    .io_outs_0(ces_30_4_io_outs_0),
    .io_outs_1(ces_30_4_io_outs_1),
    .io_outs_2(ces_30_4_io_outs_2),
    .io_outs_3(ces_30_4_io_outs_3)
  );
  Element ces_30_5 ( // @[MockArray.scala 36:52]
    .clock(ces_30_5_clock),
    .io_ins_0(ces_30_5_io_ins_0),
    .io_ins_1(ces_30_5_io_ins_1),
    .io_ins_2(ces_30_5_io_ins_2),
    .io_ins_3(ces_30_5_io_ins_3),
    .io_outs_0(ces_30_5_io_outs_0),
    .io_outs_1(ces_30_5_io_outs_1),
    .io_outs_2(ces_30_5_io_outs_2),
    .io_outs_3(ces_30_5_io_outs_3)
  );
  Element ces_30_6 ( // @[MockArray.scala 36:52]
    .clock(ces_30_6_clock),
    .io_ins_0(ces_30_6_io_ins_0),
    .io_ins_1(ces_30_6_io_ins_1),
    .io_ins_2(ces_30_6_io_ins_2),
    .io_ins_3(ces_30_6_io_ins_3),
    .io_outs_0(ces_30_6_io_outs_0),
    .io_outs_1(ces_30_6_io_outs_1),
    .io_outs_2(ces_30_6_io_outs_2),
    .io_outs_3(ces_30_6_io_outs_3)
  );
  Element ces_30_7 ( // @[MockArray.scala 36:52]
    .clock(ces_30_7_clock),
    .io_ins_0(ces_30_7_io_ins_0),
    .io_ins_1(ces_30_7_io_ins_1),
    .io_ins_2(ces_30_7_io_ins_2),
    .io_ins_3(ces_30_7_io_ins_3),
    .io_outs_0(ces_30_7_io_outs_0),
    .io_outs_1(ces_30_7_io_outs_1),
    .io_outs_2(ces_30_7_io_outs_2),
    .io_outs_3(ces_30_7_io_outs_3)
  );
  Element ces_30_8 ( // @[MockArray.scala 36:52]
    .clock(ces_30_8_clock),
    .io_ins_0(ces_30_8_io_ins_0),
    .io_ins_1(ces_30_8_io_ins_1),
    .io_ins_2(ces_30_8_io_ins_2),
    .io_ins_3(ces_30_8_io_ins_3),
    .io_outs_0(ces_30_8_io_outs_0),
    .io_outs_1(ces_30_8_io_outs_1),
    .io_outs_2(ces_30_8_io_outs_2),
    .io_outs_3(ces_30_8_io_outs_3)
  );
  Element ces_30_9 ( // @[MockArray.scala 36:52]
    .clock(ces_30_9_clock),
    .io_ins_0(ces_30_9_io_ins_0),
    .io_ins_1(ces_30_9_io_ins_1),
    .io_ins_2(ces_30_9_io_ins_2),
    .io_ins_3(ces_30_9_io_ins_3),
    .io_outs_0(ces_30_9_io_outs_0),
    .io_outs_1(ces_30_9_io_outs_1),
    .io_outs_2(ces_30_9_io_outs_2),
    .io_outs_3(ces_30_9_io_outs_3)
  );
  Element ces_30_10 ( // @[MockArray.scala 36:52]
    .clock(ces_30_10_clock),
    .io_ins_0(ces_30_10_io_ins_0),
    .io_ins_1(ces_30_10_io_ins_1),
    .io_ins_2(ces_30_10_io_ins_2),
    .io_ins_3(ces_30_10_io_ins_3),
    .io_outs_0(ces_30_10_io_outs_0),
    .io_outs_1(ces_30_10_io_outs_1),
    .io_outs_2(ces_30_10_io_outs_2),
    .io_outs_3(ces_30_10_io_outs_3)
  );
  Element ces_30_11 ( // @[MockArray.scala 36:52]
    .clock(ces_30_11_clock),
    .io_ins_0(ces_30_11_io_ins_0),
    .io_ins_1(ces_30_11_io_ins_1),
    .io_ins_2(ces_30_11_io_ins_2),
    .io_ins_3(ces_30_11_io_ins_3),
    .io_outs_0(ces_30_11_io_outs_0),
    .io_outs_1(ces_30_11_io_outs_1),
    .io_outs_2(ces_30_11_io_outs_2),
    .io_outs_3(ces_30_11_io_outs_3)
  );
  Element ces_30_12 ( // @[MockArray.scala 36:52]
    .clock(ces_30_12_clock),
    .io_ins_0(ces_30_12_io_ins_0),
    .io_ins_1(ces_30_12_io_ins_1),
    .io_ins_2(ces_30_12_io_ins_2),
    .io_ins_3(ces_30_12_io_ins_3),
    .io_outs_0(ces_30_12_io_outs_0),
    .io_outs_1(ces_30_12_io_outs_1),
    .io_outs_2(ces_30_12_io_outs_2),
    .io_outs_3(ces_30_12_io_outs_3)
  );
  Element ces_30_13 ( // @[MockArray.scala 36:52]
    .clock(ces_30_13_clock),
    .io_ins_0(ces_30_13_io_ins_0),
    .io_ins_1(ces_30_13_io_ins_1),
    .io_ins_2(ces_30_13_io_ins_2),
    .io_ins_3(ces_30_13_io_ins_3),
    .io_outs_0(ces_30_13_io_outs_0),
    .io_outs_1(ces_30_13_io_outs_1),
    .io_outs_2(ces_30_13_io_outs_2),
    .io_outs_3(ces_30_13_io_outs_3)
  );
  Element ces_30_14 ( // @[MockArray.scala 36:52]
    .clock(ces_30_14_clock),
    .io_ins_0(ces_30_14_io_ins_0),
    .io_ins_1(ces_30_14_io_ins_1),
    .io_ins_2(ces_30_14_io_ins_2),
    .io_ins_3(ces_30_14_io_ins_3),
    .io_outs_0(ces_30_14_io_outs_0),
    .io_outs_1(ces_30_14_io_outs_1),
    .io_outs_2(ces_30_14_io_outs_2),
    .io_outs_3(ces_30_14_io_outs_3)
  );
  Element ces_30_15 ( // @[MockArray.scala 36:52]
    .clock(ces_30_15_clock),
    .io_ins_0(ces_30_15_io_ins_0),
    .io_ins_1(ces_30_15_io_ins_1),
    .io_ins_2(ces_30_15_io_ins_2),
    .io_ins_3(ces_30_15_io_ins_3),
    .io_outs_0(ces_30_15_io_outs_0),
    .io_outs_1(ces_30_15_io_outs_1),
    .io_outs_2(ces_30_15_io_outs_2),
    .io_outs_3(ces_30_15_io_outs_3)
  );
  Element ces_30_16 ( // @[MockArray.scala 36:52]
    .clock(ces_30_16_clock),
    .io_ins_0(ces_30_16_io_ins_0),
    .io_ins_1(ces_30_16_io_ins_1),
    .io_ins_2(ces_30_16_io_ins_2),
    .io_ins_3(ces_30_16_io_ins_3),
    .io_outs_0(ces_30_16_io_outs_0),
    .io_outs_1(ces_30_16_io_outs_1),
    .io_outs_2(ces_30_16_io_outs_2),
    .io_outs_3(ces_30_16_io_outs_3)
  );
  Element ces_30_17 ( // @[MockArray.scala 36:52]
    .clock(ces_30_17_clock),
    .io_ins_0(ces_30_17_io_ins_0),
    .io_ins_1(ces_30_17_io_ins_1),
    .io_ins_2(ces_30_17_io_ins_2),
    .io_ins_3(ces_30_17_io_ins_3),
    .io_outs_0(ces_30_17_io_outs_0),
    .io_outs_1(ces_30_17_io_outs_1),
    .io_outs_2(ces_30_17_io_outs_2),
    .io_outs_3(ces_30_17_io_outs_3)
  );
  Element ces_30_18 ( // @[MockArray.scala 36:52]
    .clock(ces_30_18_clock),
    .io_ins_0(ces_30_18_io_ins_0),
    .io_ins_1(ces_30_18_io_ins_1),
    .io_ins_2(ces_30_18_io_ins_2),
    .io_ins_3(ces_30_18_io_ins_3),
    .io_outs_0(ces_30_18_io_outs_0),
    .io_outs_1(ces_30_18_io_outs_1),
    .io_outs_2(ces_30_18_io_outs_2),
    .io_outs_3(ces_30_18_io_outs_3)
  );
  Element ces_30_19 ( // @[MockArray.scala 36:52]
    .clock(ces_30_19_clock),
    .io_ins_0(ces_30_19_io_ins_0),
    .io_ins_1(ces_30_19_io_ins_1),
    .io_ins_2(ces_30_19_io_ins_2),
    .io_ins_3(ces_30_19_io_ins_3),
    .io_outs_0(ces_30_19_io_outs_0),
    .io_outs_1(ces_30_19_io_outs_1),
    .io_outs_2(ces_30_19_io_outs_2),
    .io_outs_3(ces_30_19_io_outs_3)
  );
  Element ces_30_20 ( // @[MockArray.scala 36:52]
    .clock(ces_30_20_clock),
    .io_ins_0(ces_30_20_io_ins_0),
    .io_ins_1(ces_30_20_io_ins_1),
    .io_ins_2(ces_30_20_io_ins_2),
    .io_ins_3(ces_30_20_io_ins_3),
    .io_outs_0(ces_30_20_io_outs_0),
    .io_outs_1(ces_30_20_io_outs_1),
    .io_outs_2(ces_30_20_io_outs_2),
    .io_outs_3(ces_30_20_io_outs_3)
  );
  Element ces_30_21 ( // @[MockArray.scala 36:52]
    .clock(ces_30_21_clock),
    .io_ins_0(ces_30_21_io_ins_0),
    .io_ins_1(ces_30_21_io_ins_1),
    .io_ins_2(ces_30_21_io_ins_2),
    .io_ins_3(ces_30_21_io_ins_3),
    .io_outs_0(ces_30_21_io_outs_0),
    .io_outs_1(ces_30_21_io_outs_1),
    .io_outs_2(ces_30_21_io_outs_2),
    .io_outs_3(ces_30_21_io_outs_3)
  );
  Element ces_30_22 ( // @[MockArray.scala 36:52]
    .clock(ces_30_22_clock),
    .io_ins_0(ces_30_22_io_ins_0),
    .io_ins_1(ces_30_22_io_ins_1),
    .io_ins_2(ces_30_22_io_ins_2),
    .io_ins_3(ces_30_22_io_ins_3),
    .io_outs_0(ces_30_22_io_outs_0),
    .io_outs_1(ces_30_22_io_outs_1),
    .io_outs_2(ces_30_22_io_outs_2),
    .io_outs_3(ces_30_22_io_outs_3)
  );
  Element ces_30_23 ( // @[MockArray.scala 36:52]
    .clock(ces_30_23_clock),
    .io_ins_0(ces_30_23_io_ins_0),
    .io_ins_1(ces_30_23_io_ins_1),
    .io_ins_2(ces_30_23_io_ins_2),
    .io_ins_3(ces_30_23_io_ins_3),
    .io_outs_0(ces_30_23_io_outs_0),
    .io_outs_1(ces_30_23_io_outs_1),
    .io_outs_2(ces_30_23_io_outs_2),
    .io_outs_3(ces_30_23_io_outs_3)
  );
  Element ces_30_24 ( // @[MockArray.scala 36:52]
    .clock(ces_30_24_clock),
    .io_ins_0(ces_30_24_io_ins_0),
    .io_ins_1(ces_30_24_io_ins_1),
    .io_ins_2(ces_30_24_io_ins_2),
    .io_ins_3(ces_30_24_io_ins_3),
    .io_outs_0(ces_30_24_io_outs_0),
    .io_outs_1(ces_30_24_io_outs_1),
    .io_outs_2(ces_30_24_io_outs_2),
    .io_outs_3(ces_30_24_io_outs_3)
  );
  Element ces_30_25 ( // @[MockArray.scala 36:52]
    .clock(ces_30_25_clock),
    .io_ins_0(ces_30_25_io_ins_0),
    .io_ins_1(ces_30_25_io_ins_1),
    .io_ins_2(ces_30_25_io_ins_2),
    .io_ins_3(ces_30_25_io_ins_3),
    .io_outs_0(ces_30_25_io_outs_0),
    .io_outs_1(ces_30_25_io_outs_1),
    .io_outs_2(ces_30_25_io_outs_2),
    .io_outs_3(ces_30_25_io_outs_3)
  );
  Element ces_30_26 ( // @[MockArray.scala 36:52]
    .clock(ces_30_26_clock),
    .io_ins_0(ces_30_26_io_ins_0),
    .io_ins_1(ces_30_26_io_ins_1),
    .io_ins_2(ces_30_26_io_ins_2),
    .io_ins_3(ces_30_26_io_ins_3),
    .io_outs_0(ces_30_26_io_outs_0),
    .io_outs_1(ces_30_26_io_outs_1),
    .io_outs_2(ces_30_26_io_outs_2),
    .io_outs_3(ces_30_26_io_outs_3)
  );
  Element ces_30_27 ( // @[MockArray.scala 36:52]
    .clock(ces_30_27_clock),
    .io_ins_0(ces_30_27_io_ins_0),
    .io_ins_1(ces_30_27_io_ins_1),
    .io_ins_2(ces_30_27_io_ins_2),
    .io_ins_3(ces_30_27_io_ins_3),
    .io_outs_0(ces_30_27_io_outs_0),
    .io_outs_1(ces_30_27_io_outs_1),
    .io_outs_2(ces_30_27_io_outs_2),
    .io_outs_3(ces_30_27_io_outs_3)
  );
  Element ces_30_28 ( // @[MockArray.scala 36:52]
    .clock(ces_30_28_clock),
    .io_ins_0(ces_30_28_io_ins_0),
    .io_ins_1(ces_30_28_io_ins_1),
    .io_ins_2(ces_30_28_io_ins_2),
    .io_ins_3(ces_30_28_io_ins_3),
    .io_outs_0(ces_30_28_io_outs_0),
    .io_outs_1(ces_30_28_io_outs_1),
    .io_outs_2(ces_30_28_io_outs_2),
    .io_outs_3(ces_30_28_io_outs_3)
  );
  Element ces_30_29 ( // @[MockArray.scala 36:52]
    .clock(ces_30_29_clock),
    .io_ins_0(ces_30_29_io_ins_0),
    .io_ins_1(ces_30_29_io_ins_1),
    .io_ins_2(ces_30_29_io_ins_2),
    .io_ins_3(ces_30_29_io_ins_3),
    .io_outs_0(ces_30_29_io_outs_0),
    .io_outs_1(ces_30_29_io_outs_1),
    .io_outs_2(ces_30_29_io_outs_2),
    .io_outs_3(ces_30_29_io_outs_3)
  );
  Element ces_30_30 ( // @[MockArray.scala 36:52]
    .clock(ces_30_30_clock),
    .io_ins_0(ces_30_30_io_ins_0),
    .io_ins_1(ces_30_30_io_ins_1),
    .io_ins_2(ces_30_30_io_ins_2),
    .io_ins_3(ces_30_30_io_ins_3),
    .io_outs_0(ces_30_30_io_outs_0),
    .io_outs_1(ces_30_30_io_outs_1),
    .io_outs_2(ces_30_30_io_outs_2),
    .io_outs_3(ces_30_30_io_outs_3)
  );
  Element ces_30_31 ( // @[MockArray.scala 36:52]
    .clock(ces_30_31_clock),
    .io_ins_0(ces_30_31_io_ins_0),
    .io_ins_1(ces_30_31_io_ins_1),
    .io_ins_2(ces_30_31_io_ins_2),
    .io_ins_3(ces_30_31_io_ins_3),
    .io_outs_0(ces_30_31_io_outs_0),
    .io_outs_1(ces_30_31_io_outs_1),
    .io_outs_2(ces_30_31_io_outs_2),
    .io_outs_3(ces_30_31_io_outs_3)
  );
  Element ces_31_0 ( // @[MockArray.scala 36:52]
    .clock(ces_31_0_clock),
    .io_ins_0(ces_31_0_io_ins_0),
    .io_ins_1(ces_31_0_io_ins_1),
    .io_ins_2(ces_31_0_io_ins_2),
    .io_ins_3(ces_31_0_io_ins_3),
    .io_outs_0(ces_31_0_io_outs_0),
    .io_outs_1(ces_31_0_io_outs_1),
    .io_outs_2(ces_31_0_io_outs_2),
    .io_outs_3(ces_31_0_io_outs_3)
  );
  Element ces_31_1 ( // @[MockArray.scala 36:52]
    .clock(ces_31_1_clock),
    .io_ins_0(ces_31_1_io_ins_0),
    .io_ins_1(ces_31_1_io_ins_1),
    .io_ins_2(ces_31_1_io_ins_2),
    .io_ins_3(ces_31_1_io_ins_3),
    .io_outs_0(ces_31_1_io_outs_0),
    .io_outs_1(ces_31_1_io_outs_1),
    .io_outs_2(ces_31_1_io_outs_2),
    .io_outs_3(ces_31_1_io_outs_3)
  );
  Element ces_31_2 ( // @[MockArray.scala 36:52]
    .clock(ces_31_2_clock),
    .io_ins_0(ces_31_2_io_ins_0),
    .io_ins_1(ces_31_2_io_ins_1),
    .io_ins_2(ces_31_2_io_ins_2),
    .io_ins_3(ces_31_2_io_ins_3),
    .io_outs_0(ces_31_2_io_outs_0),
    .io_outs_1(ces_31_2_io_outs_1),
    .io_outs_2(ces_31_2_io_outs_2),
    .io_outs_3(ces_31_2_io_outs_3)
  );
  Element ces_31_3 ( // @[MockArray.scala 36:52]
    .clock(ces_31_3_clock),
    .io_ins_0(ces_31_3_io_ins_0),
    .io_ins_1(ces_31_3_io_ins_1),
    .io_ins_2(ces_31_3_io_ins_2),
    .io_ins_3(ces_31_3_io_ins_3),
    .io_outs_0(ces_31_3_io_outs_0),
    .io_outs_1(ces_31_3_io_outs_1),
    .io_outs_2(ces_31_3_io_outs_2),
    .io_outs_3(ces_31_3_io_outs_3)
  );
  Element ces_31_4 ( // @[MockArray.scala 36:52]
    .clock(ces_31_4_clock),
    .io_ins_0(ces_31_4_io_ins_0),
    .io_ins_1(ces_31_4_io_ins_1),
    .io_ins_2(ces_31_4_io_ins_2),
    .io_ins_3(ces_31_4_io_ins_3),
    .io_outs_0(ces_31_4_io_outs_0),
    .io_outs_1(ces_31_4_io_outs_1),
    .io_outs_2(ces_31_4_io_outs_2),
    .io_outs_3(ces_31_4_io_outs_3)
  );
  Element ces_31_5 ( // @[MockArray.scala 36:52]
    .clock(ces_31_5_clock),
    .io_ins_0(ces_31_5_io_ins_0),
    .io_ins_1(ces_31_5_io_ins_1),
    .io_ins_2(ces_31_5_io_ins_2),
    .io_ins_3(ces_31_5_io_ins_3),
    .io_outs_0(ces_31_5_io_outs_0),
    .io_outs_1(ces_31_5_io_outs_1),
    .io_outs_2(ces_31_5_io_outs_2),
    .io_outs_3(ces_31_5_io_outs_3)
  );
  Element ces_31_6 ( // @[MockArray.scala 36:52]
    .clock(ces_31_6_clock),
    .io_ins_0(ces_31_6_io_ins_0),
    .io_ins_1(ces_31_6_io_ins_1),
    .io_ins_2(ces_31_6_io_ins_2),
    .io_ins_3(ces_31_6_io_ins_3),
    .io_outs_0(ces_31_6_io_outs_0),
    .io_outs_1(ces_31_6_io_outs_1),
    .io_outs_2(ces_31_6_io_outs_2),
    .io_outs_3(ces_31_6_io_outs_3)
  );
  Element ces_31_7 ( // @[MockArray.scala 36:52]
    .clock(ces_31_7_clock),
    .io_ins_0(ces_31_7_io_ins_0),
    .io_ins_1(ces_31_7_io_ins_1),
    .io_ins_2(ces_31_7_io_ins_2),
    .io_ins_3(ces_31_7_io_ins_3),
    .io_outs_0(ces_31_7_io_outs_0),
    .io_outs_1(ces_31_7_io_outs_1),
    .io_outs_2(ces_31_7_io_outs_2),
    .io_outs_3(ces_31_7_io_outs_3)
  );
  Element ces_31_8 ( // @[MockArray.scala 36:52]
    .clock(ces_31_8_clock),
    .io_ins_0(ces_31_8_io_ins_0),
    .io_ins_1(ces_31_8_io_ins_1),
    .io_ins_2(ces_31_8_io_ins_2),
    .io_ins_3(ces_31_8_io_ins_3),
    .io_outs_0(ces_31_8_io_outs_0),
    .io_outs_1(ces_31_8_io_outs_1),
    .io_outs_2(ces_31_8_io_outs_2),
    .io_outs_3(ces_31_8_io_outs_3)
  );
  Element ces_31_9 ( // @[MockArray.scala 36:52]
    .clock(ces_31_9_clock),
    .io_ins_0(ces_31_9_io_ins_0),
    .io_ins_1(ces_31_9_io_ins_1),
    .io_ins_2(ces_31_9_io_ins_2),
    .io_ins_3(ces_31_9_io_ins_3),
    .io_outs_0(ces_31_9_io_outs_0),
    .io_outs_1(ces_31_9_io_outs_1),
    .io_outs_2(ces_31_9_io_outs_2),
    .io_outs_3(ces_31_9_io_outs_3)
  );
  Element ces_31_10 ( // @[MockArray.scala 36:52]
    .clock(ces_31_10_clock),
    .io_ins_0(ces_31_10_io_ins_0),
    .io_ins_1(ces_31_10_io_ins_1),
    .io_ins_2(ces_31_10_io_ins_2),
    .io_ins_3(ces_31_10_io_ins_3),
    .io_outs_0(ces_31_10_io_outs_0),
    .io_outs_1(ces_31_10_io_outs_1),
    .io_outs_2(ces_31_10_io_outs_2),
    .io_outs_3(ces_31_10_io_outs_3)
  );
  Element ces_31_11 ( // @[MockArray.scala 36:52]
    .clock(ces_31_11_clock),
    .io_ins_0(ces_31_11_io_ins_0),
    .io_ins_1(ces_31_11_io_ins_1),
    .io_ins_2(ces_31_11_io_ins_2),
    .io_ins_3(ces_31_11_io_ins_3),
    .io_outs_0(ces_31_11_io_outs_0),
    .io_outs_1(ces_31_11_io_outs_1),
    .io_outs_2(ces_31_11_io_outs_2),
    .io_outs_3(ces_31_11_io_outs_3)
  );
  Element ces_31_12 ( // @[MockArray.scala 36:52]
    .clock(ces_31_12_clock),
    .io_ins_0(ces_31_12_io_ins_0),
    .io_ins_1(ces_31_12_io_ins_1),
    .io_ins_2(ces_31_12_io_ins_2),
    .io_ins_3(ces_31_12_io_ins_3),
    .io_outs_0(ces_31_12_io_outs_0),
    .io_outs_1(ces_31_12_io_outs_1),
    .io_outs_2(ces_31_12_io_outs_2),
    .io_outs_3(ces_31_12_io_outs_3)
  );
  Element ces_31_13 ( // @[MockArray.scala 36:52]
    .clock(ces_31_13_clock),
    .io_ins_0(ces_31_13_io_ins_0),
    .io_ins_1(ces_31_13_io_ins_1),
    .io_ins_2(ces_31_13_io_ins_2),
    .io_ins_3(ces_31_13_io_ins_3),
    .io_outs_0(ces_31_13_io_outs_0),
    .io_outs_1(ces_31_13_io_outs_1),
    .io_outs_2(ces_31_13_io_outs_2),
    .io_outs_3(ces_31_13_io_outs_3)
  );
  Element ces_31_14 ( // @[MockArray.scala 36:52]
    .clock(ces_31_14_clock),
    .io_ins_0(ces_31_14_io_ins_0),
    .io_ins_1(ces_31_14_io_ins_1),
    .io_ins_2(ces_31_14_io_ins_2),
    .io_ins_3(ces_31_14_io_ins_3),
    .io_outs_0(ces_31_14_io_outs_0),
    .io_outs_1(ces_31_14_io_outs_1),
    .io_outs_2(ces_31_14_io_outs_2),
    .io_outs_3(ces_31_14_io_outs_3)
  );
  Element ces_31_15 ( // @[MockArray.scala 36:52]
    .clock(ces_31_15_clock),
    .io_ins_0(ces_31_15_io_ins_0),
    .io_ins_1(ces_31_15_io_ins_1),
    .io_ins_2(ces_31_15_io_ins_2),
    .io_ins_3(ces_31_15_io_ins_3),
    .io_outs_0(ces_31_15_io_outs_0),
    .io_outs_1(ces_31_15_io_outs_1),
    .io_outs_2(ces_31_15_io_outs_2),
    .io_outs_3(ces_31_15_io_outs_3)
  );
  Element ces_31_16 ( // @[MockArray.scala 36:52]
    .clock(ces_31_16_clock),
    .io_ins_0(ces_31_16_io_ins_0),
    .io_ins_1(ces_31_16_io_ins_1),
    .io_ins_2(ces_31_16_io_ins_2),
    .io_ins_3(ces_31_16_io_ins_3),
    .io_outs_0(ces_31_16_io_outs_0),
    .io_outs_1(ces_31_16_io_outs_1),
    .io_outs_2(ces_31_16_io_outs_2),
    .io_outs_3(ces_31_16_io_outs_3)
  );
  Element ces_31_17 ( // @[MockArray.scala 36:52]
    .clock(ces_31_17_clock),
    .io_ins_0(ces_31_17_io_ins_0),
    .io_ins_1(ces_31_17_io_ins_1),
    .io_ins_2(ces_31_17_io_ins_2),
    .io_ins_3(ces_31_17_io_ins_3),
    .io_outs_0(ces_31_17_io_outs_0),
    .io_outs_1(ces_31_17_io_outs_1),
    .io_outs_2(ces_31_17_io_outs_2),
    .io_outs_3(ces_31_17_io_outs_3)
  );
  Element ces_31_18 ( // @[MockArray.scala 36:52]
    .clock(ces_31_18_clock),
    .io_ins_0(ces_31_18_io_ins_0),
    .io_ins_1(ces_31_18_io_ins_1),
    .io_ins_2(ces_31_18_io_ins_2),
    .io_ins_3(ces_31_18_io_ins_3),
    .io_outs_0(ces_31_18_io_outs_0),
    .io_outs_1(ces_31_18_io_outs_1),
    .io_outs_2(ces_31_18_io_outs_2),
    .io_outs_3(ces_31_18_io_outs_3)
  );
  Element ces_31_19 ( // @[MockArray.scala 36:52]
    .clock(ces_31_19_clock),
    .io_ins_0(ces_31_19_io_ins_0),
    .io_ins_1(ces_31_19_io_ins_1),
    .io_ins_2(ces_31_19_io_ins_2),
    .io_ins_3(ces_31_19_io_ins_3),
    .io_outs_0(ces_31_19_io_outs_0),
    .io_outs_1(ces_31_19_io_outs_1),
    .io_outs_2(ces_31_19_io_outs_2),
    .io_outs_3(ces_31_19_io_outs_3)
  );
  Element ces_31_20 ( // @[MockArray.scala 36:52]
    .clock(ces_31_20_clock),
    .io_ins_0(ces_31_20_io_ins_0),
    .io_ins_1(ces_31_20_io_ins_1),
    .io_ins_2(ces_31_20_io_ins_2),
    .io_ins_3(ces_31_20_io_ins_3),
    .io_outs_0(ces_31_20_io_outs_0),
    .io_outs_1(ces_31_20_io_outs_1),
    .io_outs_2(ces_31_20_io_outs_2),
    .io_outs_3(ces_31_20_io_outs_3)
  );
  Element ces_31_21 ( // @[MockArray.scala 36:52]
    .clock(ces_31_21_clock),
    .io_ins_0(ces_31_21_io_ins_0),
    .io_ins_1(ces_31_21_io_ins_1),
    .io_ins_2(ces_31_21_io_ins_2),
    .io_ins_3(ces_31_21_io_ins_3),
    .io_outs_0(ces_31_21_io_outs_0),
    .io_outs_1(ces_31_21_io_outs_1),
    .io_outs_2(ces_31_21_io_outs_2),
    .io_outs_3(ces_31_21_io_outs_3)
  );
  Element ces_31_22 ( // @[MockArray.scala 36:52]
    .clock(ces_31_22_clock),
    .io_ins_0(ces_31_22_io_ins_0),
    .io_ins_1(ces_31_22_io_ins_1),
    .io_ins_2(ces_31_22_io_ins_2),
    .io_ins_3(ces_31_22_io_ins_3),
    .io_outs_0(ces_31_22_io_outs_0),
    .io_outs_1(ces_31_22_io_outs_1),
    .io_outs_2(ces_31_22_io_outs_2),
    .io_outs_3(ces_31_22_io_outs_3)
  );
  Element ces_31_23 ( // @[MockArray.scala 36:52]
    .clock(ces_31_23_clock),
    .io_ins_0(ces_31_23_io_ins_0),
    .io_ins_1(ces_31_23_io_ins_1),
    .io_ins_2(ces_31_23_io_ins_2),
    .io_ins_3(ces_31_23_io_ins_3),
    .io_outs_0(ces_31_23_io_outs_0),
    .io_outs_1(ces_31_23_io_outs_1),
    .io_outs_2(ces_31_23_io_outs_2),
    .io_outs_3(ces_31_23_io_outs_3)
  );
  Element ces_31_24 ( // @[MockArray.scala 36:52]
    .clock(ces_31_24_clock),
    .io_ins_0(ces_31_24_io_ins_0),
    .io_ins_1(ces_31_24_io_ins_1),
    .io_ins_2(ces_31_24_io_ins_2),
    .io_ins_3(ces_31_24_io_ins_3),
    .io_outs_0(ces_31_24_io_outs_0),
    .io_outs_1(ces_31_24_io_outs_1),
    .io_outs_2(ces_31_24_io_outs_2),
    .io_outs_3(ces_31_24_io_outs_3)
  );
  Element ces_31_25 ( // @[MockArray.scala 36:52]
    .clock(ces_31_25_clock),
    .io_ins_0(ces_31_25_io_ins_0),
    .io_ins_1(ces_31_25_io_ins_1),
    .io_ins_2(ces_31_25_io_ins_2),
    .io_ins_3(ces_31_25_io_ins_3),
    .io_outs_0(ces_31_25_io_outs_0),
    .io_outs_1(ces_31_25_io_outs_1),
    .io_outs_2(ces_31_25_io_outs_2),
    .io_outs_3(ces_31_25_io_outs_3)
  );
  Element ces_31_26 ( // @[MockArray.scala 36:52]
    .clock(ces_31_26_clock),
    .io_ins_0(ces_31_26_io_ins_0),
    .io_ins_1(ces_31_26_io_ins_1),
    .io_ins_2(ces_31_26_io_ins_2),
    .io_ins_3(ces_31_26_io_ins_3),
    .io_outs_0(ces_31_26_io_outs_0),
    .io_outs_1(ces_31_26_io_outs_1),
    .io_outs_2(ces_31_26_io_outs_2),
    .io_outs_3(ces_31_26_io_outs_3)
  );
  Element ces_31_27 ( // @[MockArray.scala 36:52]
    .clock(ces_31_27_clock),
    .io_ins_0(ces_31_27_io_ins_0),
    .io_ins_1(ces_31_27_io_ins_1),
    .io_ins_2(ces_31_27_io_ins_2),
    .io_ins_3(ces_31_27_io_ins_3),
    .io_outs_0(ces_31_27_io_outs_0),
    .io_outs_1(ces_31_27_io_outs_1),
    .io_outs_2(ces_31_27_io_outs_2),
    .io_outs_3(ces_31_27_io_outs_3)
  );
  Element ces_31_28 ( // @[MockArray.scala 36:52]
    .clock(ces_31_28_clock),
    .io_ins_0(ces_31_28_io_ins_0),
    .io_ins_1(ces_31_28_io_ins_1),
    .io_ins_2(ces_31_28_io_ins_2),
    .io_ins_3(ces_31_28_io_ins_3),
    .io_outs_0(ces_31_28_io_outs_0),
    .io_outs_1(ces_31_28_io_outs_1),
    .io_outs_2(ces_31_28_io_outs_2),
    .io_outs_3(ces_31_28_io_outs_3)
  );
  Element ces_31_29 ( // @[MockArray.scala 36:52]
    .clock(ces_31_29_clock),
    .io_ins_0(ces_31_29_io_ins_0),
    .io_ins_1(ces_31_29_io_ins_1),
    .io_ins_2(ces_31_29_io_ins_2),
    .io_ins_3(ces_31_29_io_ins_3),
    .io_outs_0(ces_31_29_io_outs_0),
    .io_outs_1(ces_31_29_io_outs_1),
    .io_outs_2(ces_31_29_io_outs_2),
    .io_outs_3(ces_31_29_io_outs_3)
  );
  Element ces_31_30 ( // @[MockArray.scala 36:52]
    .clock(ces_31_30_clock),
    .io_ins_0(ces_31_30_io_ins_0),
    .io_ins_1(ces_31_30_io_ins_1),
    .io_ins_2(ces_31_30_io_ins_2),
    .io_ins_3(ces_31_30_io_ins_3),
    .io_outs_0(ces_31_30_io_outs_0),
    .io_outs_1(ces_31_30_io_outs_1),
    .io_outs_2(ces_31_30_io_outs_2),
    .io_outs_3(ces_31_30_io_outs_3)
  );
  Element ces_31_31 ( // @[MockArray.scala 36:52]
    .clock(ces_31_31_clock),
    .io_ins_0(ces_31_31_io_ins_0),
    .io_ins_1(ces_31_31_io_ins_1),
    .io_ins_2(ces_31_31_io_ins_2),
    .io_ins_3(ces_31_31_io_ins_3),
    .io_outs_0(ces_31_31_io_outs_0),
    .io_outs_1(ces_31_31_io_outs_1),
    .io_outs_2(ces_31_31_io_outs_2),
    .io_outs_3(ces_31_31_io_outs_3)
  );
  assign io_outsHorizontal_0_0 = ces_0_0_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_1 = ces_0_1_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_2 = ces_0_2_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_3 = ces_0_3_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_4 = ces_0_4_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_5 = ces_0_5_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_6 = ces_0_6_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_7 = ces_0_7_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_8 = ces_0_8_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_9 = ces_0_9_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_10 = ces_0_10_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_11 = ces_0_11_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_12 = ces_0_12_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_13 = ces_0_13_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_14 = ces_0_14_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_15 = ces_0_15_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_16 = ces_0_16_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_17 = ces_0_17_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_18 = ces_0_18_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_19 = ces_0_19_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_20 = ces_0_20_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_21 = ces_0_21_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_22 = ces_0_22_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_23 = ces_0_23_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_24 = ces_0_24_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_25 = ces_0_25_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_26 = ces_0_26_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_27 = ces_0_27_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_28 = ces_0_28_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_29 = ces_0_29_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_30 = ces_0_30_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_0_31 = ces_0_31_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_1_0 = ces_31_0_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_1 = ces_31_1_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_2 = ces_31_2_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_3 = ces_31_3_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_4 = ces_31_4_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_5 = ces_31_5_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_6 = ces_31_6_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_7 = ces_31_7_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_8 = ces_31_8_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_9 = ces_31_9_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_10 = ces_31_10_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_11 = ces_31_11_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_12 = ces_31_12_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_13 = ces_31_13_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_14 = ces_31_14_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_15 = ces_31_15_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_16 = ces_31_16_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_17 = ces_31_17_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_18 = ces_31_18_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_19 = ces_31_19_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_20 = ces_31_20_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_21 = ces_31_21_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_22 = ces_31_22_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_23 = ces_31_23_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_24 = ces_31_24_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_25 = ces_31_25_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_26 = ces_31_26_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_27 = ces_31_27_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_28 = ces_31_28_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_29 = ces_31_29_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_30 = ces_31_30_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsHorizontal_1_31 = ces_31_31_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_0 = ces_0_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_1 = ces_1_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_2 = ces_2_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_3 = ces_3_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_4 = ces_4_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_5 = ces_5_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_6 = ces_6_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_7 = ces_7_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_8 = ces_8_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_9 = ces_9_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_10 = ces_10_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_11 = ces_11_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_12 = ces_12_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_13 = ces_13_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_14 = ces_14_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_15 = ces_15_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_16 = ces_16_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_17 = ces_17_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_18 = ces_18_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_19 = ces_19_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_20 = ces_20_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_21 = ces_21_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_22 = ces_22_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_23 = ces_23_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_24 = ces_24_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_25 = ces_25_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_26 = ces_26_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_27 = ces_27_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_28 = ces_28_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_29 = ces_29_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_30 = ces_30_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_31 = ces_31_31_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_1_0 = ces_0_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_1 = ces_1_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_2 = ces_2_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_3 = ces_3_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_4 = ces_4_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_5 = ces_5_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_6 = ces_6_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_7 = ces_7_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_8 = ces_8_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_9 = ces_9_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_10 = ces_10_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_11 = ces_11_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_12 = ces_12_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_13 = ces_13_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_14 = ces_14_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_15 = ces_15_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_16 = ces_16_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_17 = ces_17_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_18 = ces_18_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_19 = ces_19_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_20 = ces_20_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_21 = ces_21_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_22 = ces_22_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_23 = ces_23_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_24 = ces_24_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_25 = ces_25_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_26 = ces_26_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_27 = ces_27_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_28 = ces_28_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_29 = ces_29_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_30 = ces_30_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_31 = ces_31_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_lsbs_0 = ces_0_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1 = ces_0_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_2 = ces_0_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_3 = ces_0_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_4 = ces_0_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_5 = ces_0_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_6 = ces_0_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_7 = ces_0_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_8 = ces_0_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_9 = ces_0_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_10 = ces_0_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_11 = ces_0_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_12 = ces_0_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_13 = ces_0_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_14 = ces_0_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_15 = ces_0_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_16 = ces_0_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_17 = ces_0_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_18 = ces_0_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_19 = ces_0_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_20 = ces_0_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_21 = ces_0_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_22 = ces_0_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_23 = ces_0_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_24 = ces_0_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_25 = ces_0_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_26 = ces_0_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_27 = ces_0_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_28 = ces_0_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_29 = ces_0_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_30 = ces_0_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_31 = ces_0_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_32 = ces_1_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_33 = ces_1_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_34 = ces_1_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_35 = ces_1_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_36 = ces_1_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_37 = ces_1_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_38 = ces_1_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_39 = ces_1_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_40 = ces_1_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_41 = ces_1_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_42 = ces_1_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_43 = ces_1_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_44 = ces_1_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_45 = ces_1_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_46 = ces_1_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_47 = ces_1_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_48 = ces_1_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_49 = ces_1_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_50 = ces_1_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_51 = ces_1_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_52 = ces_1_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_53 = ces_1_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_54 = ces_1_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_55 = ces_1_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_56 = ces_1_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_57 = ces_1_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_58 = ces_1_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_59 = ces_1_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_60 = ces_1_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_61 = ces_1_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_62 = ces_1_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_63 = ces_1_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_64 = ces_2_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_65 = ces_2_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_66 = ces_2_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_67 = ces_2_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_68 = ces_2_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_69 = ces_2_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_70 = ces_2_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_71 = ces_2_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_72 = ces_2_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_73 = ces_2_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_74 = ces_2_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_75 = ces_2_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_76 = ces_2_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_77 = ces_2_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_78 = ces_2_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_79 = ces_2_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_80 = ces_2_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_81 = ces_2_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_82 = ces_2_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_83 = ces_2_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_84 = ces_2_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_85 = ces_2_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_86 = ces_2_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_87 = ces_2_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_88 = ces_2_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_89 = ces_2_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_90 = ces_2_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_91 = ces_2_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_92 = ces_2_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_93 = ces_2_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_94 = ces_2_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_95 = ces_2_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_96 = ces_3_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_97 = ces_3_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_98 = ces_3_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_99 = ces_3_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_100 = ces_3_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_101 = ces_3_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_102 = ces_3_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_103 = ces_3_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_104 = ces_3_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_105 = ces_3_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_106 = ces_3_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_107 = ces_3_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_108 = ces_3_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_109 = ces_3_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_110 = ces_3_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_111 = ces_3_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_112 = ces_3_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_113 = ces_3_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_114 = ces_3_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_115 = ces_3_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_116 = ces_3_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_117 = ces_3_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_118 = ces_3_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_119 = ces_3_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_120 = ces_3_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_121 = ces_3_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_122 = ces_3_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_123 = ces_3_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_124 = ces_3_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_125 = ces_3_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_126 = ces_3_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_127 = ces_3_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_128 = ces_4_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_129 = ces_4_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_130 = ces_4_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_131 = ces_4_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_132 = ces_4_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_133 = ces_4_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_134 = ces_4_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_135 = ces_4_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_136 = ces_4_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_137 = ces_4_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_138 = ces_4_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_139 = ces_4_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_140 = ces_4_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_141 = ces_4_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_142 = ces_4_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_143 = ces_4_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_144 = ces_4_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_145 = ces_4_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_146 = ces_4_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_147 = ces_4_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_148 = ces_4_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_149 = ces_4_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_150 = ces_4_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_151 = ces_4_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_152 = ces_4_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_153 = ces_4_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_154 = ces_4_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_155 = ces_4_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_156 = ces_4_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_157 = ces_4_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_158 = ces_4_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_159 = ces_4_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_160 = ces_5_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_161 = ces_5_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_162 = ces_5_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_163 = ces_5_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_164 = ces_5_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_165 = ces_5_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_166 = ces_5_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_167 = ces_5_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_168 = ces_5_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_169 = ces_5_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_170 = ces_5_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_171 = ces_5_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_172 = ces_5_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_173 = ces_5_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_174 = ces_5_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_175 = ces_5_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_176 = ces_5_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_177 = ces_5_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_178 = ces_5_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_179 = ces_5_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_180 = ces_5_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_181 = ces_5_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_182 = ces_5_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_183 = ces_5_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_184 = ces_5_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_185 = ces_5_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_186 = ces_5_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_187 = ces_5_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_188 = ces_5_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_189 = ces_5_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_190 = ces_5_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_191 = ces_5_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_192 = ces_6_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_193 = ces_6_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_194 = ces_6_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_195 = ces_6_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_196 = ces_6_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_197 = ces_6_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_198 = ces_6_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_199 = ces_6_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_200 = ces_6_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_201 = ces_6_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_202 = ces_6_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_203 = ces_6_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_204 = ces_6_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_205 = ces_6_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_206 = ces_6_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_207 = ces_6_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_208 = ces_6_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_209 = ces_6_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_210 = ces_6_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_211 = ces_6_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_212 = ces_6_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_213 = ces_6_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_214 = ces_6_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_215 = ces_6_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_216 = ces_6_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_217 = ces_6_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_218 = ces_6_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_219 = ces_6_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_220 = ces_6_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_221 = ces_6_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_222 = ces_6_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_223 = ces_6_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_224 = ces_7_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_225 = ces_7_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_226 = ces_7_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_227 = ces_7_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_228 = ces_7_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_229 = ces_7_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_230 = ces_7_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_231 = ces_7_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_232 = ces_7_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_233 = ces_7_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_234 = ces_7_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_235 = ces_7_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_236 = ces_7_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_237 = ces_7_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_238 = ces_7_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_239 = ces_7_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_240 = ces_7_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_241 = ces_7_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_242 = ces_7_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_243 = ces_7_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_244 = ces_7_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_245 = ces_7_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_246 = ces_7_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_247 = ces_7_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_248 = ces_7_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_249 = ces_7_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_250 = ces_7_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_251 = ces_7_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_252 = ces_7_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_253 = ces_7_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_254 = ces_7_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_255 = ces_7_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_256 = ces_8_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_257 = ces_8_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_258 = ces_8_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_259 = ces_8_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_260 = ces_8_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_261 = ces_8_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_262 = ces_8_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_263 = ces_8_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_264 = ces_8_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_265 = ces_8_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_266 = ces_8_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_267 = ces_8_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_268 = ces_8_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_269 = ces_8_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_270 = ces_8_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_271 = ces_8_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_272 = ces_8_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_273 = ces_8_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_274 = ces_8_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_275 = ces_8_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_276 = ces_8_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_277 = ces_8_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_278 = ces_8_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_279 = ces_8_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_280 = ces_8_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_281 = ces_8_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_282 = ces_8_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_283 = ces_8_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_284 = ces_8_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_285 = ces_8_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_286 = ces_8_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_287 = ces_8_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_288 = ces_9_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_289 = ces_9_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_290 = ces_9_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_291 = ces_9_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_292 = ces_9_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_293 = ces_9_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_294 = ces_9_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_295 = ces_9_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_296 = ces_9_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_297 = ces_9_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_298 = ces_9_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_299 = ces_9_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_300 = ces_9_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_301 = ces_9_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_302 = ces_9_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_303 = ces_9_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_304 = ces_9_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_305 = ces_9_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_306 = ces_9_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_307 = ces_9_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_308 = ces_9_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_309 = ces_9_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_310 = ces_9_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_311 = ces_9_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_312 = ces_9_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_313 = ces_9_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_314 = ces_9_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_315 = ces_9_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_316 = ces_9_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_317 = ces_9_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_318 = ces_9_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_319 = ces_9_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_320 = ces_10_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_321 = ces_10_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_322 = ces_10_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_323 = ces_10_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_324 = ces_10_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_325 = ces_10_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_326 = ces_10_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_327 = ces_10_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_328 = ces_10_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_329 = ces_10_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_330 = ces_10_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_331 = ces_10_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_332 = ces_10_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_333 = ces_10_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_334 = ces_10_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_335 = ces_10_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_336 = ces_10_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_337 = ces_10_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_338 = ces_10_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_339 = ces_10_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_340 = ces_10_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_341 = ces_10_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_342 = ces_10_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_343 = ces_10_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_344 = ces_10_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_345 = ces_10_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_346 = ces_10_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_347 = ces_10_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_348 = ces_10_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_349 = ces_10_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_350 = ces_10_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_351 = ces_10_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_352 = ces_11_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_353 = ces_11_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_354 = ces_11_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_355 = ces_11_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_356 = ces_11_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_357 = ces_11_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_358 = ces_11_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_359 = ces_11_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_360 = ces_11_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_361 = ces_11_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_362 = ces_11_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_363 = ces_11_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_364 = ces_11_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_365 = ces_11_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_366 = ces_11_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_367 = ces_11_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_368 = ces_11_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_369 = ces_11_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_370 = ces_11_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_371 = ces_11_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_372 = ces_11_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_373 = ces_11_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_374 = ces_11_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_375 = ces_11_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_376 = ces_11_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_377 = ces_11_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_378 = ces_11_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_379 = ces_11_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_380 = ces_11_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_381 = ces_11_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_382 = ces_11_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_383 = ces_11_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_384 = ces_12_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_385 = ces_12_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_386 = ces_12_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_387 = ces_12_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_388 = ces_12_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_389 = ces_12_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_390 = ces_12_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_391 = ces_12_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_392 = ces_12_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_393 = ces_12_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_394 = ces_12_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_395 = ces_12_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_396 = ces_12_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_397 = ces_12_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_398 = ces_12_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_399 = ces_12_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_400 = ces_12_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_401 = ces_12_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_402 = ces_12_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_403 = ces_12_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_404 = ces_12_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_405 = ces_12_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_406 = ces_12_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_407 = ces_12_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_408 = ces_12_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_409 = ces_12_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_410 = ces_12_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_411 = ces_12_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_412 = ces_12_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_413 = ces_12_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_414 = ces_12_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_415 = ces_12_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_416 = ces_13_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_417 = ces_13_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_418 = ces_13_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_419 = ces_13_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_420 = ces_13_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_421 = ces_13_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_422 = ces_13_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_423 = ces_13_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_424 = ces_13_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_425 = ces_13_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_426 = ces_13_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_427 = ces_13_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_428 = ces_13_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_429 = ces_13_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_430 = ces_13_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_431 = ces_13_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_432 = ces_13_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_433 = ces_13_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_434 = ces_13_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_435 = ces_13_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_436 = ces_13_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_437 = ces_13_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_438 = ces_13_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_439 = ces_13_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_440 = ces_13_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_441 = ces_13_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_442 = ces_13_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_443 = ces_13_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_444 = ces_13_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_445 = ces_13_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_446 = ces_13_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_447 = ces_13_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_448 = ces_14_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_449 = ces_14_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_450 = ces_14_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_451 = ces_14_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_452 = ces_14_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_453 = ces_14_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_454 = ces_14_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_455 = ces_14_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_456 = ces_14_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_457 = ces_14_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_458 = ces_14_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_459 = ces_14_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_460 = ces_14_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_461 = ces_14_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_462 = ces_14_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_463 = ces_14_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_464 = ces_14_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_465 = ces_14_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_466 = ces_14_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_467 = ces_14_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_468 = ces_14_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_469 = ces_14_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_470 = ces_14_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_471 = ces_14_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_472 = ces_14_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_473 = ces_14_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_474 = ces_14_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_475 = ces_14_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_476 = ces_14_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_477 = ces_14_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_478 = ces_14_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_479 = ces_14_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_480 = ces_15_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_481 = ces_15_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_482 = ces_15_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_483 = ces_15_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_484 = ces_15_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_485 = ces_15_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_486 = ces_15_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_487 = ces_15_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_488 = ces_15_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_489 = ces_15_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_490 = ces_15_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_491 = ces_15_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_492 = ces_15_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_493 = ces_15_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_494 = ces_15_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_495 = ces_15_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_496 = ces_15_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_497 = ces_15_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_498 = ces_15_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_499 = ces_15_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_500 = ces_15_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_501 = ces_15_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_502 = ces_15_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_503 = ces_15_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_504 = ces_15_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_505 = ces_15_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_506 = ces_15_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_507 = ces_15_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_508 = ces_15_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_509 = ces_15_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_510 = ces_15_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_511 = ces_15_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_512 = ces_16_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_513 = ces_16_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_514 = ces_16_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_515 = ces_16_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_516 = ces_16_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_517 = ces_16_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_518 = ces_16_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_519 = ces_16_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_520 = ces_16_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_521 = ces_16_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_522 = ces_16_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_523 = ces_16_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_524 = ces_16_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_525 = ces_16_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_526 = ces_16_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_527 = ces_16_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_528 = ces_16_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_529 = ces_16_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_530 = ces_16_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_531 = ces_16_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_532 = ces_16_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_533 = ces_16_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_534 = ces_16_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_535 = ces_16_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_536 = ces_16_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_537 = ces_16_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_538 = ces_16_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_539 = ces_16_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_540 = ces_16_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_541 = ces_16_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_542 = ces_16_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_543 = ces_16_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_544 = ces_17_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_545 = ces_17_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_546 = ces_17_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_547 = ces_17_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_548 = ces_17_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_549 = ces_17_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_550 = ces_17_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_551 = ces_17_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_552 = ces_17_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_553 = ces_17_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_554 = ces_17_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_555 = ces_17_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_556 = ces_17_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_557 = ces_17_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_558 = ces_17_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_559 = ces_17_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_560 = ces_17_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_561 = ces_17_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_562 = ces_17_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_563 = ces_17_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_564 = ces_17_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_565 = ces_17_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_566 = ces_17_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_567 = ces_17_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_568 = ces_17_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_569 = ces_17_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_570 = ces_17_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_571 = ces_17_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_572 = ces_17_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_573 = ces_17_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_574 = ces_17_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_575 = ces_17_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_576 = ces_18_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_577 = ces_18_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_578 = ces_18_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_579 = ces_18_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_580 = ces_18_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_581 = ces_18_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_582 = ces_18_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_583 = ces_18_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_584 = ces_18_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_585 = ces_18_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_586 = ces_18_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_587 = ces_18_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_588 = ces_18_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_589 = ces_18_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_590 = ces_18_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_591 = ces_18_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_592 = ces_18_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_593 = ces_18_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_594 = ces_18_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_595 = ces_18_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_596 = ces_18_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_597 = ces_18_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_598 = ces_18_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_599 = ces_18_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_600 = ces_18_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_601 = ces_18_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_602 = ces_18_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_603 = ces_18_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_604 = ces_18_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_605 = ces_18_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_606 = ces_18_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_607 = ces_18_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_608 = ces_19_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_609 = ces_19_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_610 = ces_19_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_611 = ces_19_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_612 = ces_19_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_613 = ces_19_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_614 = ces_19_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_615 = ces_19_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_616 = ces_19_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_617 = ces_19_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_618 = ces_19_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_619 = ces_19_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_620 = ces_19_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_621 = ces_19_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_622 = ces_19_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_623 = ces_19_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_624 = ces_19_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_625 = ces_19_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_626 = ces_19_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_627 = ces_19_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_628 = ces_19_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_629 = ces_19_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_630 = ces_19_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_631 = ces_19_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_632 = ces_19_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_633 = ces_19_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_634 = ces_19_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_635 = ces_19_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_636 = ces_19_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_637 = ces_19_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_638 = ces_19_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_639 = ces_19_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_640 = ces_20_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_641 = ces_20_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_642 = ces_20_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_643 = ces_20_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_644 = ces_20_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_645 = ces_20_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_646 = ces_20_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_647 = ces_20_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_648 = ces_20_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_649 = ces_20_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_650 = ces_20_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_651 = ces_20_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_652 = ces_20_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_653 = ces_20_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_654 = ces_20_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_655 = ces_20_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_656 = ces_20_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_657 = ces_20_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_658 = ces_20_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_659 = ces_20_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_660 = ces_20_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_661 = ces_20_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_662 = ces_20_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_663 = ces_20_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_664 = ces_20_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_665 = ces_20_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_666 = ces_20_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_667 = ces_20_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_668 = ces_20_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_669 = ces_20_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_670 = ces_20_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_671 = ces_20_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_672 = ces_21_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_673 = ces_21_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_674 = ces_21_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_675 = ces_21_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_676 = ces_21_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_677 = ces_21_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_678 = ces_21_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_679 = ces_21_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_680 = ces_21_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_681 = ces_21_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_682 = ces_21_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_683 = ces_21_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_684 = ces_21_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_685 = ces_21_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_686 = ces_21_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_687 = ces_21_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_688 = ces_21_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_689 = ces_21_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_690 = ces_21_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_691 = ces_21_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_692 = ces_21_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_693 = ces_21_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_694 = ces_21_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_695 = ces_21_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_696 = ces_21_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_697 = ces_21_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_698 = ces_21_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_699 = ces_21_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_700 = ces_21_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_701 = ces_21_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_702 = ces_21_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_703 = ces_21_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_704 = ces_22_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_705 = ces_22_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_706 = ces_22_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_707 = ces_22_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_708 = ces_22_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_709 = ces_22_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_710 = ces_22_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_711 = ces_22_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_712 = ces_22_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_713 = ces_22_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_714 = ces_22_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_715 = ces_22_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_716 = ces_22_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_717 = ces_22_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_718 = ces_22_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_719 = ces_22_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_720 = ces_22_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_721 = ces_22_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_722 = ces_22_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_723 = ces_22_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_724 = ces_22_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_725 = ces_22_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_726 = ces_22_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_727 = ces_22_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_728 = ces_22_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_729 = ces_22_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_730 = ces_22_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_731 = ces_22_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_732 = ces_22_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_733 = ces_22_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_734 = ces_22_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_735 = ces_22_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_736 = ces_23_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_737 = ces_23_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_738 = ces_23_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_739 = ces_23_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_740 = ces_23_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_741 = ces_23_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_742 = ces_23_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_743 = ces_23_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_744 = ces_23_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_745 = ces_23_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_746 = ces_23_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_747 = ces_23_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_748 = ces_23_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_749 = ces_23_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_750 = ces_23_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_751 = ces_23_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_752 = ces_23_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_753 = ces_23_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_754 = ces_23_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_755 = ces_23_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_756 = ces_23_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_757 = ces_23_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_758 = ces_23_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_759 = ces_23_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_760 = ces_23_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_761 = ces_23_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_762 = ces_23_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_763 = ces_23_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_764 = ces_23_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_765 = ces_23_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_766 = ces_23_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_767 = ces_23_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_768 = ces_24_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_769 = ces_24_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_770 = ces_24_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_771 = ces_24_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_772 = ces_24_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_773 = ces_24_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_774 = ces_24_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_775 = ces_24_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_776 = ces_24_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_777 = ces_24_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_778 = ces_24_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_779 = ces_24_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_780 = ces_24_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_781 = ces_24_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_782 = ces_24_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_783 = ces_24_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_784 = ces_24_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_785 = ces_24_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_786 = ces_24_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_787 = ces_24_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_788 = ces_24_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_789 = ces_24_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_790 = ces_24_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_791 = ces_24_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_792 = ces_24_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_793 = ces_24_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_794 = ces_24_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_795 = ces_24_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_796 = ces_24_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_797 = ces_24_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_798 = ces_24_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_799 = ces_24_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_800 = ces_25_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_801 = ces_25_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_802 = ces_25_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_803 = ces_25_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_804 = ces_25_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_805 = ces_25_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_806 = ces_25_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_807 = ces_25_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_808 = ces_25_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_809 = ces_25_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_810 = ces_25_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_811 = ces_25_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_812 = ces_25_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_813 = ces_25_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_814 = ces_25_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_815 = ces_25_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_816 = ces_25_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_817 = ces_25_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_818 = ces_25_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_819 = ces_25_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_820 = ces_25_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_821 = ces_25_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_822 = ces_25_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_823 = ces_25_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_824 = ces_25_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_825 = ces_25_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_826 = ces_25_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_827 = ces_25_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_828 = ces_25_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_829 = ces_25_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_830 = ces_25_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_831 = ces_25_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_832 = ces_26_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_833 = ces_26_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_834 = ces_26_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_835 = ces_26_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_836 = ces_26_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_837 = ces_26_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_838 = ces_26_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_839 = ces_26_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_840 = ces_26_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_841 = ces_26_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_842 = ces_26_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_843 = ces_26_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_844 = ces_26_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_845 = ces_26_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_846 = ces_26_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_847 = ces_26_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_848 = ces_26_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_849 = ces_26_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_850 = ces_26_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_851 = ces_26_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_852 = ces_26_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_853 = ces_26_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_854 = ces_26_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_855 = ces_26_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_856 = ces_26_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_857 = ces_26_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_858 = ces_26_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_859 = ces_26_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_860 = ces_26_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_861 = ces_26_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_862 = ces_26_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_863 = ces_26_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_864 = ces_27_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_865 = ces_27_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_866 = ces_27_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_867 = ces_27_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_868 = ces_27_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_869 = ces_27_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_870 = ces_27_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_871 = ces_27_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_872 = ces_27_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_873 = ces_27_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_874 = ces_27_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_875 = ces_27_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_876 = ces_27_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_877 = ces_27_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_878 = ces_27_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_879 = ces_27_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_880 = ces_27_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_881 = ces_27_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_882 = ces_27_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_883 = ces_27_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_884 = ces_27_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_885 = ces_27_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_886 = ces_27_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_887 = ces_27_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_888 = ces_27_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_889 = ces_27_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_890 = ces_27_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_891 = ces_27_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_892 = ces_27_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_893 = ces_27_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_894 = ces_27_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_895 = ces_27_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_896 = ces_28_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_897 = ces_28_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_898 = ces_28_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_899 = ces_28_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_900 = ces_28_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_901 = ces_28_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_902 = ces_28_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_903 = ces_28_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_904 = ces_28_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_905 = ces_28_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_906 = ces_28_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_907 = ces_28_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_908 = ces_28_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_909 = ces_28_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_910 = ces_28_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_911 = ces_28_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_912 = ces_28_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_913 = ces_28_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_914 = ces_28_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_915 = ces_28_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_916 = ces_28_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_917 = ces_28_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_918 = ces_28_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_919 = ces_28_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_920 = ces_28_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_921 = ces_28_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_922 = ces_28_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_923 = ces_28_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_924 = ces_28_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_925 = ces_28_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_926 = ces_28_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_927 = ces_28_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_928 = ces_29_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_929 = ces_29_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_930 = ces_29_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_931 = ces_29_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_932 = ces_29_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_933 = ces_29_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_934 = ces_29_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_935 = ces_29_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_936 = ces_29_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_937 = ces_29_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_938 = ces_29_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_939 = ces_29_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_940 = ces_29_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_941 = ces_29_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_942 = ces_29_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_943 = ces_29_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_944 = ces_29_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_945 = ces_29_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_946 = ces_29_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_947 = ces_29_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_948 = ces_29_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_949 = ces_29_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_950 = ces_29_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_951 = ces_29_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_952 = ces_29_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_953 = ces_29_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_954 = ces_29_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_955 = ces_29_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_956 = ces_29_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_957 = ces_29_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_958 = ces_29_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_959 = ces_29_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_960 = ces_30_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_961 = ces_30_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_962 = ces_30_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_963 = ces_30_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_964 = ces_30_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_965 = ces_30_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_966 = ces_30_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_967 = ces_30_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_968 = ces_30_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_969 = ces_30_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_970 = ces_30_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_971 = ces_30_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_972 = ces_30_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_973 = ces_30_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_974 = ces_30_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_975 = ces_30_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_976 = ces_30_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_977 = ces_30_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_978 = ces_30_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_979 = ces_30_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_980 = ces_30_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_981 = ces_30_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_982 = ces_30_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_983 = ces_30_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_984 = ces_30_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_985 = ces_30_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_986 = ces_30_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_987 = ces_30_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_988 = ces_30_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_989 = ces_30_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_990 = ces_30_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_991 = ces_30_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_992 = ces_31_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_993 = ces_31_1_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_994 = ces_31_2_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_995 = ces_31_3_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_996 = ces_31_4_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_997 = ces_31_5_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_998 = ces_31_6_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_999 = ces_31_7_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1000 = ces_31_8_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1001 = ces_31_9_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1002 = ces_31_10_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1003 = ces_31_11_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1004 = ces_31_12_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1005 = ces_31_13_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1006 = ces_31_14_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1007 = ces_31_15_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1008 = ces_31_16_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1009 = ces_31_17_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1010 = ces_31_18_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1011 = ces_31_19_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1012 = ces_31_20_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1013 = ces_31_21_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1014 = ces_31_22_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1015 = ces_31_23_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1016 = ces_31_24_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1017 = ces_31_25_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1018 = ces_31_26_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1019 = ces_31_27_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1020 = ces_31_28_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1021 = ces_31_29_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1022 = ces_31_30_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1023 = ces_31_31_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign ces_0_0_clock = clock;
  assign ces_0_0_io_ins_0 = io_insHorizontal_0_0; // @[MockArray.scala 44:87]
  assign ces_0_0_io_ins_1 = ces_0_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_0_io_ins_2 = ces_1_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_0_io_ins_3 = io_insVertical_1_0; // @[MockArray.scala 47:87]
  assign ces_0_1_clock = clock;
  assign ces_0_1_io_ins_0 = io_insHorizontal_0_1; // @[MockArray.scala 44:87]
  assign ces_0_1_io_ins_1 = ces_0_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_1_io_ins_2 = ces_1_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_1_io_ins_3 = ces_0_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_2_clock = clock;
  assign ces_0_2_io_ins_0 = io_insHorizontal_0_2; // @[MockArray.scala 44:87]
  assign ces_0_2_io_ins_1 = ces_0_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_2_io_ins_2 = ces_1_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_2_io_ins_3 = ces_0_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_3_clock = clock;
  assign ces_0_3_io_ins_0 = io_insHorizontal_0_3; // @[MockArray.scala 44:87]
  assign ces_0_3_io_ins_1 = ces_0_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_3_io_ins_2 = ces_1_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_3_io_ins_3 = ces_0_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_4_clock = clock;
  assign ces_0_4_io_ins_0 = io_insHorizontal_0_4; // @[MockArray.scala 44:87]
  assign ces_0_4_io_ins_1 = ces_0_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_4_io_ins_2 = ces_1_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_4_io_ins_3 = ces_0_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_5_clock = clock;
  assign ces_0_5_io_ins_0 = io_insHorizontal_0_5; // @[MockArray.scala 44:87]
  assign ces_0_5_io_ins_1 = ces_0_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_5_io_ins_2 = ces_1_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_5_io_ins_3 = ces_0_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_6_clock = clock;
  assign ces_0_6_io_ins_0 = io_insHorizontal_0_6; // @[MockArray.scala 44:87]
  assign ces_0_6_io_ins_1 = ces_0_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_6_io_ins_2 = ces_1_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_6_io_ins_3 = ces_0_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_7_clock = clock;
  assign ces_0_7_io_ins_0 = io_insHorizontal_0_7; // @[MockArray.scala 44:87]
  assign ces_0_7_io_ins_1 = ces_0_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_7_io_ins_2 = ces_1_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_7_io_ins_3 = ces_0_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_8_clock = clock;
  assign ces_0_8_io_ins_0 = io_insHorizontal_0_8; // @[MockArray.scala 44:87]
  assign ces_0_8_io_ins_1 = ces_0_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_8_io_ins_2 = ces_1_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_8_io_ins_3 = ces_0_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_9_clock = clock;
  assign ces_0_9_io_ins_0 = io_insHorizontal_0_9; // @[MockArray.scala 44:87]
  assign ces_0_9_io_ins_1 = ces_0_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_9_io_ins_2 = ces_1_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_9_io_ins_3 = ces_0_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_10_clock = clock;
  assign ces_0_10_io_ins_0 = io_insHorizontal_0_10; // @[MockArray.scala 44:87]
  assign ces_0_10_io_ins_1 = ces_0_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_10_io_ins_2 = ces_1_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_10_io_ins_3 = ces_0_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_11_clock = clock;
  assign ces_0_11_io_ins_0 = io_insHorizontal_0_11; // @[MockArray.scala 44:87]
  assign ces_0_11_io_ins_1 = ces_0_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_11_io_ins_2 = ces_1_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_11_io_ins_3 = ces_0_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_12_clock = clock;
  assign ces_0_12_io_ins_0 = io_insHorizontal_0_12; // @[MockArray.scala 44:87]
  assign ces_0_12_io_ins_1 = ces_0_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_12_io_ins_2 = ces_1_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_12_io_ins_3 = ces_0_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_13_clock = clock;
  assign ces_0_13_io_ins_0 = io_insHorizontal_0_13; // @[MockArray.scala 44:87]
  assign ces_0_13_io_ins_1 = ces_0_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_13_io_ins_2 = ces_1_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_13_io_ins_3 = ces_0_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_14_clock = clock;
  assign ces_0_14_io_ins_0 = io_insHorizontal_0_14; // @[MockArray.scala 44:87]
  assign ces_0_14_io_ins_1 = ces_0_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_14_io_ins_2 = ces_1_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_14_io_ins_3 = ces_0_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_15_clock = clock;
  assign ces_0_15_io_ins_0 = io_insHorizontal_0_15; // @[MockArray.scala 44:87]
  assign ces_0_15_io_ins_1 = ces_0_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_15_io_ins_2 = ces_1_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_15_io_ins_3 = ces_0_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_16_clock = clock;
  assign ces_0_16_io_ins_0 = io_insHorizontal_0_16; // @[MockArray.scala 44:87]
  assign ces_0_16_io_ins_1 = ces_0_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_16_io_ins_2 = ces_1_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_16_io_ins_3 = ces_0_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_17_clock = clock;
  assign ces_0_17_io_ins_0 = io_insHorizontal_0_17; // @[MockArray.scala 44:87]
  assign ces_0_17_io_ins_1 = ces_0_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_17_io_ins_2 = ces_1_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_17_io_ins_3 = ces_0_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_18_clock = clock;
  assign ces_0_18_io_ins_0 = io_insHorizontal_0_18; // @[MockArray.scala 44:87]
  assign ces_0_18_io_ins_1 = ces_0_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_18_io_ins_2 = ces_1_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_18_io_ins_3 = ces_0_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_19_clock = clock;
  assign ces_0_19_io_ins_0 = io_insHorizontal_0_19; // @[MockArray.scala 44:87]
  assign ces_0_19_io_ins_1 = ces_0_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_19_io_ins_2 = ces_1_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_19_io_ins_3 = ces_0_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_20_clock = clock;
  assign ces_0_20_io_ins_0 = io_insHorizontal_0_20; // @[MockArray.scala 44:87]
  assign ces_0_20_io_ins_1 = ces_0_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_20_io_ins_2 = ces_1_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_20_io_ins_3 = ces_0_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_21_clock = clock;
  assign ces_0_21_io_ins_0 = io_insHorizontal_0_21; // @[MockArray.scala 44:87]
  assign ces_0_21_io_ins_1 = ces_0_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_21_io_ins_2 = ces_1_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_21_io_ins_3 = ces_0_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_22_clock = clock;
  assign ces_0_22_io_ins_0 = io_insHorizontal_0_22; // @[MockArray.scala 44:87]
  assign ces_0_22_io_ins_1 = ces_0_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_22_io_ins_2 = ces_1_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_22_io_ins_3 = ces_0_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_23_clock = clock;
  assign ces_0_23_io_ins_0 = io_insHorizontal_0_23; // @[MockArray.scala 44:87]
  assign ces_0_23_io_ins_1 = ces_0_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_23_io_ins_2 = ces_1_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_23_io_ins_3 = ces_0_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_24_clock = clock;
  assign ces_0_24_io_ins_0 = io_insHorizontal_0_24; // @[MockArray.scala 44:87]
  assign ces_0_24_io_ins_1 = ces_0_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_24_io_ins_2 = ces_1_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_24_io_ins_3 = ces_0_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_25_clock = clock;
  assign ces_0_25_io_ins_0 = io_insHorizontal_0_25; // @[MockArray.scala 44:87]
  assign ces_0_25_io_ins_1 = ces_0_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_25_io_ins_2 = ces_1_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_25_io_ins_3 = ces_0_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_26_clock = clock;
  assign ces_0_26_io_ins_0 = io_insHorizontal_0_26; // @[MockArray.scala 44:87]
  assign ces_0_26_io_ins_1 = ces_0_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_26_io_ins_2 = ces_1_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_26_io_ins_3 = ces_0_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_27_clock = clock;
  assign ces_0_27_io_ins_0 = io_insHorizontal_0_27; // @[MockArray.scala 44:87]
  assign ces_0_27_io_ins_1 = ces_0_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_27_io_ins_2 = ces_1_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_27_io_ins_3 = ces_0_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_28_clock = clock;
  assign ces_0_28_io_ins_0 = io_insHorizontal_0_28; // @[MockArray.scala 44:87]
  assign ces_0_28_io_ins_1 = ces_0_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_28_io_ins_2 = ces_1_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_28_io_ins_3 = ces_0_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_29_clock = clock;
  assign ces_0_29_io_ins_0 = io_insHorizontal_0_29; // @[MockArray.scala 44:87]
  assign ces_0_29_io_ins_1 = ces_0_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_29_io_ins_2 = ces_1_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_29_io_ins_3 = ces_0_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_30_clock = clock;
  assign ces_0_30_io_ins_0 = io_insHorizontal_0_30; // @[MockArray.scala 44:87]
  assign ces_0_30_io_ins_1 = ces_0_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_0_30_io_ins_2 = ces_1_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_30_io_ins_3 = ces_0_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_0_31_clock = clock;
  assign ces_0_31_io_ins_0 = io_insHorizontal_0_31; // @[MockArray.scala 44:87]
  assign ces_0_31_io_ins_1 = io_insVertical_0_0; // @[MockArray.scala 45:87]
  assign ces_0_31_io_ins_2 = ces_1_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_31_io_ins_3 = ces_0_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_0_clock = clock;
  assign ces_1_0_io_ins_0 = ces_0_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_0_io_ins_1 = ces_1_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_0_io_ins_2 = ces_2_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_0_io_ins_3 = io_insVertical_1_1; // @[MockArray.scala 47:87]
  assign ces_1_1_clock = clock;
  assign ces_1_1_io_ins_0 = ces_0_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_1_io_ins_1 = ces_1_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_1_io_ins_2 = ces_2_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_1_io_ins_3 = ces_1_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_2_clock = clock;
  assign ces_1_2_io_ins_0 = ces_0_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_2_io_ins_1 = ces_1_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_2_io_ins_2 = ces_2_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_2_io_ins_3 = ces_1_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_3_clock = clock;
  assign ces_1_3_io_ins_0 = ces_0_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_3_io_ins_1 = ces_1_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_3_io_ins_2 = ces_2_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_3_io_ins_3 = ces_1_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_4_clock = clock;
  assign ces_1_4_io_ins_0 = ces_0_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_4_io_ins_1 = ces_1_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_4_io_ins_2 = ces_2_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_4_io_ins_3 = ces_1_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_5_clock = clock;
  assign ces_1_5_io_ins_0 = ces_0_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_5_io_ins_1 = ces_1_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_5_io_ins_2 = ces_2_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_5_io_ins_3 = ces_1_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_6_clock = clock;
  assign ces_1_6_io_ins_0 = ces_0_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_6_io_ins_1 = ces_1_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_6_io_ins_2 = ces_2_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_6_io_ins_3 = ces_1_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_7_clock = clock;
  assign ces_1_7_io_ins_0 = ces_0_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_7_io_ins_1 = ces_1_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_7_io_ins_2 = ces_2_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_7_io_ins_3 = ces_1_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_8_clock = clock;
  assign ces_1_8_io_ins_0 = ces_0_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_8_io_ins_1 = ces_1_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_8_io_ins_2 = ces_2_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_8_io_ins_3 = ces_1_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_9_clock = clock;
  assign ces_1_9_io_ins_0 = ces_0_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_9_io_ins_1 = ces_1_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_9_io_ins_2 = ces_2_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_9_io_ins_3 = ces_1_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_10_clock = clock;
  assign ces_1_10_io_ins_0 = ces_0_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_10_io_ins_1 = ces_1_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_10_io_ins_2 = ces_2_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_10_io_ins_3 = ces_1_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_11_clock = clock;
  assign ces_1_11_io_ins_0 = ces_0_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_11_io_ins_1 = ces_1_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_11_io_ins_2 = ces_2_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_11_io_ins_3 = ces_1_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_12_clock = clock;
  assign ces_1_12_io_ins_0 = ces_0_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_12_io_ins_1 = ces_1_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_12_io_ins_2 = ces_2_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_12_io_ins_3 = ces_1_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_13_clock = clock;
  assign ces_1_13_io_ins_0 = ces_0_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_13_io_ins_1 = ces_1_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_13_io_ins_2 = ces_2_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_13_io_ins_3 = ces_1_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_14_clock = clock;
  assign ces_1_14_io_ins_0 = ces_0_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_14_io_ins_1 = ces_1_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_14_io_ins_2 = ces_2_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_14_io_ins_3 = ces_1_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_15_clock = clock;
  assign ces_1_15_io_ins_0 = ces_0_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_15_io_ins_1 = ces_1_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_15_io_ins_2 = ces_2_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_15_io_ins_3 = ces_1_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_16_clock = clock;
  assign ces_1_16_io_ins_0 = ces_0_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_16_io_ins_1 = ces_1_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_16_io_ins_2 = ces_2_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_16_io_ins_3 = ces_1_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_17_clock = clock;
  assign ces_1_17_io_ins_0 = ces_0_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_17_io_ins_1 = ces_1_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_17_io_ins_2 = ces_2_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_17_io_ins_3 = ces_1_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_18_clock = clock;
  assign ces_1_18_io_ins_0 = ces_0_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_18_io_ins_1 = ces_1_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_18_io_ins_2 = ces_2_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_18_io_ins_3 = ces_1_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_19_clock = clock;
  assign ces_1_19_io_ins_0 = ces_0_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_19_io_ins_1 = ces_1_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_19_io_ins_2 = ces_2_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_19_io_ins_3 = ces_1_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_20_clock = clock;
  assign ces_1_20_io_ins_0 = ces_0_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_20_io_ins_1 = ces_1_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_20_io_ins_2 = ces_2_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_20_io_ins_3 = ces_1_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_21_clock = clock;
  assign ces_1_21_io_ins_0 = ces_0_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_21_io_ins_1 = ces_1_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_21_io_ins_2 = ces_2_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_21_io_ins_3 = ces_1_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_22_clock = clock;
  assign ces_1_22_io_ins_0 = ces_0_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_22_io_ins_1 = ces_1_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_22_io_ins_2 = ces_2_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_22_io_ins_3 = ces_1_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_23_clock = clock;
  assign ces_1_23_io_ins_0 = ces_0_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_23_io_ins_1 = ces_1_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_23_io_ins_2 = ces_2_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_23_io_ins_3 = ces_1_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_24_clock = clock;
  assign ces_1_24_io_ins_0 = ces_0_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_24_io_ins_1 = ces_1_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_24_io_ins_2 = ces_2_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_24_io_ins_3 = ces_1_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_25_clock = clock;
  assign ces_1_25_io_ins_0 = ces_0_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_25_io_ins_1 = ces_1_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_25_io_ins_2 = ces_2_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_25_io_ins_3 = ces_1_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_26_clock = clock;
  assign ces_1_26_io_ins_0 = ces_0_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_26_io_ins_1 = ces_1_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_26_io_ins_2 = ces_2_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_26_io_ins_3 = ces_1_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_27_clock = clock;
  assign ces_1_27_io_ins_0 = ces_0_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_27_io_ins_1 = ces_1_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_27_io_ins_2 = ces_2_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_27_io_ins_3 = ces_1_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_28_clock = clock;
  assign ces_1_28_io_ins_0 = ces_0_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_28_io_ins_1 = ces_1_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_28_io_ins_2 = ces_2_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_28_io_ins_3 = ces_1_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_29_clock = clock;
  assign ces_1_29_io_ins_0 = ces_0_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_29_io_ins_1 = ces_1_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_29_io_ins_2 = ces_2_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_29_io_ins_3 = ces_1_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_30_clock = clock;
  assign ces_1_30_io_ins_0 = ces_0_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_30_io_ins_1 = ces_1_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_1_30_io_ins_2 = ces_2_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_30_io_ins_3 = ces_1_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_1_31_clock = clock;
  assign ces_1_31_io_ins_0 = ces_0_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_31_io_ins_1 = io_insVertical_0_1; // @[MockArray.scala 45:87]
  assign ces_1_31_io_ins_2 = ces_2_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_31_io_ins_3 = ces_1_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_0_clock = clock;
  assign ces_2_0_io_ins_0 = ces_1_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_0_io_ins_1 = ces_2_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_0_io_ins_2 = ces_3_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_0_io_ins_3 = io_insVertical_1_2; // @[MockArray.scala 47:87]
  assign ces_2_1_clock = clock;
  assign ces_2_1_io_ins_0 = ces_1_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_1_io_ins_1 = ces_2_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_1_io_ins_2 = ces_3_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_1_io_ins_3 = ces_2_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_2_clock = clock;
  assign ces_2_2_io_ins_0 = ces_1_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_2_io_ins_1 = ces_2_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_2_io_ins_2 = ces_3_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_2_io_ins_3 = ces_2_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_3_clock = clock;
  assign ces_2_3_io_ins_0 = ces_1_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_3_io_ins_1 = ces_2_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_3_io_ins_2 = ces_3_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_3_io_ins_3 = ces_2_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_4_clock = clock;
  assign ces_2_4_io_ins_0 = ces_1_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_4_io_ins_1 = ces_2_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_4_io_ins_2 = ces_3_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_4_io_ins_3 = ces_2_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_5_clock = clock;
  assign ces_2_5_io_ins_0 = ces_1_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_5_io_ins_1 = ces_2_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_5_io_ins_2 = ces_3_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_5_io_ins_3 = ces_2_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_6_clock = clock;
  assign ces_2_6_io_ins_0 = ces_1_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_6_io_ins_1 = ces_2_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_6_io_ins_2 = ces_3_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_6_io_ins_3 = ces_2_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_7_clock = clock;
  assign ces_2_7_io_ins_0 = ces_1_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_7_io_ins_1 = ces_2_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_7_io_ins_2 = ces_3_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_7_io_ins_3 = ces_2_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_8_clock = clock;
  assign ces_2_8_io_ins_0 = ces_1_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_8_io_ins_1 = ces_2_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_8_io_ins_2 = ces_3_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_8_io_ins_3 = ces_2_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_9_clock = clock;
  assign ces_2_9_io_ins_0 = ces_1_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_9_io_ins_1 = ces_2_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_9_io_ins_2 = ces_3_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_9_io_ins_3 = ces_2_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_10_clock = clock;
  assign ces_2_10_io_ins_0 = ces_1_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_10_io_ins_1 = ces_2_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_10_io_ins_2 = ces_3_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_10_io_ins_3 = ces_2_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_11_clock = clock;
  assign ces_2_11_io_ins_0 = ces_1_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_11_io_ins_1 = ces_2_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_11_io_ins_2 = ces_3_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_11_io_ins_3 = ces_2_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_12_clock = clock;
  assign ces_2_12_io_ins_0 = ces_1_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_12_io_ins_1 = ces_2_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_12_io_ins_2 = ces_3_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_12_io_ins_3 = ces_2_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_13_clock = clock;
  assign ces_2_13_io_ins_0 = ces_1_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_13_io_ins_1 = ces_2_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_13_io_ins_2 = ces_3_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_13_io_ins_3 = ces_2_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_14_clock = clock;
  assign ces_2_14_io_ins_0 = ces_1_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_14_io_ins_1 = ces_2_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_14_io_ins_2 = ces_3_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_14_io_ins_3 = ces_2_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_15_clock = clock;
  assign ces_2_15_io_ins_0 = ces_1_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_15_io_ins_1 = ces_2_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_15_io_ins_2 = ces_3_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_15_io_ins_3 = ces_2_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_16_clock = clock;
  assign ces_2_16_io_ins_0 = ces_1_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_16_io_ins_1 = ces_2_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_16_io_ins_2 = ces_3_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_16_io_ins_3 = ces_2_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_17_clock = clock;
  assign ces_2_17_io_ins_0 = ces_1_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_17_io_ins_1 = ces_2_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_17_io_ins_2 = ces_3_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_17_io_ins_3 = ces_2_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_18_clock = clock;
  assign ces_2_18_io_ins_0 = ces_1_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_18_io_ins_1 = ces_2_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_18_io_ins_2 = ces_3_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_18_io_ins_3 = ces_2_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_19_clock = clock;
  assign ces_2_19_io_ins_0 = ces_1_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_19_io_ins_1 = ces_2_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_19_io_ins_2 = ces_3_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_19_io_ins_3 = ces_2_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_20_clock = clock;
  assign ces_2_20_io_ins_0 = ces_1_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_20_io_ins_1 = ces_2_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_20_io_ins_2 = ces_3_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_20_io_ins_3 = ces_2_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_21_clock = clock;
  assign ces_2_21_io_ins_0 = ces_1_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_21_io_ins_1 = ces_2_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_21_io_ins_2 = ces_3_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_21_io_ins_3 = ces_2_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_22_clock = clock;
  assign ces_2_22_io_ins_0 = ces_1_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_22_io_ins_1 = ces_2_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_22_io_ins_2 = ces_3_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_22_io_ins_3 = ces_2_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_23_clock = clock;
  assign ces_2_23_io_ins_0 = ces_1_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_23_io_ins_1 = ces_2_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_23_io_ins_2 = ces_3_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_23_io_ins_3 = ces_2_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_24_clock = clock;
  assign ces_2_24_io_ins_0 = ces_1_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_24_io_ins_1 = ces_2_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_24_io_ins_2 = ces_3_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_24_io_ins_3 = ces_2_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_25_clock = clock;
  assign ces_2_25_io_ins_0 = ces_1_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_25_io_ins_1 = ces_2_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_25_io_ins_2 = ces_3_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_25_io_ins_3 = ces_2_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_26_clock = clock;
  assign ces_2_26_io_ins_0 = ces_1_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_26_io_ins_1 = ces_2_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_26_io_ins_2 = ces_3_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_26_io_ins_3 = ces_2_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_27_clock = clock;
  assign ces_2_27_io_ins_0 = ces_1_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_27_io_ins_1 = ces_2_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_27_io_ins_2 = ces_3_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_27_io_ins_3 = ces_2_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_28_clock = clock;
  assign ces_2_28_io_ins_0 = ces_1_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_28_io_ins_1 = ces_2_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_28_io_ins_2 = ces_3_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_28_io_ins_3 = ces_2_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_29_clock = clock;
  assign ces_2_29_io_ins_0 = ces_1_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_29_io_ins_1 = ces_2_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_29_io_ins_2 = ces_3_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_29_io_ins_3 = ces_2_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_30_clock = clock;
  assign ces_2_30_io_ins_0 = ces_1_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_30_io_ins_1 = ces_2_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_2_30_io_ins_2 = ces_3_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_30_io_ins_3 = ces_2_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_2_31_clock = clock;
  assign ces_2_31_io_ins_0 = ces_1_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_31_io_ins_1 = io_insVertical_0_2; // @[MockArray.scala 45:87]
  assign ces_2_31_io_ins_2 = ces_3_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_31_io_ins_3 = ces_2_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_0_clock = clock;
  assign ces_3_0_io_ins_0 = ces_2_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_0_io_ins_1 = ces_3_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_0_io_ins_2 = ces_4_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_0_io_ins_3 = io_insVertical_1_3; // @[MockArray.scala 47:87]
  assign ces_3_1_clock = clock;
  assign ces_3_1_io_ins_0 = ces_2_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_1_io_ins_1 = ces_3_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_1_io_ins_2 = ces_4_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_1_io_ins_3 = ces_3_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_2_clock = clock;
  assign ces_3_2_io_ins_0 = ces_2_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_2_io_ins_1 = ces_3_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_2_io_ins_2 = ces_4_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_2_io_ins_3 = ces_3_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_3_clock = clock;
  assign ces_3_3_io_ins_0 = ces_2_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_3_io_ins_1 = ces_3_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_3_io_ins_2 = ces_4_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_3_io_ins_3 = ces_3_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_4_clock = clock;
  assign ces_3_4_io_ins_0 = ces_2_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_4_io_ins_1 = ces_3_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_4_io_ins_2 = ces_4_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_4_io_ins_3 = ces_3_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_5_clock = clock;
  assign ces_3_5_io_ins_0 = ces_2_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_5_io_ins_1 = ces_3_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_5_io_ins_2 = ces_4_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_5_io_ins_3 = ces_3_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_6_clock = clock;
  assign ces_3_6_io_ins_0 = ces_2_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_6_io_ins_1 = ces_3_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_6_io_ins_2 = ces_4_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_6_io_ins_3 = ces_3_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_7_clock = clock;
  assign ces_3_7_io_ins_0 = ces_2_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_7_io_ins_1 = ces_3_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_7_io_ins_2 = ces_4_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_7_io_ins_3 = ces_3_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_8_clock = clock;
  assign ces_3_8_io_ins_0 = ces_2_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_8_io_ins_1 = ces_3_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_8_io_ins_2 = ces_4_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_8_io_ins_3 = ces_3_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_9_clock = clock;
  assign ces_3_9_io_ins_0 = ces_2_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_9_io_ins_1 = ces_3_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_9_io_ins_2 = ces_4_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_9_io_ins_3 = ces_3_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_10_clock = clock;
  assign ces_3_10_io_ins_0 = ces_2_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_10_io_ins_1 = ces_3_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_10_io_ins_2 = ces_4_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_10_io_ins_3 = ces_3_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_11_clock = clock;
  assign ces_3_11_io_ins_0 = ces_2_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_11_io_ins_1 = ces_3_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_11_io_ins_2 = ces_4_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_11_io_ins_3 = ces_3_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_12_clock = clock;
  assign ces_3_12_io_ins_0 = ces_2_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_12_io_ins_1 = ces_3_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_12_io_ins_2 = ces_4_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_12_io_ins_3 = ces_3_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_13_clock = clock;
  assign ces_3_13_io_ins_0 = ces_2_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_13_io_ins_1 = ces_3_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_13_io_ins_2 = ces_4_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_13_io_ins_3 = ces_3_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_14_clock = clock;
  assign ces_3_14_io_ins_0 = ces_2_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_14_io_ins_1 = ces_3_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_14_io_ins_2 = ces_4_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_14_io_ins_3 = ces_3_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_15_clock = clock;
  assign ces_3_15_io_ins_0 = ces_2_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_15_io_ins_1 = ces_3_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_15_io_ins_2 = ces_4_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_15_io_ins_3 = ces_3_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_16_clock = clock;
  assign ces_3_16_io_ins_0 = ces_2_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_16_io_ins_1 = ces_3_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_16_io_ins_2 = ces_4_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_16_io_ins_3 = ces_3_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_17_clock = clock;
  assign ces_3_17_io_ins_0 = ces_2_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_17_io_ins_1 = ces_3_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_17_io_ins_2 = ces_4_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_17_io_ins_3 = ces_3_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_18_clock = clock;
  assign ces_3_18_io_ins_0 = ces_2_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_18_io_ins_1 = ces_3_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_18_io_ins_2 = ces_4_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_18_io_ins_3 = ces_3_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_19_clock = clock;
  assign ces_3_19_io_ins_0 = ces_2_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_19_io_ins_1 = ces_3_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_19_io_ins_2 = ces_4_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_19_io_ins_3 = ces_3_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_20_clock = clock;
  assign ces_3_20_io_ins_0 = ces_2_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_20_io_ins_1 = ces_3_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_20_io_ins_2 = ces_4_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_20_io_ins_3 = ces_3_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_21_clock = clock;
  assign ces_3_21_io_ins_0 = ces_2_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_21_io_ins_1 = ces_3_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_21_io_ins_2 = ces_4_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_21_io_ins_3 = ces_3_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_22_clock = clock;
  assign ces_3_22_io_ins_0 = ces_2_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_22_io_ins_1 = ces_3_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_22_io_ins_2 = ces_4_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_22_io_ins_3 = ces_3_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_23_clock = clock;
  assign ces_3_23_io_ins_0 = ces_2_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_23_io_ins_1 = ces_3_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_23_io_ins_2 = ces_4_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_23_io_ins_3 = ces_3_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_24_clock = clock;
  assign ces_3_24_io_ins_0 = ces_2_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_24_io_ins_1 = ces_3_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_24_io_ins_2 = ces_4_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_24_io_ins_3 = ces_3_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_25_clock = clock;
  assign ces_3_25_io_ins_0 = ces_2_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_25_io_ins_1 = ces_3_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_25_io_ins_2 = ces_4_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_25_io_ins_3 = ces_3_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_26_clock = clock;
  assign ces_3_26_io_ins_0 = ces_2_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_26_io_ins_1 = ces_3_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_26_io_ins_2 = ces_4_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_26_io_ins_3 = ces_3_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_27_clock = clock;
  assign ces_3_27_io_ins_0 = ces_2_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_27_io_ins_1 = ces_3_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_27_io_ins_2 = ces_4_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_27_io_ins_3 = ces_3_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_28_clock = clock;
  assign ces_3_28_io_ins_0 = ces_2_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_28_io_ins_1 = ces_3_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_28_io_ins_2 = ces_4_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_28_io_ins_3 = ces_3_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_29_clock = clock;
  assign ces_3_29_io_ins_0 = ces_2_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_29_io_ins_1 = ces_3_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_29_io_ins_2 = ces_4_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_29_io_ins_3 = ces_3_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_30_clock = clock;
  assign ces_3_30_io_ins_0 = ces_2_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_30_io_ins_1 = ces_3_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_3_30_io_ins_2 = ces_4_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_30_io_ins_3 = ces_3_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_3_31_clock = clock;
  assign ces_3_31_io_ins_0 = ces_2_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_31_io_ins_1 = io_insVertical_0_3; // @[MockArray.scala 45:87]
  assign ces_3_31_io_ins_2 = ces_4_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_31_io_ins_3 = ces_3_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_0_clock = clock;
  assign ces_4_0_io_ins_0 = ces_3_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_0_io_ins_1 = ces_4_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_0_io_ins_2 = ces_5_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_0_io_ins_3 = io_insVertical_1_4; // @[MockArray.scala 47:87]
  assign ces_4_1_clock = clock;
  assign ces_4_1_io_ins_0 = ces_3_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_1_io_ins_1 = ces_4_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_1_io_ins_2 = ces_5_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_1_io_ins_3 = ces_4_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_2_clock = clock;
  assign ces_4_2_io_ins_0 = ces_3_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_2_io_ins_1 = ces_4_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_2_io_ins_2 = ces_5_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_2_io_ins_3 = ces_4_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_3_clock = clock;
  assign ces_4_3_io_ins_0 = ces_3_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_3_io_ins_1 = ces_4_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_3_io_ins_2 = ces_5_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_3_io_ins_3 = ces_4_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_4_clock = clock;
  assign ces_4_4_io_ins_0 = ces_3_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_4_io_ins_1 = ces_4_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_4_io_ins_2 = ces_5_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_4_io_ins_3 = ces_4_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_5_clock = clock;
  assign ces_4_5_io_ins_0 = ces_3_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_5_io_ins_1 = ces_4_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_5_io_ins_2 = ces_5_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_5_io_ins_3 = ces_4_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_6_clock = clock;
  assign ces_4_6_io_ins_0 = ces_3_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_6_io_ins_1 = ces_4_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_6_io_ins_2 = ces_5_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_6_io_ins_3 = ces_4_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_7_clock = clock;
  assign ces_4_7_io_ins_0 = ces_3_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_7_io_ins_1 = ces_4_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_7_io_ins_2 = ces_5_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_7_io_ins_3 = ces_4_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_8_clock = clock;
  assign ces_4_8_io_ins_0 = ces_3_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_8_io_ins_1 = ces_4_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_8_io_ins_2 = ces_5_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_8_io_ins_3 = ces_4_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_9_clock = clock;
  assign ces_4_9_io_ins_0 = ces_3_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_9_io_ins_1 = ces_4_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_9_io_ins_2 = ces_5_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_9_io_ins_3 = ces_4_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_10_clock = clock;
  assign ces_4_10_io_ins_0 = ces_3_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_10_io_ins_1 = ces_4_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_10_io_ins_2 = ces_5_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_10_io_ins_3 = ces_4_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_11_clock = clock;
  assign ces_4_11_io_ins_0 = ces_3_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_11_io_ins_1 = ces_4_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_11_io_ins_2 = ces_5_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_11_io_ins_3 = ces_4_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_12_clock = clock;
  assign ces_4_12_io_ins_0 = ces_3_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_12_io_ins_1 = ces_4_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_12_io_ins_2 = ces_5_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_12_io_ins_3 = ces_4_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_13_clock = clock;
  assign ces_4_13_io_ins_0 = ces_3_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_13_io_ins_1 = ces_4_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_13_io_ins_2 = ces_5_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_13_io_ins_3 = ces_4_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_14_clock = clock;
  assign ces_4_14_io_ins_0 = ces_3_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_14_io_ins_1 = ces_4_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_14_io_ins_2 = ces_5_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_14_io_ins_3 = ces_4_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_15_clock = clock;
  assign ces_4_15_io_ins_0 = ces_3_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_15_io_ins_1 = ces_4_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_15_io_ins_2 = ces_5_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_15_io_ins_3 = ces_4_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_16_clock = clock;
  assign ces_4_16_io_ins_0 = ces_3_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_16_io_ins_1 = ces_4_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_16_io_ins_2 = ces_5_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_16_io_ins_3 = ces_4_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_17_clock = clock;
  assign ces_4_17_io_ins_0 = ces_3_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_17_io_ins_1 = ces_4_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_17_io_ins_2 = ces_5_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_17_io_ins_3 = ces_4_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_18_clock = clock;
  assign ces_4_18_io_ins_0 = ces_3_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_18_io_ins_1 = ces_4_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_18_io_ins_2 = ces_5_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_18_io_ins_3 = ces_4_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_19_clock = clock;
  assign ces_4_19_io_ins_0 = ces_3_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_19_io_ins_1 = ces_4_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_19_io_ins_2 = ces_5_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_19_io_ins_3 = ces_4_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_20_clock = clock;
  assign ces_4_20_io_ins_0 = ces_3_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_20_io_ins_1 = ces_4_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_20_io_ins_2 = ces_5_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_20_io_ins_3 = ces_4_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_21_clock = clock;
  assign ces_4_21_io_ins_0 = ces_3_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_21_io_ins_1 = ces_4_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_21_io_ins_2 = ces_5_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_21_io_ins_3 = ces_4_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_22_clock = clock;
  assign ces_4_22_io_ins_0 = ces_3_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_22_io_ins_1 = ces_4_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_22_io_ins_2 = ces_5_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_22_io_ins_3 = ces_4_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_23_clock = clock;
  assign ces_4_23_io_ins_0 = ces_3_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_23_io_ins_1 = ces_4_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_23_io_ins_2 = ces_5_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_23_io_ins_3 = ces_4_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_24_clock = clock;
  assign ces_4_24_io_ins_0 = ces_3_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_24_io_ins_1 = ces_4_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_24_io_ins_2 = ces_5_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_24_io_ins_3 = ces_4_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_25_clock = clock;
  assign ces_4_25_io_ins_0 = ces_3_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_25_io_ins_1 = ces_4_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_25_io_ins_2 = ces_5_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_25_io_ins_3 = ces_4_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_26_clock = clock;
  assign ces_4_26_io_ins_0 = ces_3_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_26_io_ins_1 = ces_4_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_26_io_ins_2 = ces_5_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_26_io_ins_3 = ces_4_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_27_clock = clock;
  assign ces_4_27_io_ins_0 = ces_3_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_27_io_ins_1 = ces_4_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_27_io_ins_2 = ces_5_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_27_io_ins_3 = ces_4_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_28_clock = clock;
  assign ces_4_28_io_ins_0 = ces_3_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_28_io_ins_1 = ces_4_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_28_io_ins_2 = ces_5_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_28_io_ins_3 = ces_4_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_29_clock = clock;
  assign ces_4_29_io_ins_0 = ces_3_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_29_io_ins_1 = ces_4_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_29_io_ins_2 = ces_5_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_29_io_ins_3 = ces_4_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_30_clock = clock;
  assign ces_4_30_io_ins_0 = ces_3_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_30_io_ins_1 = ces_4_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_4_30_io_ins_2 = ces_5_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_30_io_ins_3 = ces_4_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_4_31_clock = clock;
  assign ces_4_31_io_ins_0 = ces_3_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_31_io_ins_1 = io_insVertical_0_4; // @[MockArray.scala 45:87]
  assign ces_4_31_io_ins_2 = ces_5_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_31_io_ins_3 = ces_4_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_0_clock = clock;
  assign ces_5_0_io_ins_0 = ces_4_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_0_io_ins_1 = ces_5_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_0_io_ins_2 = ces_6_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_0_io_ins_3 = io_insVertical_1_5; // @[MockArray.scala 47:87]
  assign ces_5_1_clock = clock;
  assign ces_5_1_io_ins_0 = ces_4_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_1_io_ins_1 = ces_5_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_1_io_ins_2 = ces_6_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_1_io_ins_3 = ces_5_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_2_clock = clock;
  assign ces_5_2_io_ins_0 = ces_4_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_2_io_ins_1 = ces_5_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_2_io_ins_2 = ces_6_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_2_io_ins_3 = ces_5_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_3_clock = clock;
  assign ces_5_3_io_ins_0 = ces_4_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_3_io_ins_1 = ces_5_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_3_io_ins_2 = ces_6_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_3_io_ins_3 = ces_5_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_4_clock = clock;
  assign ces_5_4_io_ins_0 = ces_4_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_4_io_ins_1 = ces_5_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_4_io_ins_2 = ces_6_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_4_io_ins_3 = ces_5_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_5_clock = clock;
  assign ces_5_5_io_ins_0 = ces_4_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_5_io_ins_1 = ces_5_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_5_io_ins_2 = ces_6_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_5_io_ins_3 = ces_5_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_6_clock = clock;
  assign ces_5_6_io_ins_0 = ces_4_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_6_io_ins_1 = ces_5_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_6_io_ins_2 = ces_6_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_6_io_ins_3 = ces_5_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_7_clock = clock;
  assign ces_5_7_io_ins_0 = ces_4_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_7_io_ins_1 = ces_5_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_7_io_ins_2 = ces_6_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_7_io_ins_3 = ces_5_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_8_clock = clock;
  assign ces_5_8_io_ins_0 = ces_4_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_8_io_ins_1 = ces_5_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_8_io_ins_2 = ces_6_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_8_io_ins_3 = ces_5_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_9_clock = clock;
  assign ces_5_9_io_ins_0 = ces_4_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_9_io_ins_1 = ces_5_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_9_io_ins_2 = ces_6_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_9_io_ins_3 = ces_5_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_10_clock = clock;
  assign ces_5_10_io_ins_0 = ces_4_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_10_io_ins_1 = ces_5_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_10_io_ins_2 = ces_6_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_10_io_ins_3 = ces_5_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_11_clock = clock;
  assign ces_5_11_io_ins_0 = ces_4_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_11_io_ins_1 = ces_5_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_11_io_ins_2 = ces_6_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_11_io_ins_3 = ces_5_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_12_clock = clock;
  assign ces_5_12_io_ins_0 = ces_4_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_12_io_ins_1 = ces_5_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_12_io_ins_2 = ces_6_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_12_io_ins_3 = ces_5_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_13_clock = clock;
  assign ces_5_13_io_ins_0 = ces_4_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_13_io_ins_1 = ces_5_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_13_io_ins_2 = ces_6_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_13_io_ins_3 = ces_5_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_14_clock = clock;
  assign ces_5_14_io_ins_0 = ces_4_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_14_io_ins_1 = ces_5_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_14_io_ins_2 = ces_6_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_14_io_ins_3 = ces_5_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_15_clock = clock;
  assign ces_5_15_io_ins_0 = ces_4_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_15_io_ins_1 = ces_5_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_15_io_ins_2 = ces_6_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_15_io_ins_3 = ces_5_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_16_clock = clock;
  assign ces_5_16_io_ins_0 = ces_4_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_16_io_ins_1 = ces_5_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_16_io_ins_2 = ces_6_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_16_io_ins_3 = ces_5_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_17_clock = clock;
  assign ces_5_17_io_ins_0 = ces_4_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_17_io_ins_1 = ces_5_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_17_io_ins_2 = ces_6_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_17_io_ins_3 = ces_5_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_18_clock = clock;
  assign ces_5_18_io_ins_0 = ces_4_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_18_io_ins_1 = ces_5_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_18_io_ins_2 = ces_6_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_18_io_ins_3 = ces_5_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_19_clock = clock;
  assign ces_5_19_io_ins_0 = ces_4_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_19_io_ins_1 = ces_5_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_19_io_ins_2 = ces_6_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_19_io_ins_3 = ces_5_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_20_clock = clock;
  assign ces_5_20_io_ins_0 = ces_4_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_20_io_ins_1 = ces_5_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_20_io_ins_2 = ces_6_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_20_io_ins_3 = ces_5_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_21_clock = clock;
  assign ces_5_21_io_ins_0 = ces_4_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_21_io_ins_1 = ces_5_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_21_io_ins_2 = ces_6_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_21_io_ins_3 = ces_5_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_22_clock = clock;
  assign ces_5_22_io_ins_0 = ces_4_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_22_io_ins_1 = ces_5_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_22_io_ins_2 = ces_6_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_22_io_ins_3 = ces_5_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_23_clock = clock;
  assign ces_5_23_io_ins_0 = ces_4_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_23_io_ins_1 = ces_5_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_23_io_ins_2 = ces_6_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_23_io_ins_3 = ces_5_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_24_clock = clock;
  assign ces_5_24_io_ins_0 = ces_4_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_24_io_ins_1 = ces_5_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_24_io_ins_2 = ces_6_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_24_io_ins_3 = ces_5_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_25_clock = clock;
  assign ces_5_25_io_ins_0 = ces_4_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_25_io_ins_1 = ces_5_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_25_io_ins_2 = ces_6_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_25_io_ins_3 = ces_5_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_26_clock = clock;
  assign ces_5_26_io_ins_0 = ces_4_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_26_io_ins_1 = ces_5_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_26_io_ins_2 = ces_6_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_26_io_ins_3 = ces_5_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_27_clock = clock;
  assign ces_5_27_io_ins_0 = ces_4_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_27_io_ins_1 = ces_5_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_27_io_ins_2 = ces_6_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_27_io_ins_3 = ces_5_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_28_clock = clock;
  assign ces_5_28_io_ins_0 = ces_4_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_28_io_ins_1 = ces_5_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_28_io_ins_2 = ces_6_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_28_io_ins_3 = ces_5_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_29_clock = clock;
  assign ces_5_29_io_ins_0 = ces_4_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_29_io_ins_1 = ces_5_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_29_io_ins_2 = ces_6_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_29_io_ins_3 = ces_5_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_30_clock = clock;
  assign ces_5_30_io_ins_0 = ces_4_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_30_io_ins_1 = ces_5_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_5_30_io_ins_2 = ces_6_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_30_io_ins_3 = ces_5_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_5_31_clock = clock;
  assign ces_5_31_io_ins_0 = ces_4_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_31_io_ins_1 = io_insVertical_0_5; // @[MockArray.scala 45:87]
  assign ces_5_31_io_ins_2 = ces_6_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_31_io_ins_3 = ces_5_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_0_clock = clock;
  assign ces_6_0_io_ins_0 = ces_5_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_0_io_ins_1 = ces_6_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_0_io_ins_2 = ces_7_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_0_io_ins_3 = io_insVertical_1_6; // @[MockArray.scala 47:87]
  assign ces_6_1_clock = clock;
  assign ces_6_1_io_ins_0 = ces_5_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_1_io_ins_1 = ces_6_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_1_io_ins_2 = ces_7_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_1_io_ins_3 = ces_6_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_2_clock = clock;
  assign ces_6_2_io_ins_0 = ces_5_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_2_io_ins_1 = ces_6_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_2_io_ins_2 = ces_7_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_2_io_ins_3 = ces_6_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_3_clock = clock;
  assign ces_6_3_io_ins_0 = ces_5_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_3_io_ins_1 = ces_6_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_3_io_ins_2 = ces_7_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_3_io_ins_3 = ces_6_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_4_clock = clock;
  assign ces_6_4_io_ins_0 = ces_5_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_4_io_ins_1 = ces_6_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_4_io_ins_2 = ces_7_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_4_io_ins_3 = ces_6_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_5_clock = clock;
  assign ces_6_5_io_ins_0 = ces_5_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_5_io_ins_1 = ces_6_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_5_io_ins_2 = ces_7_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_5_io_ins_3 = ces_6_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_6_clock = clock;
  assign ces_6_6_io_ins_0 = ces_5_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_6_io_ins_1 = ces_6_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_6_io_ins_2 = ces_7_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_6_io_ins_3 = ces_6_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_7_clock = clock;
  assign ces_6_7_io_ins_0 = ces_5_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_7_io_ins_1 = ces_6_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_7_io_ins_2 = ces_7_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_7_io_ins_3 = ces_6_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_8_clock = clock;
  assign ces_6_8_io_ins_0 = ces_5_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_8_io_ins_1 = ces_6_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_8_io_ins_2 = ces_7_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_8_io_ins_3 = ces_6_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_9_clock = clock;
  assign ces_6_9_io_ins_0 = ces_5_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_9_io_ins_1 = ces_6_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_9_io_ins_2 = ces_7_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_9_io_ins_3 = ces_6_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_10_clock = clock;
  assign ces_6_10_io_ins_0 = ces_5_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_10_io_ins_1 = ces_6_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_10_io_ins_2 = ces_7_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_10_io_ins_3 = ces_6_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_11_clock = clock;
  assign ces_6_11_io_ins_0 = ces_5_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_11_io_ins_1 = ces_6_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_11_io_ins_2 = ces_7_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_11_io_ins_3 = ces_6_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_12_clock = clock;
  assign ces_6_12_io_ins_0 = ces_5_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_12_io_ins_1 = ces_6_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_12_io_ins_2 = ces_7_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_12_io_ins_3 = ces_6_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_13_clock = clock;
  assign ces_6_13_io_ins_0 = ces_5_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_13_io_ins_1 = ces_6_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_13_io_ins_2 = ces_7_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_13_io_ins_3 = ces_6_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_14_clock = clock;
  assign ces_6_14_io_ins_0 = ces_5_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_14_io_ins_1 = ces_6_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_14_io_ins_2 = ces_7_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_14_io_ins_3 = ces_6_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_15_clock = clock;
  assign ces_6_15_io_ins_0 = ces_5_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_15_io_ins_1 = ces_6_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_15_io_ins_2 = ces_7_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_15_io_ins_3 = ces_6_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_16_clock = clock;
  assign ces_6_16_io_ins_0 = ces_5_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_16_io_ins_1 = ces_6_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_16_io_ins_2 = ces_7_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_16_io_ins_3 = ces_6_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_17_clock = clock;
  assign ces_6_17_io_ins_0 = ces_5_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_17_io_ins_1 = ces_6_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_17_io_ins_2 = ces_7_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_17_io_ins_3 = ces_6_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_18_clock = clock;
  assign ces_6_18_io_ins_0 = ces_5_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_18_io_ins_1 = ces_6_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_18_io_ins_2 = ces_7_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_18_io_ins_3 = ces_6_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_19_clock = clock;
  assign ces_6_19_io_ins_0 = ces_5_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_19_io_ins_1 = ces_6_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_19_io_ins_2 = ces_7_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_19_io_ins_3 = ces_6_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_20_clock = clock;
  assign ces_6_20_io_ins_0 = ces_5_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_20_io_ins_1 = ces_6_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_20_io_ins_2 = ces_7_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_20_io_ins_3 = ces_6_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_21_clock = clock;
  assign ces_6_21_io_ins_0 = ces_5_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_21_io_ins_1 = ces_6_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_21_io_ins_2 = ces_7_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_21_io_ins_3 = ces_6_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_22_clock = clock;
  assign ces_6_22_io_ins_0 = ces_5_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_22_io_ins_1 = ces_6_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_22_io_ins_2 = ces_7_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_22_io_ins_3 = ces_6_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_23_clock = clock;
  assign ces_6_23_io_ins_0 = ces_5_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_23_io_ins_1 = ces_6_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_23_io_ins_2 = ces_7_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_23_io_ins_3 = ces_6_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_24_clock = clock;
  assign ces_6_24_io_ins_0 = ces_5_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_24_io_ins_1 = ces_6_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_24_io_ins_2 = ces_7_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_24_io_ins_3 = ces_6_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_25_clock = clock;
  assign ces_6_25_io_ins_0 = ces_5_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_25_io_ins_1 = ces_6_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_25_io_ins_2 = ces_7_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_25_io_ins_3 = ces_6_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_26_clock = clock;
  assign ces_6_26_io_ins_0 = ces_5_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_26_io_ins_1 = ces_6_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_26_io_ins_2 = ces_7_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_26_io_ins_3 = ces_6_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_27_clock = clock;
  assign ces_6_27_io_ins_0 = ces_5_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_27_io_ins_1 = ces_6_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_27_io_ins_2 = ces_7_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_27_io_ins_3 = ces_6_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_28_clock = clock;
  assign ces_6_28_io_ins_0 = ces_5_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_28_io_ins_1 = ces_6_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_28_io_ins_2 = ces_7_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_28_io_ins_3 = ces_6_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_29_clock = clock;
  assign ces_6_29_io_ins_0 = ces_5_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_29_io_ins_1 = ces_6_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_29_io_ins_2 = ces_7_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_29_io_ins_3 = ces_6_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_30_clock = clock;
  assign ces_6_30_io_ins_0 = ces_5_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_30_io_ins_1 = ces_6_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_6_30_io_ins_2 = ces_7_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_30_io_ins_3 = ces_6_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_6_31_clock = clock;
  assign ces_6_31_io_ins_0 = ces_5_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_31_io_ins_1 = io_insVertical_0_6; // @[MockArray.scala 45:87]
  assign ces_6_31_io_ins_2 = ces_7_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_31_io_ins_3 = ces_6_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_0_clock = clock;
  assign ces_7_0_io_ins_0 = ces_6_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_0_io_ins_1 = ces_7_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_0_io_ins_2 = ces_8_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_0_io_ins_3 = io_insVertical_1_7; // @[MockArray.scala 47:87]
  assign ces_7_1_clock = clock;
  assign ces_7_1_io_ins_0 = ces_6_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_1_io_ins_1 = ces_7_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_1_io_ins_2 = ces_8_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_1_io_ins_3 = ces_7_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_2_clock = clock;
  assign ces_7_2_io_ins_0 = ces_6_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_2_io_ins_1 = ces_7_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_2_io_ins_2 = ces_8_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_2_io_ins_3 = ces_7_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_3_clock = clock;
  assign ces_7_3_io_ins_0 = ces_6_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_3_io_ins_1 = ces_7_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_3_io_ins_2 = ces_8_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_3_io_ins_3 = ces_7_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_4_clock = clock;
  assign ces_7_4_io_ins_0 = ces_6_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_4_io_ins_1 = ces_7_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_4_io_ins_2 = ces_8_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_4_io_ins_3 = ces_7_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_5_clock = clock;
  assign ces_7_5_io_ins_0 = ces_6_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_5_io_ins_1 = ces_7_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_5_io_ins_2 = ces_8_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_5_io_ins_3 = ces_7_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_6_clock = clock;
  assign ces_7_6_io_ins_0 = ces_6_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_6_io_ins_1 = ces_7_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_6_io_ins_2 = ces_8_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_6_io_ins_3 = ces_7_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_7_clock = clock;
  assign ces_7_7_io_ins_0 = ces_6_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_7_io_ins_1 = ces_7_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_7_io_ins_2 = ces_8_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_7_io_ins_3 = ces_7_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_8_clock = clock;
  assign ces_7_8_io_ins_0 = ces_6_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_8_io_ins_1 = ces_7_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_8_io_ins_2 = ces_8_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_8_io_ins_3 = ces_7_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_9_clock = clock;
  assign ces_7_9_io_ins_0 = ces_6_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_9_io_ins_1 = ces_7_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_9_io_ins_2 = ces_8_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_9_io_ins_3 = ces_7_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_10_clock = clock;
  assign ces_7_10_io_ins_0 = ces_6_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_10_io_ins_1 = ces_7_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_10_io_ins_2 = ces_8_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_10_io_ins_3 = ces_7_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_11_clock = clock;
  assign ces_7_11_io_ins_0 = ces_6_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_11_io_ins_1 = ces_7_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_11_io_ins_2 = ces_8_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_11_io_ins_3 = ces_7_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_12_clock = clock;
  assign ces_7_12_io_ins_0 = ces_6_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_12_io_ins_1 = ces_7_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_12_io_ins_2 = ces_8_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_12_io_ins_3 = ces_7_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_13_clock = clock;
  assign ces_7_13_io_ins_0 = ces_6_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_13_io_ins_1 = ces_7_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_13_io_ins_2 = ces_8_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_13_io_ins_3 = ces_7_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_14_clock = clock;
  assign ces_7_14_io_ins_0 = ces_6_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_14_io_ins_1 = ces_7_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_14_io_ins_2 = ces_8_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_14_io_ins_3 = ces_7_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_15_clock = clock;
  assign ces_7_15_io_ins_0 = ces_6_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_15_io_ins_1 = ces_7_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_15_io_ins_2 = ces_8_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_15_io_ins_3 = ces_7_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_16_clock = clock;
  assign ces_7_16_io_ins_0 = ces_6_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_16_io_ins_1 = ces_7_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_16_io_ins_2 = ces_8_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_16_io_ins_3 = ces_7_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_17_clock = clock;
  assign ces_7_17_io_ins_0 = ces_6_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_17_io_ins_1 = ces_7_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_17_io_ins_2 = ces_8_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_17_io_ins_3 = ces_7_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_18_clock = clock;
  assign ces_7_18_io_ins_0 = ces_6_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_18_io_ins_1 = ces_7_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_18_io_ins_2 = ces_8_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_18_io_ins_3 = ces_7_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_19_clock = clock;
  assign ces_7_19_io_ins_0 = ces_6_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_19_io_ins_1 = ces_7_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_19_io_ins_2 = ces_8_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_19_io_ins_3 = ces_7_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_20_clock = clock;
  assign ces_7_20_io_ins_0 = ces_6_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_20_io_ins_1 = ces_7_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_20_io_ins_2 = ces_8_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_20_io_ins_3 = ces_7_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_21_clock = clock;
  assign ces_7_21_io_ins_0 = ces_6_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_21_io_ins_1 = ces_7_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_21_io_ins_2 = ces_8_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_21_io_ins_3 = ces_7_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_22_clock = clock;
  assign ces_7_22_io_ins_0 = ces_6_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_22_io_ins_1 = ces_7_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_22_io_ins_2 = ces_8_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_22_io_ins_3 = ces_7_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_23_clock = clock;
  assign ces_7_23_io_ins_0 = ces_6_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_23_io_ins_1 = ces_7_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_23_io_ins_2 = ces_8_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_23_io_ins_3 = ces_7_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_24_clock = clock;
  assign ces_7_24_io_ins_0 = ces_6_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_24_io_ins_1 = ces_7_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_24_io_ins_2 = ces_8_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_24_io_ins_3 = ces_7_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_25_clock = clock;
  assign ces_7_25_io_ins_0 = ces_6_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_25_io_ins_1 = ces_7_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_25_io_ins_2 = ces_8_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_25_io_ins_3 = ces_7_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_26_clock = clock;
  assign ces_7_26_io_ins_0 = ces_6_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_26_io_ins_1 = ces_7_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_26_io_ins_2 = ces_8_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_26_io_ins_3 = ces_7_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_27_clock = clock;
  assign ces_7_27_io_ins_0 = ces_6_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_27_io_ins_1 = ces_7_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_27_io_ins_2 = ces_8_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_27_io_ins_3 = ces_7_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_28_clock = clock;
  assign ces_7_28_io_ins_0 = ces_6_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_28_io_ins_1 = ces_7_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_28_io_ins_2 = ces_8_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_28_io_ins_3 = ces_7_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_29_clock = clock;
  assign ces_7_29_io_ins_0 = ces_6_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_29_io_ins_1 = ces_7_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_29_io_ins_2 = ces_8_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_29_io_ins_3 = ces_7_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_30_clock = clock;
  assign ces_7_30_io_ins_0 = ces_6_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_30_io_ins_1 = ces_7_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_7_30_io_ins_2 = ces_8_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_30_io_ins_3 = ces_7_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_7_31_clock = clock;
  assign ces_7_31_io_ins_0 = ces_6_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_31_io_ins_1 = io_insVertical_0_7; // @[MockArray.scala 45:87]
  assign ces_7_31_io_ins_2 = ces_8_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_31_io_ins_3 = ces_7_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_0_clock = clock;
  assign ces_8_0_io_ins_0 = ces_7_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_0_io_ins_1 = ces_8_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_0_io_ins_2 = ces_9_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_0_io_ins_3 = io_insVertical_1_8; // @[MockArray.scala 47:87]
  assign ces_8_1_clock = clock;
  assign ces_8_1_io_ins_0 = ces_7_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_1_io_ins_1 = ces_8_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_1_io_ins_2 = ces_9_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_1_io_ins_3 = ces_8_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_2_clock = clock;
  assign ces_8_2_io_ins_0 = ces_7_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_2_io_ins_1 = ces_8_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_2_io_ins_2 = ces_9_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_2_io_ins_3 = ces_8_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_3_clock = clock;
  assign ces_8_3_io_ins_0 = ces_7_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_3_io_ins_1 = ces_8_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_3_io_ins_2 = ces_9_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_3_io_ins_3 = ces_8_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_4_clock = clock;
  assign ces_8_4_io_ins_0 = ces_7_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_4_io_ins_1 = ces_8_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_4_io_ins_2 = ces_9_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_4_io_ins_3 = ces_8_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_5_clock = clock;
  assign ces_8_5_io_ins_0 = ces_7_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_5_io_ins_1 = ces_8_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_5_io_ins_2 = ces_9_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_5_io_ins_3 = ces_8_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_6_clock = clock;
  assign ces_8_6_io_ins_0 = ces_7_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_6_io_ins_1 = ces_8_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_6_io_ins_2 = ces_9_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_6_io_ins_3 = ces_8_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_7_clock = clock;
  assign ces_8_7_io_ins_0 = ces_7_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_7_io_ins_1 = ces_8_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_7_io_ins_2 = ces_9_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_7_io_ins_3 = ces_8_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_8_clock = clock;
  assign ces_8_8_io_ins_0 = ces_7_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_8_io_ins_1 = ces_8_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_8_io_ins_2 = ces_9_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_8_io_ins_3 = ces_8_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_9_clock = clock;
  assign ces_8_9_io_ins_0 = ces_7_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_9_io_ins_1 = ces_8_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_9_io_ins_2 = ces_9_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_9_io_ins_3 = ces_8_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_10_clock = clock;
  assign ces_8_10_io_ins_0 = ces_7_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_10_io_ins_1 = ces_8_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_10_io_ins_2 = ces_9_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_10_io_ins_3 = ces_8_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_11_clock = clock;
  assign ces_8_11_io_ins_0 = ces_7_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_11_io_ins_1 = ces_8_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_11_io_ins_2 = ces_9_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_11_io_ins_3 = ces_8_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_12_clock = clock;
  assign ces_8_12_io_ins_0 = ces_7_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_12_io_ins_1 = ces_8_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_12_io_ins_2 = ces_9_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_12_io_ins_3 = ces_8_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_13_clock = clock;
  assign ces_8_13_io_ins_0 = ces_7_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_13_io_ins_1 = ces_8_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_13_io_ins_2 = ces_9_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_13_io_ins_3 = ces_8_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_14_clock = clock;
  assign ces_8_14_io_ins_0 = ces_7_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_14_io_ins_1 = ces_8_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_14_io_ins_2 = ces_9_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_14_io_ins_3 = ces_8_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_15_clock = clock;
  assign ces_8_15_io_ins_0 = ces_7_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_15_io_ins_1 = ces_8_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_15_io_ins_2 = ces_9_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_15_io_ins_3 = ces_8_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_16_clock = clock;
  assign ces_8_16_io_ins_0 = ces_7_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_16_io_ins_1 = ces_8_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_16_io_ins_2 = ces_9_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_16_io_ins_3 = ces_8_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_17_clock = clock;
  assign ces_8_17_io_ins_0 = ces_7_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_17_io_ins_1 = ces_8_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_17_io_ins_2 = ces_9_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_17_io_ins_3 = ces_8_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_18_clock = clock;
  assign ces_8_18_io_ins_0 = ces_7_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_18_io_ins_1 = ces_8_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_18_io_ins_2 = ces_9_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_18_io_ins_3 = ces_8_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_19_clock = clock;
  assign ces_8_19_io_ins_0 = ces_7_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_19_io_ins_1 = ces_8_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_19_io_ins_2 = ces_9_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_19_io_ins_3 = ces_8_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_20_clock = clock;
  assign ces_8_20_io_ins_0 = ces_7_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_20_io_ins_1 = ces_8_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_20_io_ins_2 = ces_9_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_20_io_ins_3 = ces_8_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_21_clock = clock;
  assign ces_8_21_io_ins_0 = ces_7_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_21_io_ins_1 = ces_8_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_21_io_ins_2 = ces_9_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_21_io_ins_3 = ces_8_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_22_clock = clock;
  assign ces_8_22_io_ins_0 = ces_7_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_22_io_ins_1 = ces_8_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_22_io_ins_2 = ces_9_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_22_io_ins_3 = ces_8_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_23_clock = clock;
  assign ces_8_23_io_ins_0 = ces_7_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_23_io_ins_1 = ces_8_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_23_io_ins_2 = ces_9_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_23_io_ins_3 = ces_8_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_24_clock = clock;
  assign ces_8_24_io_ins_0 = ces_7_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_24_io_ins_1 = ces_8_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_24_io_ins_2 = ces_9_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_24_io_ins_3 = ces_8_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_25_clock = clock;
  assign ces_8_25_io_ins_0 = ces_7_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_25_io_ins_1 = ces_8_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_25_io_ins_2 = ces_9_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_25_io_ins_3 = ces_8_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_26_clock = clock;
  assign ces_8_26_io_ins_0 = ces_7_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_26_io_ins_1 = ces_8_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_26_io_ins_2 = ces_9_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_26_io_ins_3 = ces_8_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_27_clock = clock;
  assign ces_8_27_io_ins_0 = ces_7_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_27_io_ins_1 = ces_8_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_27_io_ins_2 = ces_9_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_27_io_ins_3 = ces_8_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_28_clock = clock;
  assign ces_8_28_io_ins_0 = ces_7_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_28_io_ins_1 = ces_8_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_28_io_ins_2 = ces_9_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_28_io_ins_3 = ces_8_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_29_clock = clock;
  assign ces_8_29_io_ins_0 = ces_7_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_29_io_ins_1 = ces_8_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_29_io_ins_2 = ces_9_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_29_io_ins_3 = ces_8_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_30_clock = clock;
  assign ces_8_30_io_ins_0 = ces_7_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_30_io_ins_1 = ces_8_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_8_30_io_ins_2 = ces_9_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_30_io_ins_3 = ces_8_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_8_31_clock = clock;
  assign ces_8_31_io_ins_0 = ces_7_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_31_io_ins_1 = io_insVertical_0_8; // @[MockArray.scala 45:87]
  assign ces_8_31_io_ins_2 = ces_9_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_31_io_ins_3 = ces_8_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_0_clock = clock;
  assign ces_9_0_io_ins_0 = ces_8_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_0_io_ins_1 = ces_9_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_0_io_ins_2 = ces_10_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_0_io_ins_3 = io_insVertical_1_9; // @[MockArray.scala 47:87]
  assign ces_9_1_clock = clock;
  assign ces_9_1_io_ins_0 = ces_8_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_1_io_ins_1 = ces_9_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_1_io_ins_2 = ces_10_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_1_io_ins_3 = ces_9_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_2_clock = clock;
  assign ces_9_2_io_ins_0 = ces_8_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_2_io_ins_1 = ces_9_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_2_io_ins_2 = ces_10_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_2_io_ins_3 = ces_9_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_3_clock = clock;
  assign ces_9_3_io_ins_0 = ces_8_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_3_io_ins_1 = ces_9_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_3_io_ins_2 = ces_10_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_3_io_ins_3 = ces_9_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_4_clock = clock;
  assign ces_9_4_io_ins_0 = ces_8_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_4_io_ins_1 = ces_9_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_4_io_ins_2 = ces_10_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_4_io_ins_3 = ces_9_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_5_clock = clock;
  assign ces_9_5_io_ins_0 = ces_8_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_5_io_ins_1 = ces_9_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_5_io_ins_2 = ces_10_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_5_io_ins_3 = ces_9_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_6_clock = clock;
  assign ces_9_6_io_ins_0 = ces_8_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_6_io_ins_1 = ces_9_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_6_io_ins_2 = ces_10_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_6_io_ins_3 = ces_9_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_7_clock = clock;
  assign ces_9_7_io_ins_0 = ces_8_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_7_io_ins_1 = ces_9_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_7_io_ins_2 = ces_10_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_7_io_ins_3 = ces_9_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_8_clock = clock;
  assign ces_9_8_io_ins_0 = ces_8_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_8_io_ins_1 = ces_9_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_8_io_ins_2 = ces_10_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_8_io_ins_3 = ces_9_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_9_clock = clock;
  assign ces_9_9_io_ins_0 = ces_8_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_9_io_ins_1 = ces_9_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_9_io_ins_2 = ces_10_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_9_io_ins_3 = ces_9_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_10_clock = clock;
  assign ces_9_10_io_ins_0 = ces_8_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_10_io_ins_1 = ces_9_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_10_io_ins_2 = ces_10_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_10_io_ins_3 = ces_9_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_11_clock = clock;
  assign ces_9_11_io_ins_0 = ces_8_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_11_io_ins_1 = ces_9_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_11_io_ins_2 = ces_10_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_11_io_ins_3 = ces_9_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_12_clock = clock;
  assign ces_9_12_io_ins_0 = ces_8_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_12_io_ins_1 = ces_9_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_12_io_ins_2 = ces_10_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_12_io_ins_3 = ces_9_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_13_clock = clock;
  assign ces_9_13_io_ins_0 = ces_8_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_13_io_ins_1 = ces_9_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_13_io_ins_2 = ces_10_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_13_io_ins_3 = ces_9_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_14_clock = clock;
  assign ces_9_14_io_ins_0 = ces_8_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_14_io_ins_1 = ces_9_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_14_io_ins_2 = ces_10_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_14_io_ins_3 = ces_9_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_15_clock = clock;
  assign ces_9_15_io_ins_0 = ces_8_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_15_io_ins_1 = ces_9_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_15_io_ins_2 = ces_10_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_15_io_ins_3 = ces_9_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_16_clock = clock;
  assign ces_9_16_io_ins_0 = ces_8_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_16_io_ins_1 = ces_9_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_16_io_ins_2 = ces_10_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_16_io_ins_3 = ces_9_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_17_clock = clock;
  assign ces_9_17_io_ins_0 = ces_8_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_17_io_ins_1 = ces_9_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_17_io_ins_2 = ces_10_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_17_io_ins_3 = ces_9_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_18_clock = clock;
  assign ces_9_18_io_ins_0 = ces_8_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_18_io_ins_1 = ces_9_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_18_io_ins_2 = ces_10_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_18_io_ins_3 = ces_9_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_19_clock = clock;
  assign ces_9_19_io_ins_0 = ces_8_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_19_io_ins_1 = ces_9_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_19_io_ins_2 = ces_10_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_19_io_ins_3 = ces_9_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_20_clock = clock;
  assign ces_9_20_io_ins_0 = ces_8_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_20_io_ins_1 = ces_9_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_20_io_ins_2 = ces_10_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_20_io_ins_3 = ces_9_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_21_clock = clock;
  assign ces_9_21_io_ins_0 = ces_8_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_21_io_ins_1 = ces_9_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_21_io_ins_2 = ces_10_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_21_io_ins_3 = ces_9_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_22_clock = clock;
  assign ces_9_22_io_ins_0 = ces_8_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_22_io_ins_1 = ces_9_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_22_io_ins_2 = ces_10_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_22_io_ins_3 = ces_9_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_23_clock = clock;
  assign ces_9_23_io_ins_0 = ces_8_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_23_io_ins_1 = ces_9_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_23_io_ins_2 = ces_10_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_23_io_ins_3 = ces_9_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_24_clock = clock;
  assign ces_9_24_io_ins_0 = ces_8_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_24_io_ins_1 = ces_9_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_24_io_ins_2 = ces_10_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_24_io_ins_3 = ces_9_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_25_clock = clock;
  assign ces_9_25_io_ins_0 = ces_8_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_25_io_ins_1 = ces_9_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_25_io_ins_2 = ces_10_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_25_io_ins_3 = ces_9_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_26_clock = clock;
  assign ces_9_26_io_ins_0 = ces_8_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_26_io_ins_1 = ces_9_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_26_io_ins_2 = ces_10_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_26_io_ins_3 = ces_9_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_27_clock = clock;
  assign ces_9_27_io_ins_0 = ces_8_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_27_io_ins_1 = ces_9_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_27_io_ins_2 = ces_10_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_27_io_ins_3 = ces_9_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_28_clock = clock;
  assign ces_9_28_io_ins_0 = ces_8_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_28_io_ins_1 = ces_9_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_28_io_ins_2 = ces_10_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_28_io_ins_3 = ces_9_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_29_clock = clock;
  assign ces_9_29_io_ins_0 = ces_8_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_29_io_ins_1 = ces_9_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_29_io_ins_2 = ces_10_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_29_io_ins_3 = ces_9_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_30_clock = clock;
  assign ces_9_30_io_ins_0 = ces_8_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_30_io_ins_1 = ces_9_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_9_30_io_ins_2 = ces_10_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_30_io_ins_3 = ces_9_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_9_31_clock = clock;
  assign ces_9_31_io_ins_0 = ces_8_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_31_io_ins_1 = io_insVertical_0_9; // @[MockArray.scala 45:87]
  assign ces_9_31_io_ins_2 = ces_10_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_31_io_ins_3 = ces_9_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_0_clock = clock;
  assign ces_10_0_io_ins_0 = ces_9_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_0_io_ins_1 = ces_10_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_0_io_ins_2 = ces_11_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_0_io_ins_3 = io_insVertical_1_10; // @[MockArray.scala 47:87]
  assign ces_10_1_clock = clock;
  assign ces_10_1_io_ins_0 = ces_9_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_1_io_ins_1 = ces_10_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_1_io_ins_2 = ces_11_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_1_io_ins_3 = ces_10_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_2_clock = clock;
  assign ces_10_2_io_ins_0 = ces_9_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_2_io_ins_1 = ces_10_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_2_io_ins_2 = ces_11_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_2_io_ins_3 = ces_10_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_3_clock = clock;
  assign ces_10_3_io_ins_0 = ces_9_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_3_io_ins_1 = ces_10_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_3_io_ins_2 = ces_11_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_3_io_ins_3 = ces_10_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_4_clock = clock;
  assign ces_10_4_io_ins_0 = ces_9_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_4_io_ins_1 = ces_10_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_4_io_ins_2 = ces_11_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_4_io_ins_3 = ces_10_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_5_clock = clock;
  assign ces_10_5_io_ins_0 = ces_9_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_5_io_ins_1 = ces_10_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_5_io_ins_2 = ces_11_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_5_io_ins_3 = ces_10_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_6_clock = clock;
  assign ces_10_6_io_ins_0 = ces_9_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_6_io_ins_1 = ces_10_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_6_io_ins_2 = ces_11_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_6_io_ins_3 = ces_10_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_7_clock = clock;
  assign ces_10_7_io_ins_0 = ces_9_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_7_io_ins_1 = ces_10_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_7_io_ins_2 = ces_11_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_7_io_ins_3 = ces_10_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_8_clock = clock;
  assign ces_10_8_io_ins_0 = ces_9_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_8_io_ins_1 = ces_10_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_8_io_ins_2 = ces_11_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_8_io_ins_3 = ces_10_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_9_clock = clock;
  assign ces_10_9_io_ins_0 = ces_9_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_9_io_ins_1 = ces_10_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_9_io_ins_2 = ces_11_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_9_io_ins_3 = ces_10_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_10_clock = clock;
  assign ces_10_10_io_ins_0 = ces_9_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_10_io_ins_1 = ces_10_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_10_io_ins_2 = ces_11_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_10_io_ins_3 = ces_10_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_11_clock = clock;
  assign ces_10_11_io_ins_0 = ces_9_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_11_io_ins_1 = ces_10_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_11_io_ins_2 = ces_11_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_11_io_ins_3 = ces_10_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_12_clock = clock;
  assign ces_10_12_io_ins_0 = ces_9_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_12_io_ins_1 = ces_10_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_12_io_ins_2 = ces_11_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_12_io_ins_3 = ces_10_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_13_clock = clock;
  assign ces_10_13_io_ins_0 = ces_9_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_13_io_ins_1 = ces_10_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_13_io_ins_2 = ces_11_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_13_io_ins_3 = ces_10_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_14_clock = clock;
  assign ces_10_14_io_ins_0 = ces_9_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_14_io_ins_1 = ces_10_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_14_io_ins_2 = ces_11_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_14_io_ins_3 = ces_10_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_15_clock = clock;
  assign ces_10_15_io_ins_0 = ces_9_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_15_io_ins_1 = ces_10_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_15_io_ins_2 = ces_11_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_15_io_ins_3 = ces_10_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_16_clock = clock;
  assign ces_10_16_io_ins_0 = ces_9_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_16_io_ins_1 = ces_10_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_16_io_ins_2 = ces_11_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_16_io_ins_3 = ces_10_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_17_clock = clock;
  assign ces_10_17_io_ins_0 = ces_9_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_17_io_ins_1 = ces_10_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_17_io_ins_2 = ces_11_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_17_io_ins_3 = ces_10_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_18_clock = clock;
  assign ces_10_18_io_ins_0 = ces_9_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_18_io_ins_1 = ces_10_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_18_io_ins_2 = ces_11_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_18_io_ins_3 = ces_10_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_19_clock = clock;
  assign ces_10_19_io_ins_0 = ces_9_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_19_io_ins_1 = ces_10_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_19_io_ins_2 = ces_11_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_19_io_ins_3 = ces_10_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_20_clock = clock;
  assign ces_10_20_io_ins_0 = ces_9_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_20_io_ins_1 = ces_10_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_20_io_ins_2 = ces_11_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_20_io_ins_3 = ces_10_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_21_clock = clock;
  assign ces_10_21_io_ins_0 = ces_9_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_21_io_ins_1 = ces_10_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_21_io_ins_2 = ces_11_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_21_io_ins_3 = ces_10_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_22_clock = clock;
  assign ces_10_22_io_ins_0 = ces_9_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_22_io_ins_1 = ces_10_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_22_io_ins_2 = ces_11_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_22_io_ins_3 = ces_10_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_23_clock = clock;
  assign ces_10_23_io_ins_0 = ces_9_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_23_io_ins_1 = ces_10_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_23_io_ins_2 = ces_11_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_23_io_ins_3 = ces_10_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_24_clock = clock;
  assign ces_10_24_io_ins_0 = ces_9_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_24_io_ins_1 = ces_10_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_24_io_ins_2 = ces_11_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_24_io_ins_3 = ces_10_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_25_clock = clock;
  assign ces_10_25_io_ins_0 = ces_9_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_25_io_ins_1 = ces_10_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_25_io_ins_2 = ces_11_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_25_io_ins_3 = ces_10_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_26_clock = clock;
  assign ces_10_26_io_ins_0 = ces_9_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_26_io_ins_1 = ces_10_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_26_io_ins_2 = ces_11_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_26_io_ins_3 = ces_10_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_27_clock = clock;
  assign ces_10_27_io_ins_0 = ces_9_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_27_io_ins_1 = ces_10_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_27_io_ins_2 = ces_11_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_27_io_ins_3 = ces_10_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_28_clock = clock;
  assign ces_10_28_io_ins_0 = ces_9_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_28_io_ins_1 = ces_10_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_28_io_ins_2 = ces_11_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_28_io_ins_3 = ces_10_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_29_clock = clock;
  assign ces_10_29_io_ins_0 = ces_9_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_29_io_ins_1 = ces_10_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_29_io_ins_2 = ces_11_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_29_io_ins_3 = ces_10_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_30_clock = clock;
  assign ces_10_30_io_ins_0 = ces_9_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_30_io_ins_1 = ces_10_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_10_30_io_ins_2 = ces_11_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_30_io_ins_3 = ces_10_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_10_31_clock = clock;
  assign ces_10_31_io_ins_0 = ces_9_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_31_io_ins_1 = io_insVertical_0_10; // @[MockArray.scala 45:87]
  assign ces_10_31_io_ins_2 = ces_11_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_31_io_ins_3 = ces_10_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_0_clock = clock;
  assign ces_11_0_io_ins_0 = ces_10_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_0_io_ins_1 = ces_11_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_0_io_ins_2 = ces_12_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_0_io_ins_3 = io_insVertical_1_11; // @[MockArray.scala 47:87]
  assign ces_11_1_clock = clock;
  assign ces_11_1_io_ins_0 = ces_10_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_1_io_ins_1 = ces_11_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_1_io_ins_2 = ces_12_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_1_io_ins_3 = ces_11_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_2_clock = clock;
  assign ces_11_2_io_ins_0 = ces_10_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_2_io_ins_1 = ces_11_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_2_io_ins_2 = ces_12_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_2_io_ins_3 = ces_11_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_3_clock = clock;
  assign ces_11_3_io_ins_0 = ces_10_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_3_io_ins_1 = ces_11_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_3_io_ins_2 = ces_12_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_3_io_ins_3 = ces_11_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_4_clock = clock;
  assign ces_11_4_io_ins_0 = ces_10_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_4_io_ins_1 = ces_11_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_4_io_ins_2 = ces_12_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_4_io_ins_3 = ces_11_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_5_clock = clock;
  assign ces_11_5_io_ins_0 = ces_10_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_5_io_ins_1 = ces_11_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_5_io_ins_2 = ces_12_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_5_io_ins_3 = ces_11_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_6_clock = clock;
  assign ces_11_6_io_ins_0 = ces_10_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_6_io_ins_1 = ces_11_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_6_io_ins_2 = ces_12_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_6_io_ins_3 = ces_11_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_7_clock = clock;
  assign ces_11_7_io_ins_0 = ces_10_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_7_io_ins_1 = ces_11_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_7_io_ins_2 = ces_12_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_7_io_ins_3 = ces_11_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_8_clock = clock;
  assign ces_11_8_io_ins_0 = ces_10_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_8_io_ins_1 = ces_11_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_8_io_ins_2 = ces_12_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_8_io_ins_3 = ces_11_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_9_clock = clock;
  assign ces_11_9_io_ins_0 = ces_10_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_9_io_ins_1 = ces_11_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_9_io_ins_2 = ces_12_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_9_io_ins_3 = ces_11_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_10_clock = clock;
  assign ces_11_10_io_ins_0 = ces_10_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_10_io_ins_1 = ces_11_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_10_io_ins_2 = ces_12_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_10_io_ins_3 = ces_11_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_11_clock = clock;
  assign ces_11_11_io_ins_0 = ces_10_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_11_io_ins_1 = ces_11_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_11_io_ins_2 = ces_12_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_11_io_ins_3 = ces_11_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_12_clock = clock;
  assign ces_11_12_io_ins_0 = ces_10_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_12_io_ins_1 = ces_11_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_12_io_ins_2 = ces_12_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_12_io_ins_3 = ces_11_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_13_clock = clock;
  assign ces_11_13_io_ins_0 = ces_10_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_13_io_ins_1 = ces_11_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_13_io_ins_2 = ces_12_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_13_io_ins_3 = ces_11_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_14_clock = clock;
  assign ces_11_14_io_ins_0 = ces_10_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_14_io_ins_1 = ces_11_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_14_io_ins_2 = ces_12_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_14_io_ins_3 = ces_11_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_15_clock = clock;
  assign ces_11_15_io_ins_0 = ces_10_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_15_io_ins_1 = ces_11_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_15_io_ins_2 = ces_12_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_15_io_ins_3 = ces_11_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_16_clock = clock;
  assign ces_11_16_io_ins_0 = ces_10_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_16_io_ins_1 = ces_11_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_16_io_ins_2 = ces_12_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_16_io_ins_3 = ces_11_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_17_clock = clock;
  assign ces_11_17_io_ins_0 = ces_10_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_17_io_ins_1 = ces_11_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_17_io_ins_2 = ces_12_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_17_io_ins_3 = ces_11_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_18_clock = clock;
  assign ces_11_18_io_ins_0 = ces_10_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_18_io_ins_1 = ces_11_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_18_io_ins_2 = ces_12_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_18_io_ins_3 = ces_11_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_19_clock = clock;
  assign ces_11_19_io_ins_0 = ces_10_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_19_io_ins_1 = ces_11_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_19_io_ins_2 = ces_12_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_19_io_ins_3 = ces_11_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_20_clock = clock;
  assign ces_11_20_io_ins_0 = ces_10_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_20_io_ins_1 = ces_11_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_20_io_ins_2 = ces_12_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_20_io_ins_3 = ces_11_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_21_clock = clock;
  assign ces_11_21_io_ins_0 = ces_10_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_21_io_ins_1 = ces_11_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_21_io_ins_2 = ces_12_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_21_io_ins_3 = ces_11_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_22_clock = clock;
  assign ces_11_22_io_ins_0 = ces_10_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_22_io_ins_1 = ces_11_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_22_io_ins_2 = ces_12_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_22_io_ins_3 = ces_11_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_23_clock = clock;
  assign ces_11_23_io_ins_0 = ces_10_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_23_io_ins_1 = ces_11_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_23_io_ins_2 = ces_12_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_23_io_ins_3 = ces_11_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_24_clock = clock;
  assign ces_11_24_io_ins_0 = ces_10_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_24_io_ins_1 = ces_11_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_24_io_ins_2 = ces_12_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_24_io_ins_3 = ces_11_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_25_clock = clock;
  assign ces_11_25_io_ins_0 = ces_10_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_25_io_ins_1 = ces_11_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_25_io_ins_2 = ces_12_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_25_io_ins_3 = ces_11_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_26_clock = clock;
  assign ces_11_26_io_ins_0 = ces_10_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_26_io_ins_1 = ces_11_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_26_io_ins_2 = ces_12_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_26_io_ins_3 = ces_11_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_27_clock = clock;
  assign ces_11_27_io_ins_0 = ces_10_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_27_io_ins_1 = ces_11_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_27_io_ins_2 = ces_12_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_27_io_ins_3 = ces_11_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_28_clock = clock;
  assign ces_11_28_io_ins_0 = ces_10_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_28_io_ins_1 = ces_11_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_28_io_ins_2 = ces_12_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_28_io_ins_3 = ces_11_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_29_clock = clock;
  assign ces_11_29_io_ins_0 = ces_10_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_29_io_ins_1 = ces_11_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_29_io_ins_2 = ces_12_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_29_io_ins_3 = ces_11_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_30_clock = clock;
  assign ces_11_30_io_ins_0 = ces_10_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_30_io_ins_1 = ces_11_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_11_30_io_ins_2 = ces_12_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_30_io_ins_3 = ces_11_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_11_31_clock = clock;
  assign ces_11_31_io_ins_0 = ces_10_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_31_io_ins_1 = io_insVertical_0_11; // @[MockArray.scala 45:87]
  assign ces_11_31_io_ins_2 = ces_12_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_31_io_ins_3 = ces_11_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_0_clock = clock;
  assign ces_12_0_io_ins_0 = ces_11_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_0_io_ins_1 = ces_12_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_0_io_ins_2 = ces_13_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_0_io_ins_3 = io_insVertical_1_12; // @[MockArray.scala 47:87]
  assign ces_12_1_clock = clock;
  assign ces_12_1_io_ins_0 = ces_11_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_1_io_ins_1 = ces_12_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_1_io_ins_2 = ces_13_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_1_io_ins_3 = ces_12_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_2_clock = clock;
  assign ces_12_2_io_ins_0 = ces_11_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_2_io_ins_1 = ces_12_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_2_io_ins_2 = ces_13_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_2_io_ins_3 = ces_12_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_3_clock = clock;
  assign ces_12_3_io_ins_0 = ces_11_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_3_io_ins_1 = ces_12_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_3_io_ins_2 = ces_13_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_3_io_ins_3 = ces_12_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_4_clock = clock;
  assign ces_12_4_io_ins_0 = ces_11_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_4_io_ins_1 = ces_12_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_4_io_ins_2 = ces_13_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_4_io_ins_3 = ces_12_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_5_clock = clock;
  assign ces_12_5_io_ins_0 = ces_11_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_5_io_ins_1 = ces_12_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_5_io_ins_2 = ces_13_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_5_io_ins_3 = ces_12_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_6_clock = clock;
  assign ces_12_6_io_ins_0 = ces_11_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_6_io_ins_1 = ces_12_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_6_io_ins_2 = ces_13_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_6_io_ins_3 = ces_12_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_7_clock = clock;
  assign ces_12_7_io_ins_0 = ces_11_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_7_io_ins_1 = ces_12_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_7_io_ins_2 = ces_13_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_7_io_ins_3 = ces_12_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_8_clock = clock;
  assign ces_12_8_io_ins_0 = ces_11_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_8_io_ins_1 = ces_12_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_8_io_ins_2 = ces_13_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_8_io_ins_3 = ces_12_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_9_clock = clock;
  assign ces_12_9_io_ins_0 = ces_11_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_9_io_ins_1 = ces_12_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_9_io_ins_2 = ces_13_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_9_io_ins_3 = ces_12_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_10_clock = clock;
  assign ces_12_10_io_ins_0 = ces_11_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_10_io_ins_1 = ces_12_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_10_io_ins_2 = ces_13_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_10_io_ins_3 = ces_12_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_11_clock = clock;
  assign ces_12_11_io_ins_0 = ces_11_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_11_io_ins_1 = ces_12_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_11_io_ins_2 = ces_13_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_11_io_ins_3 = ces_12_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_12_clock = clock;
  assign ces_12_12_io_ins_0 = ces_11_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_12_io_ins_1 = ces_12_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_12_io_ins_2 = ces_13_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_12_io_ins_3 = ces_12_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_13_clock = clock;
  assign ces_12_13_io_ins_0 = ces_11_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_13_io_ins_1 = ces_12_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_13_io_ins_2 = ces_13_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_13_io_ins_3 = ces_12_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_14_clock = clock;
  assign ces_12_14_io_ins_0 = ces_11_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_14_io_ins_1 = ces_12_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_14_io_ins_2 = ces_13_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_14_io_ins_3 = ces_12_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_15_clock = clock;
  assign ces_12_15_io_ins_0 = ces_11_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_15_io_ins_1 = ces_12_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_15_io_ins_2 = ces_13_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_15_io_ins_3 = ces_12_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_16_clock = clock;
  assign ces_12_16_io_ins_0 = ces_11_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_16_io_ins_1 = ces_12_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_16_io_ins_2 = ces_13_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_16_io_ins_3 = ces_12_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_17_clock = clock;
  assign ces_12_17_io_ins_0 = ces_11_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_17_io_ins_1 = ces_12_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_17_io_ins_2 = ces_13_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_17_io_ins_3 = ces_12_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_18_clock = clock;
  assign ces_12_18_io_ins_0 = ces_11_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_18_io_ins_1 = ces_12_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_18_io_ins_2 = ces_13_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_18_io_ins_3 = ces_12_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_19_clock = clock;
  assign ces_12_19_io_ins_0 = ces_11_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_19_io_ins_1 = ces_12_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_19_io_ins_2 = ces_13_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_19_io_ins_3 = ces_12_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_20_clock = clock;
  assign ces_12_20_io_ins_0 = ces_11_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_20_io_ins_1 = ces_12_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_20_io_ins_2 = ces_13_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_20_io_ins_3 = ces_12_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_21_clock = clock;
  assign ces_12_21_io_ins_0 = ces_11_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_21_io_ins_1 = ces_12_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_21_io_ins_2 = ces_13_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_21_io_ins_3 = ces_12_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_22_clock = clock;
  assign ces_12_22_io_ins_0 = ces_11_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_22_io_ins_1 = ces_12_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_22_io_ins_2 = ces_13_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_22_io_ins_3 = ces_12_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_23_clock = clock;
  assign ces_12_23_io_ins_0 = ces_11_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_23_io_ins_1 = ces_12_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_23_io_ins_2 = ces_13_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_23_io_ins_3 = ces_12_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_24_clock = clock;
  assign ces_12_24_io_ins_0 = ces_11_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_24_io_ins_1 = ces_12_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_24_io_ins_2 = ces_13_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_24_io_ins_3 = ces_12_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_25_clock = clock;
  assign ces_12_25_io_ins_0 = ces_11_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_25_io_ins_1 = ces_12_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_25_io_ins_2 = ces_13_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_25_io_ins_3 = ces_12_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_26_clock = clock;
  assign ces_12_26_io_ins_0 = ces_11_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_26_io_ins_1 = ces_12_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_26_io_ins_2 = ces_13_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_26_io_ins_3 = ces_12_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_27_clock = clock;
  assign ces_12_27_io_ins_0 = ces_11_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_27_io_ins_1 = ces_12_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_27_io_ins_2 = ces_13_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_27_io_ins_3 = ces_12_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_28_clock = clock;
  assign ces_12_28_io_ins_0 = ces_11_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_28_io_ins_1 = ces_12_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_28_io_ins_2 = ces_13_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_28_io_ins_3 = ces_12_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_29_clock = clock;
  assign ces_12_29_io_ins_0 = ces_11_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_29_io_ins_1 = ces_12_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_29_io_ins_2 = ces_13_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_29_io_ins_3 = ces_12_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_30_clock = clock;
  assign ces_12_30_io_ins_0 = ces_11_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_30_io_ins_1 = ces_12_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_12_30_io_ins_2 = ces_13_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_30_io_ins_3 = ces_12_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_12_31_clock = clock;
  assign ces_12_31_io_ins_0 = ces_11_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_31_io_ins_1 = io_insVertical_0_12; // @[MockArray.scala 45:87]
  assign ces_12_31_io_ins_2 = ces_13_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_31_io_ins_3 = ces_12_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_0_clock = clock;
  assign ces_13_0_io_ins_0 = ces_12_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_0_io_ins_1 = ces_13_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_0_io_ins_2 = ces_14_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_0_io_ins_3 = io_insVertical_1_13; // @[MockArray.scala 47:87]
  assign ces_13_1_clock = clock;
  assign ces_13_1_io_ins_0 = ces_12_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_1_io_ins_1 = ces_13_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_1_io_ins_2 = ces_14_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_1_io_ins_3 = ces_13_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_2_clock = clock;
  assign ces_13_2_io_ins_0 = ces_12_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_2_io_ins_1 = ces_13_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_2_io_ins_2 = ces_14_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_2_io_ins_3 = ces_13_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_3_clock = clock;
  assign ces_13_3_io_ins_0 = ces_12_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_3_io_ins_1 = ces_13_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_3_io_ins_2 = ces_14_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_3_io_ins_3 = ces_13_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_4_clock = clock;
  assign ces_13_4_io_ins_0 = ces_12_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_4_io_ins_1 = ces_13_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_4_io_ins_2 = ces_14_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_4_io_ins_3 = ces_13_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_5_clock = clock;
  assign ces_13_5_io_ins_0 = ces_12_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_5_io_ins_1 = ces_13_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_5_io_ins_2 = ces_14_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_5_io_ins_3 = ces_13_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_6_clock = clock;
  assign ces_13_6_io_ins_0 = ces_12_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_6_io_ins_1 = ces_13_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_6_io_ins_2 = ces_14_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_6_io_ins_3 = ces_13_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_7_clock = clock;
  assign ces_13_7_io_ins_0 = ces_12_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_7_io_ins_1 = ces_13_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_7_io_ins_2 = ces_14_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_7_io_ins_3 = ces_13_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_8_clock = clock;
  assign ces_13_8_io_ins_0 = ces_12_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_8_io_ins_1 = ces_13_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_8_io_ins_2 = ces_14_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_8_io_ins_3 = ces_13_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_9_clock = clock;
  assign ces_13_9_io_ins_0 = ces_12_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_9_io_ins_1 = ces_13_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_9_io_ins_2 = ces_14_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_9_io_ins_3 = ces_13_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_10_clock = clock;
  assign ces_13_10_io_ins_0 = ces_12_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_10_io_ins_1 = ces_13_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_10_io_ins_2 = ces_14_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_10_io_ins_3 = ces_13_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_11_clock = clock;
  assign ces_13_11_io_ins_0 = ces_12_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_11_io_ins_1 = ces_13_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_11_io_ins_2 = ces_14_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_11_io_ins_3 = ces_13_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_12_clock = clock;
  assign ces_13_12_io_ins_0 = ces_12_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_12_io_ins_1 = ces_13_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_12_io_ins_2 = ces_14_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_12_io_ins_3 = ces_13_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_13_clock = clock;
  assign ces_13_13_io_ins_0 = ces_12_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_13_io_ins_1 = ces_13_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_13_io_ins_2 = ces_14_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_13_io_ins_3 = ces_13_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_14_clock = clock;
  assign ces_13_14_io_ins_0 = ces_12_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_14_io_ins_1 = ces_13_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_14_io_ins_2 = ces_14_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_14_io_ins_3 = ces_13_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_15_clock = clock;
  assign ces_13_15_io_ins_0 = ces_12_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_15_io_ins_1 = ces_13_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_15_io_ins_2 = ces_14_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_15_io_ins_3 = ces_13_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_16_clock = clock;
  assign ces_13_16_io_ins_0 = ces_12_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_16_io_ins_1 = ces_13_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_16_io_ins_2 = ces_14_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_16_io_ins_3 = ces_13_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_17_clock = clock;
  assign ces_13_17_io_ins_0 = ces_12_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_17_io_ins_1 = ces_13_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_17_io_ins_2 = ces_14_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_17_io_ins_3 = ces_13_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_18_clock = clock;
  assign ces_13_18_io_ins_0 = ces_12_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_18_io_ins_1 = ces_13_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_18_io_ins_2 = ces_14_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_18_io_ins_3 = ces_13_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_19_clock = clock;
  assign ces_13_19_io_ins_0 = ces_12_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_19_io_ins_1 = ces_13_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_19_io_ins_2 = ces_14_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_19_io_ins_3 = ces_13_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_20_clock = clock;
  assign ces_13_20_io_ins_0 = ces_12_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_20_io_ins_1 = ces_13_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_20_io_ins_2 = ces_14_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_20_io_ins_3 = ces_13_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_21_clock = clock;
  assign ces_13_21_io_ins_0 = ces_12_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_21_io_ins_1 = ces_13_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_21_io_ins_2 = ces_14_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_21_io_ins_3 = ces_13_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_22_clock = clock;
  assign ces_13_22_io_ins_0 = ces_12_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_22_io_ins_1 = ces_13_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_22_io_ins_2 = ces_14_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_22_io_ins_3 = ces_13_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_23_clock = clock;
  assign ces_13_23_io_ins_0 = ces_12_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_23_io_ins_1 = ces_13_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_23_io_ins_2 = ces_14_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_23_io_ins_3 = ces_13_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_24_clock = clock;
  assign ces_13_24_io_ins_0 = ces_12_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_24_io_ins_1 = ces_13_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_24_io_ins_2 = ces_14_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_24_io_ins_3 = ces_13_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_25_clock = clock;
  assign ces_13_25_io_ins_0 = ces_12_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_25_io_ins_1 = ces_13_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_25_io_ins_2 = ces_14_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_25_io_ins_3 = ces_13_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_26_clock = clock;
  assign ces_13_26_io_ins_0 = ces_12_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_26_io_ins_1 = ces_13_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_26_io_ins_2 = ces_14_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_26_io_ins_3 = ces_13_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_27_clock = clock;
  assign ces_13_27_io_ins_0 = ces_12_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_27_io_ins_1 = ces_13_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_27_io_ins_2 = ces_14_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_27_io_ins_3 = ces_13_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_28_clock = clock;
  assign ces_13_28_io_ins_0 = ces_12_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_28_io_ins_1 = ces_13_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_28_io_ins_2 = ces_14_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_28_io_ins_3 = ces_13_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_29_clock = clock;
  assign ces_13_29_io_ins_0 = ces_12_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_29_io_ins_1 = ces_13_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_29_io_ins_2 = ces_14_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_29_io_ins_3 = ces_13_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_30_clock = clock;
  assign ces_13_30_io_ins_0 = ces_12_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_30_io_ins_1 = ces_13_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_13_30_io_ins_2 = ces_14_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_30_io_ins_3 = ces_13_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_13_31_clock = clock;
  assign ces_13_31_io_ins_0 = ces_12_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_31_io_ins_1 = io_insVertical_0_13; // @[MockArray.scala 45:87]
  assign ces_13_31_io_ins_2 = ces_14_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_31_io_ins_3 = ces_13_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_0_clock = clock;
  assign ces_14_0_io_ins_0 = ces_13_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_0_io_ins_1 = ces_14_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_0_io_ins_2 = ces_15_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_0_io_ins_3 = io_insVertical_1_14; // @[MockArray.scala 47:87]
  assign ces_14_1_clock = clock;
  assign ces_14_1_io_ins_0 = ces_13_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_1_io_ins_1 = ces_14_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_1_io_ins_2 = ces_15_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_1_io_ins_3 = ces_14_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_2_clock = clock;
  assign ces_14_2_io_ins_0 = ces_13_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_2_io_ins_1 = ces_14_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_2_io_ins_2 = ces_15_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_2_io_ins_3 = ces_14_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_3_clock = clock;
  assign ces_14_3_io_ins_0 = ces_13_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_3_io_ins_1 = ces_14_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_3_io_ins_2 = ces_15_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_3_io_ins_3 = ces_14_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_4_clock = clock;
  assign ces_14_4_io_ins_0 = ces_13_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_4_io_ins_1 = ces_14_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_4_io_ins_2 = ces_15_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_4_io_ins_3 = ces_14_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_5_clock = clock;
  assign ces_14_5_io_ins_0 = ces_13_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_5_io_ins_1 = ces_14_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_5_io_ins_2 = ces_15_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_5_io_ins_3 = ces_14_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_6_clock = clock;
  assign ces_14_6_io_ins_0 = ces_13_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_6_io_ins_1 = ces_14_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_6_io_ins_2 = ces_15_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_6_io_ins_3 = ces_14_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_7_clock = clock;
  assign ces_14_7_io_ins_0 = ces_13_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_7_io_ins_1 = ces_14_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_7_io_ins_2 = ces_15_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_7_io_ins_3 = ces_14_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_8_clock = clock;
  assign ces_14_8_io_ins_0 = ces_13_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_8_io_ins_1 = ces_14_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_8_io_ins_2 = ces_15_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_8_io_ins_3 = ces_14_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_9_clock = clock;
  assign ces_14_9_io_ins_0 = ces_13_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_9_io_ins_1 = ces_14_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_9_io_ins_2 = ces_15_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_9_io_ins_3 = ces_14_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_10_clock = clock;
  assign ces_14_10_io_ins_0 = ces_13_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_10_io_ins_1 = ces_14_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_10_io_ins_2 = ces_15_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_10_io_ins_3 = ces_14_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_11_clock = clock;
  assign ces_14_11_io_ins_0 = ces_13_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_11_io_ins_1 = ces_14_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_11_io_ins_2 = ces_15_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_11_io_ins_3 = ces_14_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_12_clock = clock;
  assign ces_14_12_io_ins_0 = ces_13_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_12_io_ins_1 = ces_14_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_12_io_ins_2 = ces_15_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_12_io_ins_3 = ces_14_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_13_clock = clock;
  assign ces_14_13_io_ins_0 = ces_13_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_13_io_ins_1 = ces_14_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_13_io_ins_2 = ces_15_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_13_io_ins_3 = ces_14_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_14_clock = clock;
  assign ces_14_14_io_ins_0 = ces_13_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_14_io_ins_1 = ces_14_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_14_io_ins_2 = ces_15_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_14_io_ins_3 = ces_14_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_15_clock = clock;
  assign ces_14_15_io_ins_0 = ces_13_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_15_io_ins_1 = ces_14_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_15_io_ins_2 = ces_15_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_15_io_ins_3 = ces_14_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_16_clock = clock;
  assign ces_14_16_io_ins_0 = ces_13_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_16_io_ins_1 = ces_14_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_16_io_ins_2 = ces_15_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_16_io_ins_3 = ces_14_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_17_clock = clock;
  assign ces_14_17_io_ins_0 = ces_13_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_17_io_ins_1 = ces_14_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_17_io_ins_2 = ces_15_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_17_io_ins_3 = ces_14_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_18_clock = clock;
  assign ces_14_18_io_ins_0 = ces_13_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_18_io_ins_1 = ces_14_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_18_io_ins_2 = ces_15_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_18_io_ins_3 = ces_14_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_19_clock = clock;
  assign ces_14_19_io_ins_0 = ces_13_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_19_io_ins_1 = ces_14_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_19_io_ins_2 = ces_15_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_19_io_ins_3 = ces_14_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_20_clock = clock;
  assign ces_14_20_io_ins_0 = ces_13_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_20_io_ins_1 = ces_14_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_20_io_ins_2 = ces_15_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_20_io_ins_3 = ces_14_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_21_clock = clock;
  assign ces_14_21_io_ins_0 = ces_13_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_21_io_ins_1 = ces_14_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_21_io_ins_2 = ces_15_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_21_io_ins_3 = ces_14_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_22_clock = clock;
  assign ces_14_22_io_ins_0 = ces_13_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_22_io_ins_1 = ces_14_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_22_io_ins_2 = ces_15_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_22_io_ins_3 = ces_14_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_23_clock = clock;
  assign ces_14_23_io_ins_0 = ces_13_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_23_io_ins_1 = ces_14_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_23_io_ins_2 = ces_15_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_23_io_ins_3 = ces_14_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_24_clock = clock;
  assign ces_14_24_io_ins_0 = ces_13_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_24_io_ins_1 = ces_14_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_24_io_ins_2 = ces_15_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_24_io_ins_3 = ces_14_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_25_clock = clock;
  assign ces_14_25_io_ins_0 = ces_13_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_25_io_ins_1 = ces_14_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_25_io_ins_2 = ces_15_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_25_io_ins_3 = ces_14_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_26_clock = clock;
  assign ces_14_26_io_ins_0 = ces_13_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_26_io_ins_1 = ces_14_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_26_io_ins_2 = ces_15_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_26_io_ins_3 = ces_14_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_27_clock = clock;
  assign ces_14_27_io_ins_0 = ces_13_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_27_io_ins_1 = ces_14_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_27_io_ins_2 = ces_15_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_27_io_ins_3 = ces_14_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_28_clock = clock;
  assign ces_14_28_io_ins_0 = ces_13_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_28_io_ins_1 = ces_14_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_28_io_ins_2 = ces_15_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_28_io_ins_3 = ces_14_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_29_clock = clock;
  assign ces_14_29_io_ins_0 = ces_13_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_29_io_ins_1 = ces_14_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_29_io_ins_2 = ces_15_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_29_io_ins_3 = ces_14_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_30_clock = clock;
  assign ces_14_30_io_ins_0 = ces_13_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_30_io_ins_1 = ces_14_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_14_30_io_ins_2 = ces_15_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_30_io_ins_3 = ces_14_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_14_31_clock = clock;
  assign ces_14_31_io_ins_0 = ces_13_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_31_io_ins_1 = io_insVertical_0_14; // @[MockArray.scala 45:87]
  assign ces_14_31_io_ins_2 = ces_15_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_31_io_ins_3 = ces_14_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_0_clock = clock;
  assign ces_15_0_io_ins_0 = ces_14_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_0_io_ins_1 = ces_15_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_0_io_ins_2 = ces_16_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_0_io_ins_3 = io_insVertical_1_15; // @[MockArray.scala 47:87]
  assign ces_15_1_clock = clock;
  assign ces_15_1_io_ins_0 = ces_14_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_1_io_ins_1 = ces_15_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_1_io_ins_2 = ces_16_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_1_io_ins_3 = ces_15_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_2_clock = clock;
  assign ces_15_2_io_ins_0 = ces_14_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_2_io_ins_1 = ces_15_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_2_io_ins_2 = ces_16_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_2_io_ins_3 = ces_15_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_3_clock = clock;
  assign ces_15_3_io_ins_0 = ces_14_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_3_io_ins_1 = ces_15_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_3_io_ins_2 = ces_16_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_3_io_ins_3 = ces_15_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_4_clock = clock;
  assign ces_15_4_io_ins_0 = ces_14_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_4_io_ins_1 = ces_15_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_4_io_ins_2 = ces_16_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_4_io_ins_3 = ces_15_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_5_clock = clock;
  assign ces_15_5_io_ins_0 = ces_14_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_5_io_ins_1 = ces_15_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_5_io_ins_2 = ces_16_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_5_io_ins_3 = ces_15_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_6_clock = clock;
  assign ces_15_6_io_ins_0 = ces_14_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_6_io_ins_1 = ces_15_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_6_io_ins_2 = ces_16_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_6_io_ins_3 = ces_15_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_7_clock = clock;
  assign ces_15_7_io_ins_0 = ces_14_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_7_io_ins_1 = ces_15_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_7_io_ins_2 = ces_16_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_7_io_ins_3 = ces_15_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_8_clock = clock;
  assign ces_15_8_io_ins_0 = ces_14_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_8_io_ins_1 = ces_15_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_8_io_ins_2 = ces_16_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_8_io_ins_3 = ces_15_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_9_clock = clock;
  assign ces_15_9_io_ins_0 = ces_14_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_9_io_ins_1 = ces_15_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_9_io_ins_2 = ces_16_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_9_io_ins_3 = ces_15_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_10_clock = clock;
  assign ces_15_10_io_ins_0 = ces_14_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_10_io_ins_1 = ces_15_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_10_io_ins_2 = ces_16_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_10_io_ins_3 = ces_15_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_11_clock = clock;
  assign ces_15_11_io_ins_0 = ces_14_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_11_io_ins_1 = ces_15_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_11_io_ins_2 = ces_16_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_11_io_ins_3 = ces_15_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_12_clock = clock;
  assign ces_15_12_io_ins_0 = ces_14_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_12_io_ins_1 = ces_15_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_12_io_ins_2 = ces_16_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_12_io_ins_3 = ces_15_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_13_clock = clock;
  assign ces_15_13_io_ins_0 = ces_14_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_13_io_ins_1 = ces_15_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_13_io_ins_2 = ces_16_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_13_io_ins_3 = ces_15_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_14_clock = clock;
  assign ces_15_14_io_ins_0 = ces_14_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_14_io_ins_1 = ces_15_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_14_io_ins_2 = ces_16_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_14_io_ins_3 = ces_15_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_15_clock = clock;
  assign ces_15_15_io_ins_0 = ces_14_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_15_io_ins_1 = ces_15_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_15_io_ins_2 = ces_16_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_15_io_ins_3 = ces_15_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_16_clock = clock;
  assign ces_15_16_io_ins_0 = ces_14_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_16_io_ins_1 = ces_15_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_16_io_ins_2 = ces_16_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_16_io_ins_3 = ces_15_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_17_clock = clock;
  assign ces_15_17_io_ins_0 = ces_14_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_17_io_ins_1 = ces_15_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_17_io_ins_2 = ces_16_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_17_io_ins_3 = ces_15_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_18_clock = clock;
  assign ces_15_18_io_ins_0 = ces_14_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_18_io_ins_1 = ces_15_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_18_io_ins_2 = ces_16_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_18_io_ins_3 = ces_15_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_19_clock = clock;
  assign ces_15_19_io_ins_0 = ces_14_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_19_io_ins_1 = ces_15_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_19_io_ins_2 = ces_16_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_19_io_ins_3 = ces_15_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_20_clock = clock;
  assign ces_15_20_io_ins_0 = ces_14_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_20_io_ins_1 = ces_15_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_20_io_ins_2 = ces_16_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_20_io_ins_3 = ces_15_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_21_clock = clock;
  assign ces_15_21_io_ins_0 = ces_14_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_21_io_ins_1 = ces_15_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_21_io_ins_2 = ces_16_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_21_io_ins_3 = ces_15_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_22_clock = clock;
  assign ces_15_22_io_ins_0 = ces_14_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_22_io_ins_1 = ces_15_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_22_io_ins_2 = ces_16_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_22_io_ins_3 = ces_15_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_23_clock = clock;
  assign ces_15_23_io_ins_0 = ces_14_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_23_io_ins_1 = ces_15_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_23_io_ins_2 = ces_16_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_23_io_ins_3 = ces_15_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_24_clock = clock;
  assign ces_15_24_io_ins_0 = ces_14_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_24_io_ins_1 = ces_15_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_24_io_ins_2 = ces_16_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_24_io_ins_3 = ces_15_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_25_clock = clock;
  assign ces_15_25_io_ins_0 = ces_14_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_25_io_ins_1 = ces_15_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_25_io_ins_2 = ces_16_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_25_io_ins_3 = ces_15_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_26_clock = clock;
  assign ces_15_26_io_ins_0 = ces_14_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_26_io_ins_1 = ces_15_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_26_io_ins_2 = ces_16_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_26_io_ins_3 = ces_15_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_27_clock = clock;
  assign ces_15_27_io_ins_0 = ces_14_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_27_io_ins_1 = ces_15_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_27_io_ins_2 = ces_16_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_27_io_ins_3 = ces_15_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_28_clock = clock;
  assign ces_15_28_io_ins_0 = ces_14_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_28_io_ins_1 = ces_15_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_28_io_ins_2 = ces_16_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_28_io_ins_3 = ces_15_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_29_clock = clock;
  assign ces_15_29_io_ins_0 = ces_14_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_29_io_ins_1 = ces_15_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_29_io_ins_2 = ces_16_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_29_io_ins_3 = ces_15_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_30_clock = clock;
  assign ces_15_30_io_ins_0 = ces_14_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_30_io_ins_1 = ces_15_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_15_30_io_ins_2 = ces_16_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_30_io_ins_3 = ces_15_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_15_31_clock = clock;
  assign ces_15_31_io_ins_0 = ces_14_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_31_io_ins_1 = io_insVertical_0_15; // @[MockArray.scala 45:87]
  assign ces_15_31_io_ins_2 = ces_16_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_31_io_ins_3 = ces_15_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_0_clock = clock;
  assign ces_16_0_io_ins_0 = ces_15_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_0_io_ins_1 = ces_16_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_0_io_ins_2 = ces_17_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_0_io_ins_3 = io_insVertical_1_16; // @[MockArray.scala 47:87]
  assign ces_16_1_clock = clock;
  assign ces_16_1_io_ins_0 = ces_15_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_1_io_ins_1 = ces_16_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_1_io_ins_2 = ces_17_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_1_io_ins_3 = ces_16_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_2_clock = clock;
  assign ces_16_2_io_ins_0 = ces_15_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_2_io_ins_1 = ces_16_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_2_io_ins_2 = ces_17_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_2_io_ins_3 = ces_16_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_3_clock = clock;
  assign ces_16_3_io_ins_0 = ces_15_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_3_io_ins_1 = ces_16_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_3_io_ins_2 = ces_17_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_3_io_ins_3 = ces_16_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_4_clock = clock;
  assign ces_16_4_io_ins_0 = ces_15_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_4_io_ins_1 = ces_16_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_4_io_ins_2 = ces_17_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_4_io_ins_3 = ces_16_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_5_clock = clock;
  assign ces_16_5_io_ins_0 = ces_15_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_5_io_ins_1 = ces_16_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_5_io_ins_2 = ces_17_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_5_io_ins_3 = ces_16_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_6_clock = clock;
  assign ces_16_6_io_ins_0 = ces_15_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_6_io_ins_1 = ces_16_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_6_io_ins_2 = ces_17_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_6_io_ins_3 = ces_16_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_7_clock = clock;
  assign ces_16_7_io_ins_0 = ces_15_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_7_io_ins_1 = ces_16_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_7_io_ins_2 = ces_17_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_7_io_ins_3 = ces_16_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_8_clock = clock;
  assign ces_16_8_io_ins_0 = ces_15_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_8_io_ins_1 = ces_16_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_8_io_ins_2 = ces_17_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_8_io_ins_3 = ces_16_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_9_clock = clock;
  assign ces_16_9_io_ins_0 = ces_15_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_9_io_ins_1 = ces_16_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_9_io_ins_2 = ces_17_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_9_io_ins_3 = ces_16_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_10_clock = clock;
  assign ces_16_10_io_ins_0 = ces_15_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_10_io_ins_1 = ces_16_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_10_io_ins_2 = ces_17_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_10_io_ins_3 = ces_16_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_11_clock = clock;
  assign ces_16_11_io_ins_0 = ces_15_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_11_io_ins_1 = ces_16_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_11_io_ins_2 = ces_17_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_11_io_ins_3 = ces_16_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_12_clock = clock;
  assign ces_16_12_io_ins_0 = ces_15_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_12_io_ins_1 = ces_16_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_12_io_ins_2 = ces_17_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_12_io_ins_3 = ces_16_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_13_clock = clock;
  assign ces_16_13_io_ins_0 = ces_15_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_13_io_ins_1 = ces_16_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_13_io_ins_2 = ces_17_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_13_io_ins_3 = ces_16_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_14_clock = clock;
  assign ces_16_14_io_ins_0 = ces_15_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_14_io_ins_1 = ces_16_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_14_io_ins_2 = ces_17_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_14_io_ins_3 = ces_16_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_15_clock = clock;
  assign ces_16_15_io_ins_0 = ces_15_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_15_io_ins_1 = ces_16_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_15_io_ins_2 = ces_17_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_15_io_ins_3 = ces_16_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_16_clock = clock;
  assign ces_16_16_io_ins_0 = ces_15_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_16_io_ins_1 = ces_16_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_16_io_ins_2 = ces_17_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_16_io_ins_3 = ces_16_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_17_clock = clock;
  assign ces_16_17_io_ins_0 = ces_15_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_17_io_ins_1 = ces_16_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_17_io_ins_2 = ces_17_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_17_io_ins_3 = ces_16_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_18_clock = clock;
  assign ces_16_18_io_ins_0 = ces_15_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_18_io_ins_1 = ces_16_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_18_io_ins_2 = ces_17_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_18_io_ins_3 = ces_16_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_19_clock = clock;
  assign ces_16_19_io_ins_0 = ces_15_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_19_io_ins_1 = ces_16_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_19_io_ins_2 = ces_17_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_19_io_ins_3 = ces_16_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_20_clock = clock;
  assign ces_16_20_io_ins_0 = ces_15_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_20_io_ins_1 = ces_16_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_20_io_ins_2 = ces_17_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_20_io_ins_3 = ces_16_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_21_clock = clock;
  assign ces_16_21_io_ins_0 = ces_15_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_21_io_ins_1 = ces_16_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_21_io_ins_2 = ces_17_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_21_io_ins_3 = ces_16_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_22_clock = clock;
  assign ces_16_22_io_ins_0 = ces_15_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_22_io_ins_1 = ces_16_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_22_io_ins_2 = ces_17_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_22_io_ins_3 = ces_16_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_23_clock = clock;
  assign ces_16_23_io_ins_0 = ces_15_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_23_io_ins_1 = ces_16_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_23_io_ins_2 = ces_17_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_23_io_ins_3 = ces_16_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_24_clock = clock;
  assign ces_16_24_io_ins_0 = ces_15_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_24_io_ins_1 = ces_16_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_24_io_ins_2 = ces_17_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_24_io_ins_3 = ces_16_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_25_clock = clock;
  assign ces_16_25_io_ins_0 = ces_15_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_25_io_ins_1 = ces_16_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_25_io_ins_2 = ces_17_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_25_io_ins_3 = ces_16_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_26_clock = clock;
  assign ces_16_26_io_ins_0 = ces_15_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_26_io_ins_1 = ces_16_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_26_io_ins_2 = ces_17_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_26_io_ins_3 = ces_16_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_27_clock = clock;
  assign ces_16_27_io_ins_0 = ces_15_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_27_io_ins_1 = ces_16_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_27_io_ins_2 = ces_17_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_27_io_ins_3 = ces_16_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_28_clock = clock;
  assign ces_16_28_io_ins_0 = ces_15_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_28_io_ins_1 = ces_16_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_28_io_ins_2 = ces_17_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_28_io_ins_3 = ces_16_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_29_clock = clock;
  assign ces_16_29_io_ins_0 = ces_15_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_29_io_ins_1 = ces_16_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_29_io_ins_2 = ces_17_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_29_io_ins_3 = ces_16_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_30_clock = clock;
  assign ces_16_30_io_ins_0 = ces_15_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_30_io_ins_1 = ces_16_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_16_30_io_ins_2 = ces_17_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_30_io_ins_3 = ces_16_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_16_31_clock = clock;
  assign ces_16_31_io_ins_0 = ces_15_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_31_io_ins_1 = io_insVertical_0_16; // @[MockArray.scala 45:87]
  assign ces_16_31_io_ins_2 = ces_17_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_31_io_ins_3 = ces_16_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_0_clock = clock;
  assign ces_17_0_io_ins_0 = ces_16_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_0_io_ins_1 = ces_17_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_0_io_ins_2 = ces_18_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_0_io_ins_3 = io_insVertical_1_17; // @[MockArray.scala 47:87]
  assign ces_17_1_clock = clock;
  assign ces_17_1_io_ins_0 = ces_16_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_1_io_ins_1 = ces_17_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_1_io_ins_2 = ces_18_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_1_io_ins_3 = ces_17_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_2_clock = clock;
  assign ces_17_2_io_ins_0 = ces_16_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_2_io_ins_1 = ces_17_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_2_io_ins_2 = ces_18_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_2_io_ins_3 = ces_17_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_3_clock = clock;
  assign ces_17_3_io_ins_0 = ces_16_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_3_io_ins_1 = ces_17_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_3_io_ins_2 = ces_18_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_3_io_ins_3 = ces_17_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_4_clock = clock;
  assign ces_17_4_io_ins_0 = ces_16_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_4_io_ins_1 = ces_17_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_4_io_ins_2 = ces_18_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_4_io_ins_3 = ces_17_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_5_clock = clock;
  assign ces_17_5_io_ins_0 = ces_16_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_5_io_ins_1 = ces_17_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_5_io_ins_2 = ces_18_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_5_io_ins_3 = ces_17_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_6_clock = clock;
  assign ces_17_6_io_ins_0 = ces_16_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_6_io_ins_1 = ces_17_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_6_io_ins_2 = ces_18_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_6_io_ins_3 = ces_17_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_7_clock = clock;
  assign ces_17_7_io_ins_0 = ces_16_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_7_io_ins_1 = ces_17_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_7_io_ins_2 = ces_18_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_7_io_ins_3 = ces_17_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_8_clock = clock;
  assign ces_17_8_io_ins_0 = ces_16_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_8_io_ins_1 = ces_17_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_8_io_ins_2 = ces_18_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_8_io_ins_3 = ces_17_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_9_clock = clock;
  assign ces_17_9_io_ins_0 = ces_16_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_9_io_ins_1 = ces_17_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_9_io_ins_2 = ces_18_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_9_io_ins_3 = ces_17_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_10_clock = clock;
  assign ces_17_10_io_ins_0 = ces_16_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_10_io_ins_1 = ces_17_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_10_io_ins_2 = ces_18_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_10_io_ins_3 = ces_17_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_11_clock = clock;
  assign ces_17_11_io_ins_0 = ces_16_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_11_io_ins_1 = ces_17_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_11_io_ins_2 = ces_18_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_11_io_ins_3 = ces_17_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_12_clock = clock;
  assign ces_17_12_io_ins_0 = ces_16_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_12_io_ins_1 = ces_17_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_12_io_ins_2 = ces_18_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_12_io_ins_3 = ces_17_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_13_clock = clock;
  assign ces_17_13_io_ins_0 = ces_16_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_13_io_ins_1 = ces_17_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_13_io_ins_2 = ces_18_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_13_io_ins_3 = ces_17_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_14_clock = clock;
  assign ces_17_14_io_ins_0 = ces_16_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_14_io_ins_1 = ces_17_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_14_io_ins_2 = ces_18_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_14_io_ins_3 = ces_17_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_15_clock = clock;
  assign ces_17_15_io_ins_0 = ces_16_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_15_io_ins_1 = ces_17_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_15_io_ins_2 = ces_18_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_15_io_ins_3 = ces_17_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_16_clock = clock;
  assign ces_17_16_io_ins_0 = ces_16_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_16_io_ins_1 = ces_17_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_16_io_ins_2 = ces_18_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_16_io_ins_3 = ces_17_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_17_clock = clock;
  assign ces_17_17_io_ins_0 = ces_16_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_17_io_ins_1 = ces_17_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_17_io_ins_2 = ces_18_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_17_io_ins_3 = ces_17_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_18_clock = clock;
  assign ces_17_18_io_ins_0 = ces_16_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_18_io_ins_1 = ces_17_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_18_io_ins_2 = ces_18_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_18_io_ins_3 = ces_17_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_19_clock = clock;
  assign ces_17_19_io_ins_0 = ces_16_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_19_io_ins_1 = ces_17_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_19_io_ins_2 = ces_18_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_19_io_ins_3 = ces_17_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_20_clock = clock;
  assign ces_17_20_io_ins_0 = ces_16_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_20_io_ins_1 = ces_17_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_20_io_ins_2 = ces_18_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_20_io_ins_3 = ces_17_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_21_clock = clock;
  assign ces_17_21_io_ins_0 = ces_16_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_21_io_ins_1 = ces_17_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_21_io_ins_2 = ces_18_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_21_io_ins_3 = ces_17_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_22_clock = clock;
  assign ces_17_22_io_ins_0 = ces_16_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_22_io_ins_1 = ces_17_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_22_io_ins_2 = ces_18_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_22_io_ins_3 = ces_17_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_23_clock = clock;
  assign ces_17_23_io_ins_0 = ces_16_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_23_io_ins_1 = ces_17_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_23_io_ins_2 = ces_18_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_23_io_ins_3 = ces_17_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_24_clock = clock;
  assign ces_17_24_io_ins_0 = ces_16_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_24_io_ins_1 = ces_17_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_24_io_ins_2 = ces_18_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_24_io_ins_3 = ces_17_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_25_clock = clock;
  assign ces_17_25_io_ins_0 = ces_16_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_25_io_ins_1 = ces_17_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_25_io_ins_2 = ces_18_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_25_io_ins_3 = ces_17_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_26_clock = clock;
  assign ces_17_26_io_ins_0 = ces_16_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_26_io_ins_1 = ces_17_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_26_io_ins_2 = ces_18_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_26_io_ins_3 = ces_17_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_27_clock = clock;
  assign ces_17_27_io_ins_0 = ces_16_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_27_io_ins_1 = ces_17_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_27_io_ins_2 = ces_18_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_27_io_ins_3 = ces_17_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_28_clock = clock;
  assign ces_17_28_io_ins_0 = ces_16_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_28_io_ins_1 = ces_17_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_28_io_ins_2 = ces_18_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_28_io_ins_3 = ces_17_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_29_clock = clock;
  assign ces_17_29_io_ins_0 = ces_16_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_29_io_ins_1 = ces_17_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_29_io_ins_2 = ces_18_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_29_io_ins_3 = ces_17_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_30_clock = clock;
  assign ces_17_30_io_ins_0 = ces_16_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_30_io_ins_1 = ces_17_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_17_30_io_ins_2 = ces_18_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_30_io_ins_3 = ces_17_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_17_31_clock = clock;
  assign ces_17_31_io_ins_0 = ces_16_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_31_io_ins_1 = io_insVertical_0_17; // @[MockArray.scala 45:87]
  assign ces_17_31_io_ins_2 = ces_18_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_31_io_ins_3 = ces_17_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_0_clock = clock;
  assign ces_18_0_io_ins_0 = ces_17_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_0_io_ins_1 = ces_18_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_0_io_ins_2 = ces_19_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_0_io_ins_3 = io_insVertical_1_18; // @[MockArray.scala 47:87]
  assign ces_18_1_clock = clock;
  assign ces_18_1_io_ins_0 = ces_17_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_1_io_ins_1 = ces_18_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_1_io_ins_2 = ces_19_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_1_io_ins_3 = ces_18_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_2_clock = clock;
  assign ces_18_2_io_ins_0 = ces_17_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_2_io_ins_1 = ces_18_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_2_io_ins_2 = ces_19_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_2_io_ins_3 = ces_18_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_3_clock = clock;
  assign ces_18_3_io_ins_0 = ces_17_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_3_io_ins_1 = ces_18_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_3_io_ins_2 = ces_19_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_3_io_ins_3 = ces_18_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_4_clock = clock;
  assign ces_18_4_io_ins_0 = ces_17_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_4_io_ins_1 = ces_18_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_4_io_ins_2 = ces_19_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_4_io_ins_3 = ces_18_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_5_clock = clock;
  assign ces_18_5_io_ins_0 = ces_17_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_5_io_ins_1 = ces_18_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_5_io_ins_2 = ces_19_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_5_io_ins_3 = ces_18_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_6_clock = clock;
  assign ces_18_6_io_ins_0 = ces_17_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_6_io_ins_1 = ces_18_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_6_io_ins_2 = ces_19_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_6_io_ins_3 = ces_18_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_7_clock = clock;
  assign ces_18_7_io_ins_0 = ces_17_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_7_io_ins_1 = ces_18_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_7_io_ins_2 = ces_19_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_7_io_ins_3 = ces_18_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_8_clock = clock;
  assign ces_18_8_io_ins_0 = ces_17_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_8_io_ins_1 = ces_18_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_8_io_ins_2 = ces_19_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_8_io_ins_3 = ces_18_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_9_clock = clock;
  assign ces_18_9_io_ins_0 = ces_17_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_9_io_ins_1 = ces_18_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_9_io_ins_2 = ces_19_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_9_io_ins_3 = ces_18_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_10_clock = clock;
  assign ces_18_10_io_ins_0 = ces_17_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_10_io_ins_1 = ces_18_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_10_io_ins_2 = ces_19_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_10_io_ins_3 = ces_18_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_11_clock = clock;
  assign ces_18_11_io_ins_0 = ces_17_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_11_io_ins_1 = ces_18_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_11_io_ins_2 = ces_19_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_11_io_ins_3 = ces_18_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_12_clock = clock;
  assign ces_18_12_io_ins_0 = ces_17_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_12_io_ins_1 = ces_18_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_12_io_ins_2 = ces_19_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_12_io_ins_3 = ces_18_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_13_clock = clock;
  assign ces_18_13_io_ins_0 = ces_17_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_13_io_ins_1 = ces_18_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_13_io_ins_2 = ces_19_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_13_io_ins_3 = ces_18_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_14_clock = clock;
  assign ces_18_14_io_ins_0 = ces_17_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_14_io_ins_1 = ces_18_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_14_io_ins_2 = ces_19_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_14_io_ins_3 = ces_18_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_15_clock = clock;
  assign ces_18_15_io_ins_0 = ces_17_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_15_io_ins_1 = ces_18_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_15_io_ins_2 = ces_19_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_15_io_ins_3 = ces_18_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_16_clock = clock;
  assign ces_18_16_io_ins_0 = ces_17_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_16_io_ins_1 = ces_18_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_16_io_ins_2 = ces_19_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_16_io_ins_3 = ces_18_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_17_clock = clock;
  assign ces_18_17_io_ins_0 = ces_17_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_17_io_ins_1 = ces_18_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_17_io_ins_2 = ces_19_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_17_io_ins_3 = ces_18_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_18_clock = clock;
  assign ces_18_18_io_ins_0 = ces_17_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_18_io_ins_1 = ces_18_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_18_io_ins_2 = ces_19_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_18_io_ins_3 = ces_18_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_19_clock = clock;
  assign ces_18_19_io_ins_0 = ces_17_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_19_io_ins_1 = ces_18_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_19_io_ins_2 = ces_19_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_19_io_ins_3 = ces_18_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_20_clock = clock;
  assign ces_18_20_io_ins_0 = ces_17_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_20_io_ins_1 = ces_18_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_20_io_ins_2 = ces_19_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_20_io_ins_3 = ces_18_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_21_clock = clock;
  assign ces_18_21_io_ins_0 = ces_17_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_21_io_ins_1 = ces_18_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_21_io_ins_2 = ces_19_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_21_io_ins_3 = ces_18_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_22_clock = clock;
  assign ces_18_22_io_ins_0 = ces_17_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_22_io_ins_1 = ces_18_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_22_io_ins_2 = ces_19_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_22_io_ins_3 = ces_18_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_23_clock = clock;
  assign ces_18_23_io_ins_0 = ces_17_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_23_io_ins_1 = ces_18_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_23_io_ins_2 = ces_19_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_23_io_ins_3 = ces_18_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_24_clock = clock;
  assign ces_18_24_io_ins_0 = ces_17_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_24_io_ins_1 = ces_18_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_24_io_ins_2 = ces_19_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_24_io_ins_3 = ces_18_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_25_clock = clock;
  assign ces_18_25_io_ins_0 = ces_17_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_25_io_ins_1 = ces_18_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_25_io_ins_2 = ces_19_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_25_io_ins_3 = ces_18_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_26_clock = clock;
  assign ces_18_26_io_ins_0 = ces_17_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_26_io_ins_1 = ces_18_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_26_io_ins_2 = ces_19_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_26_io_ins_3 = ces_18_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_27_clock = clock;
  assign ces_18_27_io_ins_0 = ces_17_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_27_io_ins_1 = ces_18_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_27_io_ins_2 = ces_19_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_27_io_ins_3 = ces_18_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_28_clock = clock;
  assign ces_18_28_io_ins_0 = ces_17_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_28_io_ins_1 = ces_18_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_28_io_ins_2 = ces_19_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_28_io_ins_3 = ces_18_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_29_clock = clock;
  assign ces_18_29_io_ins_0 = ces_17_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_29_io_ins_1 = ces_18_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_29_io_ins_2 = ces_19_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_29_io_ins_3 = ces_18_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_30_clock = clock;
  assign ces_18_30_io_ins_0 = ces_17_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_30_io_ins_1 = ces_18_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_18_30_io_ins_2 = ces_19_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_30_io_ins_3 = ces_18_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_18_31_clock = clock;
  assign ces_18_31_io_ins_0 = ces_17_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_31_io_ins_1 = io_insVertical_0_18; // @[MockArray.scala 45:87]
  assign ces_18_31_io_ins_2 = ces_19_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_31_io_ins_3 = ces_18_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_0_clock = clock;
  assign ces_19_0_io_ins_0 = ces_18_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_0_io_ins_1 = ces_19_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_0_io_ins_2 = ces_20_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_0_io_ins_3 = io_insVertical_1_19; // @[MockArray.scala 47:87]
  assign ces_19_1_clock = clock;
  assign ces_19_1_io_ins_0 = ces_18_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_1_io_ins_1 = ces_19_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_1_io_ins_2 = ces_20_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_1_io_ins_3 = ces_19_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_2_clock = clock;
  assign ces_19_2_io_ins_0 = ces_18_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_2_io_ins_1 = ces_19_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_2_io_ins_2 = ces_20_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_2_io_ins_3 = ces_19_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_3_clock = clock;
  assign ces_19_3_io_ins_0 = ces_18_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_3_io_ins_1 = ces_19_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_3_io_ins_2 = ces_20_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_3_io_ins_3 = ces_19_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_4_clock = clock;
  assign ces_19_4_io_ins_0 = ces_18_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_4_io_ins_1 = ces_19_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_4_io_ins_2 = ces_20_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_4_io_ins_3 = ces_19_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_5_clock = clock;
  assign ces_19_5_io_ins_0 = ces_18_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_5_io_ins_1 = ces_19_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_5_io_ins_2 = ces_20_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_5_io_ins_3 = ces_19_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_6_clock = clock;
  assign ces_19_6_io_ins_0 = ces_18_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_6_io_ins_1 = ces_19_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_6_io_ins_2 = ces_20_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_6_io_ins_3 = ces_19_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_7_clock = clock;
  assign ces_19_7_io_ins_0 = ces_18_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_7_io_ins_1 = ces_19_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_7_io_ins_2 = ces_20_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_7_io_ins_3 = ces_19_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_8_clock = clock;
  assign ces_19_8_io_ins_0 = ces_18_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_8_io_ins_1 = ces_19_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_8_io_ins_2 = ces_20_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_8_io_ins_3 = ces_19_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_9_clock = clock;
  assign ces_19_9_io_ins_0 = ces_18_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_9_io_ins_1 = ces_19_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_9_io_ins_2 = ces_20_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_9_io_ins_3 = ces_19_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_10_clock = clock;
  assign ces_19_10_io_ins_0 = ces_18_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_10_io_ins_1 = ces_19_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_10_io_ins_2 = ces_20_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_10_io_ins_3 = ces_19_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_11_clock = clock;
  assign ces_19_11_io_ins_0 = ces_18_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_11_io_ins_1 = ces_19_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_11_io_ins_2 = ces_20_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_11_io_ins_3 = ces_19_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_12_clock = clock;
  assign ces_19_12_io_ins_0 = ces_18_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_12_io_ins_1 = ces_19_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_12_io_ins_2 = ces_20_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_12_io_ins_3 = ces_19_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_13_clock = clock;
  assign ces_19_13_io_ins_0 = ces_18_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_13_io_ins_1 = ces_19_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_13_io_ins_2 = ces_20_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_13_io_ins_3 = ces_19_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_14_clock = clock;
  assign ces_19_14_io_ins_0 = ces_18_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_14_io_ins_1 = ces_19_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_14_io_ins_2 = ces_20_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_14_io_ins_3 = ces_19_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_15_clock = clock;
  assign ces_19_15_io_ins_0 = ces_18_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_15_io_ins_1 = ces_19_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_15_io_ins_2 = ces_20_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_15_io_ins_3 = ces_19_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_16_clock = clock;
  assign ces_19_16_io_ins_0 = ces_18_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_16_io_ins_1 = ces_19_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_16_io_ins_2 = ces_20_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_16_io_ins_3 = ces_19_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_17_clock = clock;
  assign ces_19_17_io_ins_0 = ces_18_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_17_io_ins_1 = ces_19_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_17_io_ins_2 = ces_20_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_17_io_ins_3 = ces_19_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_18_clock = clock;
  assign ces_19_18_io_ins_0 = ces_18_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_18_io_ins_1 = ces_19_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_18_io_ins_2 = ces_20_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_18_io_ins_3 = ces_19_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_19_clock = clock;
  assign ces_19_19_io_ins_0 = ces_18_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_19_io_ins_1 = ces_19_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_19_io_ins_2 = ces_20_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_19_io_ins_3 = ces_19_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_20_clock = clock;
  assign ces_19_20_io_ins_0 = ces_18_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_20_io_ins_1 = ces_19_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_20_io_ins_2 = ces_20_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_20_io_ins_3 = ces_19_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_21_clock = clock;
  assign ces_19_21_io_ins_0 = ces_18_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_21_io_ins_1 = ces_19_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_21_io_ins_2 = ces_20_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_21_io_ins_3 = ces_19_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_22_clock = clock;
  assign ces_19_22_io_ins_0 = ces_18_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_22_io_ins_1 = ces_19_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_22_io_ins_2 = ces_20_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_22_io_ins_3 = ces_19_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_23_clock = clock;
  assign ces_19_23_io_ins_0 = ces_18_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_23_io_ins_1 = ces_19_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_23_io_ins_2 = ces_20_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_23_io_ins_3 = ces_19_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_24_clock = clock;
  assign ces_19_24_io_ins_0 = ces_18_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_24_io_ins_1 = ces_19_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_24_io_ins_2 = ces_20_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_24_io_ins_3 = ces_19_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_25_clock = clock;
  assign ces_19_25_io_ins_0 = ces_18_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_25_io_ins_1 = ces_19_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_25_io_ins_2 = ces_20_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_25_io_ins_3 = ces_19_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_26_clock = clock;
  assign ces_19_26_io_ins_0 = ces_18_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_26_io_ins_1 = ces_19_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_26_io_ins_2 = ces_20_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_26_io_ins_3 = ces_19_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_27_clock = clock;
  assign ces_19_27_io_ins_0 = ces_18_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_27_io_ins_1 = ces_19_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_27_io_ins_2 = ces_20_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_27_io_ins_3 = ces_19_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_28_clock = clock;
  assign ces_19_28_io_ins_0 = ces_18_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_28_io_ins_1 = ces_19_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_28_io_ins_2 = ces_20_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_28_io_ins_3 = ces_19_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_29_clock = clock;
  assign ces_19_29_io_ins_0 = ces_18_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_29_io_ins_1 = ces_19_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_29_io_ins_2 = ces_20_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_29_io_ins_3 = ces_19_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_30_clock = clock;
  assign ces_19_30_io_ins_0 = ces_18_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_30_io_ins_1 = ces_19_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_19_30_io_ins_2 = ces_20_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_30_io_ins_3 = ces_19_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_19_31_clock = clock;
  assign ces_19_31_io_ins_0 = ces_18_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_31_io_ins_1 = io_insVertical_0_19; // @[MockArray.scala 45:87]
  assign ces_19_31_io_ins_2 = ces_20_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_31_io_ins_3 = ces_19_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_0_clock = clock;
  assign ces_20_0_io_ins_0 = ces_19_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_0_io_ins_1 = ces_20_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_0_io_ins_2 = ces_21_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_0_io_ins_3 = io_insVertical_1_20; // @[MockArray.scala 47:87]
  assign ces_20_1_clock = clock;
  assign ces_20_1_io_ins_0 = ces_19_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_1_io_ins_1 = ces_20_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_1_io_ins_2 = ces_21_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_1_io_ins_3 = ces_20_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_2_clock = clock;
  assign ces_20_2_io_ins_0 = ces_19_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_2_io_ins_1 = ces_20_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_2_io_ins_2 = ces_21_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_2_io_ins_3 = ces_20_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_3_clock = clock;
  assign ces_20_3_io_ins_0 = ces_19_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_3_io_ins_1 = ces_20_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_3_io_ins_2 = ces_21_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_3_io_ins_3 = ces_20_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_4_clock = clock;
  assign ces_20_4_io_ins_0 = ces_19_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_4_io_ins_1 = ces_20_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_4_io_ins_2 = ces_21_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_4_io_ins_3 = ces_20_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_5_clock = clock;
  assign ces_20_5_io_ins_0 = ces_19_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_5_io_ins_1 = ces_20_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_5_io_ins_2 = ces_21_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_5_io_ins_3 = ces_20_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_6_clock = clock;
  assign ces_20_6_io_ins_0 = ces_19_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_6_io_ins_1 = ces_20_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_6_io_ins_2 = ces_21_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_6_io_ins_3 = ces_20_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_7_clock = clock;
  assign ces_20_7_io_ins_0 = ces_19_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_7_io_ins_1 = ces_20_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_7_io_ins_2 = ces_21_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_7_io_ins_3 = ces_20_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_8_clock = clock;
  assign ces_20_8_io_ins_0 = ces_19_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_8_io_ins_1 = ces_20_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_8_io_ins_2 = ces_21_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_8_io_ins_3 = ces_20_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_9_clock = clock;
  assign ces_20_9_io_ins_0 = ces_19_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_9_io_ins_1 = ces_20_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_9_io_ins_2 = ces_21_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_9_io_ins_3 = ces_20_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_10_clock = clock;
  assign ces_20_10_io_ins_0 = ces_19_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_10_io_ins_1 = ces_20_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_10_io_ins_2 = ces_21_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_10_io_ins_3 = ces_20_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_11_clock = clock;
  assign ces_20_11_io_ins_0 = ces_19_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_11_io_ins_1 = ces_20_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_11_io_ins_2 = ces_21_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_11_io_ins_3 = ces_20_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_12_clock = clock;
  assign ces_20_12_io_ins_0 = ces_19_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_12_io_ins_1 = ces_20_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_12_io_ins_2 = ces_21_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_12_io_ins_3 = ces_20_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_13_clock = clock;
  assign ces_20_13_io_ins_0 = ces_19_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_13_io_ins_1 = ces_20_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_13_io_ins_2 = ces_21_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_13_io_ins_3 = ces_20_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_14_clock = clock;
  assign ces_20_14_io_ins_0 = ces_19_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_14_io_ins_1 = ces_20_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_14_io_ins_2 = ces_21_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_14_io_ins_3 = ces_20_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_15_clock = clock;
  assign ces_20_15_io_ins_0 = ces_19_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_15_io_ins_1 = ces_20_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_15_io_ins_2 = ces_21_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_15_io_ins_3 = ces_20_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_16_clock = clock;
  assign ces_20_16_io_ins_0 = ces_19_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_16_io_ins_1 = ces_20_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_16_io_ins_2 = ces_21_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_16_io_ins_3 = ces_20_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_17_clock = clock;
  assign ces_20_17_io_ins_0 = ces_19_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_17_io_ins_1 = ces_20_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_17_io_ins_2 = ces_21_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_17_io_ins_3 = ces_20_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_18_clock = clock;
  assign ces_20_18_io_ins_0 = ces_19_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_18_io_ins_1 = ces_20_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_18_io_ins_2 = ces_21_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_18_io_ins_3 = ces_20_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_19_clock = clock;
  assign ces_20_19_io_ins_0 = ces_19_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_19_io_ins_1 = ces_20_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_19_io_ins_2 = ces_21_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_19_io_ins_3 = ces_20_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_20_clock = clock;
  assign ces_20_20_io_ins_0 = ces_19_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_20_io_ins_1 = ces_20_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_20_io_ins_2 = ces_21_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_20_io_ins_3 = ces_20_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_21_clock = clock;
  assign ces_20_21_io_ins_0 = ces_19_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_21_io_ins_1 = ces_20_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_21_io_ins_2 = ces_21_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_21_io_ins_3 = ces_20_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_22_clock = clock;
  assign ces_20_22_io_ins_0 = ces_19_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_22_io_ins_1 = ces_20_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_22_io_ins_2 = ces_21_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_22_io_ins_3 = ces_20_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_23_clock = clock;
  assign ces_20_23_io_ins_0 = ces_19_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_23_io_ins_1 = ces_20_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_23_io_ins_2 = ces_21_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_23_io_ins_3 = ces_20_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_24_clock = clock;
  assign ces_20_24_io_ins_0 = ces_19_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_24_io_ins_1 = ces_20_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_24_io_ins_2 = ces_21_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_24_io_ins_3 = ces_20_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_25_clock = clock;
  assign ces_20_25_io_ins_0 = ces_19_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_25_io_ins_1 = ces_20_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_25_io_ins_2 = ces_21_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_25_io_ins_3 = ces_20_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_26_clock = clock;
  assign ces_20_26_io_ins_0 = ces_19_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_26_io_ins_1 = ces_20_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_26_io_ins_2 = ces_21_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_26_io_ins_3 = ces_20_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_27_clock = clock;
  assign ces_20_27_io_ins_0 = ces_19_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_27_io_ins_1 = ces_20_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_27_io_ins_2 = ces_21_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_27_io_ins_3 = ces_20_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_28_clock = clock;
  assign ces_20_28_io_ins_0 = ces_19_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_28_io_ins_1 = ces_20_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_28_io_ins_2 = ces_21_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_28_io_ins_3 = ces_20_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_29_clock = clock;
  assign ces_20_29_io_ins_0 = ces_19_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_29_io_ins_1 = ces_20_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_29_io_ins_2 = ces_21_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_29_io_ins_3 = ces_20_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_30_clock = clock;
  assign ces_20_30_io_ins_0 = ces_19_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_30_io_ins_1 = ces_20_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_20_30_io_ins_2 = ces_21_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_30_io_ins_3 = ces_20_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_20_31_clock = clock;
  assign ces_20_31_io_ins_0 = ces_19_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_31_io_ins_1 = io_insVertical_0_20; // @[MockArray.scala 45:87]
  assign ces_20_31_io_ins_2 = ces_21_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_31_io_ins_3 = ces_20_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_0_clock = clock;
  assign ces_21_0_io_ins_0 = ces_20_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_0_io_ins_1 = ces_21_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_0_io_ins_2 = ces_22_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_0_io_ins_3 = io_insVertical_1_21; // @[MockArray.scala 47:87]
  assign ces_21_1_clock = clock;
  assign ces_21_1_io_ins_0 = ces_20_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_1_io_ins_1 = ces_21_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_1_io_ins_2 = ces_22_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_1_io_ins_3 = ces_21_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_2_clock = clock;
  assign ces_21_2_io_ins_0 = ces_20_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_2_io_ins_1 = ces_21_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_2_io_ins_2 = ces_22_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_2_io_ins_3 = ces_21_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_3_clock = clock;
  assign ces_21_3_io_ins_0 = ces_20_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_3_io_ins_1 = ces_21_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_3_io_ins_2 = ces_22_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_3_io_ins_3 = ces_21_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_4_clock = clock;
  assign ces_21_4_io_ins_0 = ces_20_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_4_io_ins_1 = ces_21_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_4_io_ins_2 = ces_22_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_4_io_ins_3 = ces_21_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_5_clock = clock;
  assign ces_21_5_io_ins_0 = ces_20_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_5_io_ins_1 = ces_21_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_5_io_ins_2 = ces_22_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_5_io_ins_3 = ces_21_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_6_clock = clock;
  assign ces_21_6_io_ins_0 = ces_20_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_6_io_ins_1 = ces_21_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_6_io_ins_2 = ces_22_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_6_io_ins_3 = ces_21_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_7_clock = clock;
  assign ces_21_7_io_ins_0 = ces_20_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_7_io_ins_1 = ces_21_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_7_io_ins_2 = ces_22_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_7_io_ins_3 = ces_21_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_8_clock = clock;
  assign ces_21_8_io_ins_0 = ces_20_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_8_io_ins_1 = ces_21_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_8_io_ins_2 = ces_22_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_8_io_ins_3 = ces_21_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_9_clock = clock;
  assign ces_21_9_io_ins_0 = ces_20_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_9_io_ins_1 = ces_21_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_9_io_ins_2 = ces_22_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_9_io_ins_3 = ces_21_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_10_clock = clock;
  assign ces_21_10_io_ins_0 = ces_20_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_10_io_ins_1 = ces_21_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_10_io_ins_2 = ces_22_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_10_io_ins_3 = ces_21_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_11_clock = clock;
  assign ces_21_11_io_ins_0 = ces_20_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_11_io_ins_1 = ces_21_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_11_io_ins_2 = ces_22_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_11_io_ins_3 = ces_21_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_12_clock = clock;
  assign ces_21_12_io_ins_0 = ces_20_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_12_io_ins_1 = ces_21_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_12_io_ins_2 = ces_22_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_12_io_ins_3 = ces_21_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_13_clock = clock;
  assign ces_21_13_io_ins_0 = ces_20_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_13_io_ins_1 = ces_21_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_13_io_ins_2 = ces_22_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_13_io_ins_3 = ces_21_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_14_clock = clock;
  assign ces_21_14_io_ins_0 = ces_20_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_14_io_ins_1 = ces_21_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_14_io_ins_2 = ces_22_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_14_io_ins_3 = ces_21_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_15_clock = clock;
  assign ces_21_15_io_ins_0 = ces_20_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_15_io_ins_1 = ces_21_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_15_io_ins_2 = ces_22_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_15_io_ins_3 = ces_21_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_16_clock = clock;
  assign ces_21_16_io_ins_0 = ces_20_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_16_io_ins_1 = ces_21_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_16_io_ins_2 = ces_22_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_16_io_ins_3 = ces_21_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_17_clock = clock;
  assign ces_21_17_io_ins_0 = ces_20_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_17_io_ins_1 = ces_21_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_17_io_ins_2 = ces_22_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_17_io_ins_3 = ces_21_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_18_clock = clock;
  assign ces_21_18_io_ins_0 = ces_20_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_18_io_ins_1 = ces_21_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_18_io_ins_2 = ces_22_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_18_io_ins_3 = ces_21_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_19_clock = clock;
  assign ces_21_19_io_ins_0 = ces_20_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_19_io_ins_1 = ces_21_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_19_io_ins_2 = ces_22_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_19_io_ins_3 = ces_21_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_20_clock = clock;
  assign ces_21_20_io_ins_0 = ces_20_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_20_io_ins_1 = ces_21_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_20_io_ins_2 = ces_22_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_20_io_ins_3 = ces_21_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_21_clock = clock;
  assign ces_21_21_io_ins_0 = ces_20_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_21_io_ins_1 = ces_21_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_21_io_ins_2 = ces_22_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_21_io_ins_3 = ces_21_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_22_clock = clock;
  assign ces_21_22_io_ins_0 = ces_20_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_22_io_ins_1 = ces_21_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_22_io_ins_2 = ces_22_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_22_io_ins_3 = ces_21_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_23_clock = clock;
  assign ces_21_23_io_ins_0 = ces_20_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_23_io_ins_1 = ces_21_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_23_io_ins_2 = ces_22_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_23_io_ins_3 = ces_21_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_24_clock = clock;
  assign ces_21_24_io_ins_0 = ces_20_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_24_io_ins_1 = ces_21_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_24_io_ins_2 = ces_22_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_24_io_ins_3 = ces_21_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_25_clock = clock;
  assign ces_21_25_io_ins_0 = ces_20_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_25_io_ins_1 = ces_21_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_25_io_ins_2 = ces_22_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_25_io_ins_3 = ces_21_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_26_clock = clock;
  assign ces_21_26_io_ins_0 = ces_20_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_26_io_ins_1 = ces_21_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_26_io_ins_2 = ces_22_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_26_io_ins_3 = ces_21_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_27_clock = clock;
  assign ces_21_27_io_ins_0 = ces_20_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_27_io_ins_1 = ces_21_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_27_io_ins_2 = ces_22_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_27_io_ins_3 = ces_21_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_28_clock = clock;
  assign ces_21_28_io_ins_0 = ces_20_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_28_io_ins_1 = ces_21_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_28_io_ins_2 = ces_22_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_28_io_ins_3 = ces_21_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_29_clock = clock;
  assign ces_21_29_io_ins_0 = ces_20_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_29_io_ins_1 = ces_21_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_29_io_ins_2 = ces_22_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_29_io_ins_3 = ces_21_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_30_clock = clock;
  assign ces_21_30_io_ins_0 = ces_20_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_30_io_ins_1 = ces_21_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_21_30_io_ins_2 = ces_22_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_30_io_ins_3 = ces_21_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_21_31_clock = clock;
  assign ces_21_31_io_ins_0 = ces_20_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_31_io_ins_1 = io_insVertical_0_21; // @[MockArray.scala 45:87]
  assign ces_21_31_io_ins_2 = ces_22_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_31_io_ins_3 = ces_21_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_0_clock = clock;
  assign ces_22_0_io_ins_0 = ces_21_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_0_io_ins_1 = ces_22_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_0_io_ins_2 = ces_23_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_0_io_ins_3 = io_insVertical_1_22; // @[MockArray.scala 47:87]
  assign ces_22_1_clock = clock;
  assign ces_22_1_io_ins_0 = ces_21_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_1_io_ins_1 = ces_22_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_1_io_ins_2 = ces_23_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_1_io_ins_3 = ces_22_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_2_clock = clock;
  assign ces_22_2_io_ins_0 = ces_21_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_2_io_ins_1 = ces_22_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_2_io_ins_2 = ces_23_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_2_io_ins_3 = ces_22_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_3_clock = clock;
  assign ces_22_3_io_ins_0 = ces_21_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_3_io_ins_1 = ces_22_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_3_io_ins_2 = ces_23_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_3_io_ins_3 = ces_22_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_4_clock = clock;
  assign ces_22_4_io_ins_0 = ces_21_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_4_io_ins_1 = ces_22_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_4_io_ins_2 = ces_23_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_4_io_ins_3 = ces_22_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_5_clock = clock;
  assign ces_22_5_io_ins_0 = ces_21_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_5_io_ins_1 = ces_22_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_5_io_ins_2 = ces_23_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_5_io_ins_3 = ces_22_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_6_clock = clock;
  assign ces_22_6_io_ins_0 = ces_21_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_6_io_ins_1 = ces_22_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_6_io_ins_2 = ces_23_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_6_io_ins_3 = ces_22_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_7_clock = clock;
  assign ces_22_7_io_ins_0 = ces_21_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_7_io_ins_1 = ces_22_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_7_io_ins_2 = ces_23_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_7_io_ins_3 = ces_22_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_8_clock = clock;
  assign ces_22_8_io_ins_0 = ces_21_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_8_io_ins_1 = ces_22_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_8_io_ins_2 = ces_23_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_8_io_ins_3 = ces_22_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_9_clock = clock;
  assign ces_22_9_io_ins_0 = ces_21_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_9_io_ins_1 = ces_22_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_9_io_ins_2 = ces_23_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_9_io_ins_3 = ces_22_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_10_clock = clock;
  assign ces_22_10_io_ins_0 = ces_21_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_10_io_ins_1 = ces_22_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_10_io_ins_2 = ces_23_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_10_io_ins_3 = ces_22_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_11_clock = clock;
  assign ces_22_11_io_ins_0 = ces_21_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_11_io_ins_1 = ces_22_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_11_io_ins_2 = ces_23_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_11_io_ins_3 = ces_22_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_12_clock = clock;
  assign ces_22_12_io_ins_0 = ces_21_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_12_io_ins_1 = ces_22_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_12_io_ins_2 = ces_23_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_12_io_ins_3 = ces_22_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_13_clock = clock;
  assign ces_22_13_io_ins_0 = ces_21_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_13_io_ins_1 = ces_22_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_13_io_ins_2 = ces_23_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_13_io_ins_3 = ces_22_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_14_clock = clock;
  assign ces_22_14_io_ins_0 = ces_21_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_14_io_ins_1 = ces_22_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_14_io_ins_2 = ces_23_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_14_io_ins_3 = ces_22_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_15_clock = clock;
  assign ces_22_15_io_ins_0 = ces_21_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_15_io_ins_1 = ces_22_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_15_io_ins_2 = ces_23_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_15_io_ins_3 = ces_22_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_16_clock = clock;
  assign ces_22_16_io_ins_0 = ces_21_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_16_io_ins_1 = ces_22_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_16_io_ins_2 = ces_23_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_16_io_ins_3 = ces_22_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_17_clock = clock;
  assign ces_22_17_io_ins_0 = ces_21_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_17_io_ins_1 = ces_22_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_17_io_ins_2 = ces_23_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_17_io_ins_3 = ces_22_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_18_clock = clock;
  assign ces_22_18_io_ins_0 = ces_21_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_18_io_ins_1 = ces_22_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_18_io_ins_2 = ces_23_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_18_io_ins_3 = ces_22_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_19_clock = clock;
  assign ces_22_19_io_ins_0 = ces_21_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_19_io_ins_1 = ces_22_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_19_io_ins_2 = ces_23_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_19_io_ins_3 = ces_22_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_20_clock = clock;
  assign ces_22_20_io_ins_0 = ces_21_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_20_io_ins_1 = ces_22_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_20_io_ins_2 = ces_23_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_20_io_ins_3 = ces_22_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_21_clock = clock;
  assign ces_22_21_io_ins_0 = ces_21_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_21_io_ins_1 = ces_22_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_21_io_ins_2 = ces_23_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_21_io_ins_3 = ces_22_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_22_clock = clock;
  assign ces_22_22_io_ins_0 = ces_21_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_22_io_ins_1 = ces_22_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_22_io_ins_2 = ces_23_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_22_io_ins_3 = ces_22_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_23_clock = clock;
  assign ces_22_23_io_ins_0 = ces_21_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_23_io_ins_1 = ces_22_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_23_io_ins_2 = ces_23_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_23_io_ins_3 = ces_22_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_24_clock = clock;
  assign ces_22_24_io_ins_0 = ces_21_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_24_io_ins_1 = ces_22_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_24_io_ins_2 = ces_23_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_24_io_ins_3 = ces_22_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_25_clock = clock;
  assign ces_22_25_io_ins_0 = ces_21_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_25_io_ins_1 = ces_22_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_25_io_ins_2 = ces_23_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_25_io_ins_3 = ces_22_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_26_clock = clock;
  assign ces_22_26_io_ins_0 = ces_21_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_26_io_ins_1 = ces_22_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_26_io_ins_2 = ces_23_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_26_io_ins_3 = ces_22_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_27_clock = clock;
  assign ces_22_27_io_ins_0 = ces_21_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_27_io_ins_1 = ces_22_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_27_io_ins_2 = ces_23_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_27_io_ins_3 = ces_22_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_28_clock = clock;
  assign ces_22_28_io_ins_0 = ces_21_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_28_io_ins_1 = ces_22_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_28_io_ins_2 = ces_23_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_28_io_ins_3 = ces_22_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_29_clock = clock;
  assign ces_22_29_io_ins_0 = ces_21_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_29_io_ins_1 = ces_22_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_29_io_ins_2 = ces_23_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_29_io_ins_3 = ces_22_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_30_clock = clock;
  assign ces_22_30_io_ins_0 = ces_21_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_30_io_ins_1 = ces_22_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_22_30_io_ins_2 = ces_23_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_30_io_ins_3 = ces_22_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_22_31_clock = clock;
  assign ces_22_31_io_ins_0 = ces_21_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_31_io_ins_1 = io_insVertical_0_22; // @[MockArray.scala 45:87]
  assign ces_22_31_io_ins_2 = ces_23_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_31_io_ins_3 = ces_22_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_0_clock = clock;
  assign ces_23_0_io_ins_0 = ces_22_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_0_io_ins_1 = ces_23_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_0_io_ins_2 = ces_24_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_0_io_ins_3 = io_insVertical_1_23; // @[MockArray.scala 47:87]
  assign ces_23_1_clock = clock;
  assign ces_23_1_io_ins_0 = ces_22_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_1_io_ins_1 = ces_23_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_1_io_ins_2 = ces_24_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_1_io_ins_3 = ces_23_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_2_clock = clock;
  assign ces_23_2_io_ins_0 = ces_22_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_2_io_ins_1 = ces_23_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_2_io_ins_2 = ces_24_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_2_io_ins_3 = ces_23_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_3_clock = clock;
  assign ces_23_3_io_ins_0 = ces_22_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_3_io_ins_1 = ces_23_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_3_io_ins_2 = ces_24_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_3_io_ins_3 = ces_23_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_4_clock = clock;
  assign ces_23_4_io_ins_0 = ces_22_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_4_io_ins_1 = ces_23_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_4_io_ins_2 = ces_24_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_4_io_ins_3 = ces_23_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_5_clock = clock;
  assign ces_23_5_io_ins_0 = ces_22_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_5_io_ins_1 = ces_23_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_5_io_ins_2 = ces_24_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_5_io_ins_3 = ces_23_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_6_clock = clock;
  assign ces_23_6_io_ins_0 = ces_22_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_6_io_ins_1 = ces_23_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_6_io_ins_2 = ces_24_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_6_io_ins_3 = ces_23_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_7_clock = clock;
  assign ces_23_7_io_ins_0 = ces_22_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_7_io_ins_1 = ces_23_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_7_io_ins_2 = ces_24_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_7_io_ins_3 = ces_23_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_8_clock = clock;
  assign ces_23_8_io_ins_0 = ces_22_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_8_io_ins_1 = ces_23_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_8_io_ins_2 = ces_24_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_8_io_ins_3 = ces_23_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_9_clock = clock;
  assign ces_23_9_io_ins_0 = ces_22_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_9_io_ins_1 = ces_23_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_9_io_ins_2 = ces_24_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_9_io_ins_3 = ces_23_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_10_clock = clock;
  assign ces_23_10_io_ins_0 = ces_22_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_10_io_ins_1 = ces_23_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_10_io_ins_2 = ces_24_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_10_io_ins_3 = ces_23_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_11_clock = clock;
  assign ces_23_11_io_ins_0 = ces_22_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_11_io_ins_1 = ces_23_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_11_io_ins_2 = ces_24_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_11_io_ins_3 = ces_23_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_12_clock = clock;
  assign ces_23_12_io_ins_0 = ces_22_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_12_io_ins_1 = ces_23_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_12_io_ins_2 = ces_24_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_12_io_ins_3 = ces_23_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_13_clock = clock;
  assign ces_23_13_io_ins_0 = ces_22_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_13_io_ins_1 = ces_23_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_13_io_ins_2 = ces_24_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_13_io_ins_3 = ces_23_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_14_clock = clock;
  assign ces_23_14_io_ins_0 = ces_22_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_14_io_ins_1 = ces_23_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_14_io_ins_2 = ces_24_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_14_io_ins_3 = ces_23_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_15_clock = clock;
  assign ces_23_15_io_ins_0 = ces_22_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_15_io_ins_1 = ces_23_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_15_io_ins_2 = ces_24_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_15_io_ins_3 = ces_23_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_16_clock = clock;
  assign ces_23_16_io_ins_0 = ces_22_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_16_io_ins_1 = ces_23_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_16_io_ins_2 = ces_24_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_16_io_ins_3 = ces_23_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_17_clock = clock;
  assign ces_23_17_io_ins_0 = ces_22_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_17_io_ins_1 = ces_23_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_17_io_ins_2 = ces_24_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_17_io_ins_3 = ces_23_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_18_clock = clock;
  assign ces_23_18_io_ins_0 = ces_22_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_18_io_ins_1 = ces_23_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_18_io_ins_2 = ces_24_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_18_io_ins_3 = ces_23_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_19_clock = clock;
  assign ces_23_19_io_ins_0 = ces_22_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_19_io_ins_1 = ces_23_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_19_io_ins_2 = ces_24_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_19_io_ins_3 = ces_23_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_20_clock = clock;
  assign ces_23_20_io_ins_0 = ces_22_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_20_io_ins_1 = ces_23_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_20_io_ins_2 = ces_24_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_20_io_ins_3 = ces_23_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_21_clock = clock;
  assign ces_23_21_io_ins_0 = ces_22_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_21_io_ins_1 = ces_23_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_21_io_ins_2 = ces_24_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_21_io_ins_3 = ces_23_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_22_clock = clock;
  assign ces_23_22_io_ins_0 = ces_22_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_22_io_ins_1 = ces_23_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_22_io_ins_2 = ces_24_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_22_io_ins_3 = ces_23_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_23_clock = clock;
  assign ces_23_23_io_ins_0 = ces_22_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_23_io_ins_1 = ces_23_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_23_io_ins_2 = ces_24_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_23_io_ins_3 = ces_23_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_24_clock = clock;
  assign ces_23_24_io_ins_0 = ces_22_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_24_io_ins_1 = ces_23_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_24_io_ins_2 = ces_24_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_24_io_ins_3 = ces_23_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_25_clock = clock;
  assign ces_23_25_io_ins_0 = ces_22_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_25_io_ins_1 = ces_23_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_25_io_ins_2 = ces_24_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_25_io_ins_3 = ces_23_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_26_clock = clock;
  assign ces_23_26_io_ins_0 = ces_22_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_26_io_ins_1 = ces_23_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_26_io_ins_2 = ces_24_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_26_io_ins_3 = ces_23_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_27_clock = clock;
  assign ces_23_27_io_ins_0 = ces_22_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_27_io_ins_1 = ces_23_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_27_io_ins_2 = ces_24_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_27_io_ins_3 = ces_23_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_28_clock = clock;
  assign ces_23_28_io_ins_0 = ces_22_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_28_io_ins_1 = ces_23_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_28_io_ins_2 = ces_24_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_28_io_ins_3 = ces_23_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_29_clock = clock;
  assign ces_23_29_io_ins_0 = ces_22_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_29_io_ins_1 = ces_23_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_29_io_ins_2 = ces_24_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_29_io_ins_3 = ces_23_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_30_clock = clock;
  assign ces_23_30_io_ins_0 = ces_22_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_30_io_ins_1 = ces_23_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_23_30_io_ins_2 = ces_24_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_30_io_ins_3 = ces_23_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_23_31_clock = clock;
  assign ces_23_31_io_ins_0 = ces_22_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_31_io_ins_1 = io_insVertical_0_23; // @[MockArray.scala 45:87]
  assign ces_23_31_io_ins_2 = ces_24_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_31_io_ins_3 = ces_23_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_0_clock = clock;
  assign ces_24_0_io_ins_0 = ces_23_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_0_io_ins_1 = ces_24_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_0_io_ins_2 = ces_25_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_0_io_ins_3 = io_insVertical_1_24; // @[MockArray.scala 47:87]
  assign ces_24_1_clock = clock;
  assign ces_24_1_io_ins_0 = ces_23_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_1_io_ins_1 = ces_24_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_1_io_ins_2 = ces_25_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_1_io_ins_3 = ces_24_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_2_clock = clock;
  assign ces_24_2_io_ins_0 = ces_23_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_2_io_ins_1 = ces_24_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_2_io_ins_2 = ces_25_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_2_io_ins_3 = ces_24_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_3_clock = clock;
  assign ces_24_3_io_ins_0 = ces_23_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_3_io_ins_1 = ces_24_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_3_io_ins_2 = ces_25_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_3_io_ins_3 = ces_24_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_4_clock = clock;
  assign ces_24_4_io_ins_0 = ces_23_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_4_io_ins_1 = ces_24_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_4_io_ins_2 = ces_25_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_4_io_ins_3 = ces_24_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_5_clock = clock;
  assign ces_24_5_io_ins_0 = ces_23_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_5_io_ins_1 = ces_24_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_5_io_ins_2 = ces_25_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_5_io_ins_3 = ces_24_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_6_clock = clock;
  assign ces_24_6_io_ins_0 = ces_23_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_6_io_ins_1 = ces_24_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_6_io_ins_2 = ces_25_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_6_io_ins_3 = ces_24_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_7_clock = clock;
  assign ces_24_7_io_ins_0 = ces_23_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_7_io_ins_1 = ces_24_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_7_io_ins_2 = ces_25_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_7_io_ins_3 = ces_24_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_8_clock = clock;
  assign ces_24_8_io_ins_0 = ces_23_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_8_io_ins_1 = ces_24_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_8_io_ins_2 = ces_25_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_8_io_ins_3 = ces_24_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_9_clock = clock;
  assign ces_24_9_io_ins_0 = ces_23_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_9_io_ins_1 = ces_24_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_9_io_ins_2 = ces_25_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_9_io_ins_3 = ces_24_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_10_clock = clock;
  assign ces_24_10_io_ins_0 = ces_23_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_10_io_ins_1 = ces_24_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_10_io_ins_2 = ces_25_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_10_io_ins_3 = ces_24_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_11_clock = clock;
  assign ces_24_11_io_ins_0 = ces_23_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_11_io_ins_1 = ces_24_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_11_io_ins_2 = ces_25_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_11_io_ins_3 = ces_24_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_12_clock = clock;
  assign ces_24_12_io_ins_0 = ces_23_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_12_io_ins_1 = ces_24_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_12_io_ins_2 = ces_25_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_12_io_ins_3 = ces_24_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_13_clock = clock;
  assign ces_24_13_io_ins_0 = ces_23_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_13_io_ins_1 = ces_24_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_13_io_ins_2 = ces_25_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_13_io_ins_3 = ces_24_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_14_clock = clock;
  assign ces_24_14_io_ins_0 = ces_23_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_14_io_ins_1 = ces_24_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_14_io_ins_2 = ces_25_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_14_io_ins_3 = ces_24_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_15_clock = clock;
  assign ces_24_15_io_ins_0 = ces_23_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_15_io_ins_1 = ces_24_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_15_io_ins_2 = ces_25_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_15_io_ins_3 = ces_24_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_16_clock = clock;
  assign ces_24_16_io_ins_0 = ces_23_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_16_io_ins_1 = ces_24_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_16_io_ins_2 = ces_25_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_16_io_ins_3 = ces_24_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_17_clock = clock;
  assign ces_24_17_io_ins_0 = ces_23_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_17_io_ins_1 = ces_24_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_17_io_ins_2 = ces_25_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_17_io_ins_3 = ces_24_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_18_clock = clock;
  assign ces_24_18_io_ins_0 = ces_23_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_18_io_ins_1 = ces_24_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_18_io_ins_2 = ces_25_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_18_io_ins_3 = ces_24_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_19_clock = clock;
  assign ces_24_19_io_ins_0 = ces_23_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_19_io_ins_1 = ces_24_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_19_io_ins_2 = ces_25_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_19_io_ins_3 = ces_24_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_20_clock = clock;
  assign ces_24_20_io_ins_0 = ces_23_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_20_io_ins_1 = ces_24_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_20_io_ins_2 = ces_25_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_20_io_ins_3 = ces_24_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_21_clock = clock;
  assign ces_24_21_io_ins_0 = ces_23_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_21_io_ins_1 = ces_24_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_21_io_ins_2 = ces_25_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_21_io_ins_3 = ces_24_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_22_clock = clock;
  assign ces_24_22_io_ins_0 = ces_23_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_22_io_ins_1 = ces_24_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_22_io_ins_2 = ces_25_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_22_io_ins_3 = ces_24_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_23_clock = clock;
  assign ces_24_23_io_ins_0 = ces_23_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_23_io_ins_1 = ces_24_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_23_io_ins_2 = ces_25_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_23_io_ins_3 = ces_24_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_24_clock = clock;
  assign ces_24_24_io_ins_0 = ces_23_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_24_io_ins_1 = ces_24_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_24_io_ins_2 = ces_25_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_24_io_ins_3 = ces_24_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_25_clock = clock;
  assign ces_24_25_io_ins_0 = ces_23_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_25_io_ins_1 = ces_24_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_25_io_ins_2 = ces_25_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_25_io_ins_3 = ces_24_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_26_clock = clock;
  assign ces_24_26_io_ins_0 = ces_23_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_26_io_ins_1 = ces_24_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_26_io_ins_2 = ces_25_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_26_io_ins_3 = ces_24_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_27_clock = clock;
  assign ces_24_27_io_ins_0 = ces_23_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_27_io_ins_1 = ces_24_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_27_io_ins_2 = ces_25_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_27_io_ins_3 = ces_24_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_28_clock = clock;
  assign ces_24_28_io_ins_0 = ces_23_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_28_io_ins_1 = ces_24_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_28_io_ins_2 = ces_25_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_28_io_ins_3 = ces_24_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_29_clock = clock;
  assign ces_24_29_io_ins_0 = ces_23_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_29_io_ins_1 = ces_24_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_29_io_ins_2 = ces_25_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_29_io_ins_3 = ces_24_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_30_clock = clock;
  assign ces_24_30_io_ins_0 = ces_23_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_30_io_ins_1 = ces_24_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_24_30_io_ins_2 = ces_25_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_30_io_ins_3 = ces_24_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_24_31_clock = clock;
  assign ces_24_31_io_ins_0 = ces_23_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_31_io_ins_1 = io_insVertical_0_24; // @[MockArray.scala 45:87]
  assign ces_24_31_io_ins_2 = ces_25_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_31_io_ins_3 = ces_24_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_0_clock = clock;
  assign ces_25_0_io_ins_0 = ces_24_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_0_io_ins_1 = ces_25_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_0_io_ins_2 = ces_26_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_0_io_ins_3 = io_insVertical_1_25; // @[MockArray.scala 47:87]
  assign ces_25_1_clock = clock;
  assign ces_25_1_io_ins_0 = ces_24_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_1_io_ins_1 = ces_25_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_1_io_ins_2 = ces_26_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_1_io_ins_3 = ces_25_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_2_clock = clock;
  assign ces_25_2_io_ins_0 = ces_24_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_2_io_ins_1 = ces_25_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_2_io_ins_2 = ces_26_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_2_io_ins_3 = ces_25_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_3_clock = clock;
  assign ces_25_3_io_ins_0 = ces_24_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_3_io_ins_1 = ces_25_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_3_io_ins_2 = ces_26_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_3_io_ins_3 = ces_25_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_4_clock = clock;
  assign ces_25_4_io_ins_0 = ces_24_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_4_io_ins_1 = ces_25_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_4_io_ins_2 = ces_26_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_4_io_ins_3 = ces_25_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_5_clock = clock;
  assign ces_25_5_io_ins_0 = ces_24_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_5_io_ins_1 = ces_25_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_5_io_ins_2 = ces_26_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_5_io_ins_3 = ces_25_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_6_clock = clock;
  assign ces_25_6_io_ins_0 = ces_24_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_6_io_ins_1 = ces_25_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_6_io_ins_2 = ces_26_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_6_io_ins_3 = ces_25_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_7_clock = clock;
  assign ces_25_7_io_ins_0 = ces_24_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_7_io_ins_1 = ces_25_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_7_io_ins_2 = ces_26_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_7_io_ins_3 = ces_25_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_8_clock = clock;
  assign ces_25_8_io_ins_0 = ces_24_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_8_io_ins_1 = ces_25_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_8_io_ins_2 = ces_26_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_8_io_ins_3 = ces_25_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_9_clock = clock;
  assign ces_25_9_io_ins_0 = ces_24_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_9_io_ins_1 = ces_25_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_9_io_ins_2 = ces_26_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_9_io_ins_3 = ces_25_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_10_clock = clock;
  assign ces_25_10_io_ins_0 = ces_24_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_10_io_ins_1 = ces_25_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_10_io_ins_2 = ces_26_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_10_io_ins_3 = ces_25_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_11_clock = clock;
  assign ces_25_11_io_ins_0 = ces_24_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_11_io_ins_1 = ces_25_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_11_io_ins_2 = ces_26_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_11_io_ins_3 = ces_25_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_12_clock = clock;
  assign ces_25_12_io_ins_0 = ces_24_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_12_io_ins_1 = ces_25_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_12_io_ins_2 = ces_26_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_12_io_ins_3 = ces_25_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_13_clock = clock;
  assign ces_25_13_io_ins_0 = ces_24_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_13_io_ins_1 = ces_25_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_13_io_ins_2 = ces_26_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_13_io_ins_3 = ces_25_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_14_clock = clock;
  assign ces_25_14_io_ins_0 = ces_24_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_14_io_ins_1 = ces_25_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_14_io_ins_2 = ces_26_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_14_io_ins_3 = ces_25_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_15_clock = clock;
  assign ces_25_15_io_ins_0 = ces_24_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_15_io_ins_1 = ces_25_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_15_io_ins_2 = ces_26_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_15_io_ins_3 = ces_25_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_16_clock = clock;
  assign ces_25_16_io_ins_0 = ces_24_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_16_io_ins_1 = ces_25_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_16_io_ins_2 = ces_26_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_16_io_ins_3 = ces_25_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_17_clock = clock;
  assign ces_25_17_io_ins_0 = ces_24_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_17_io_ins_1 = ces_25_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_17_io_ins_2 = ces_26_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_17_io_ins_3 = ces_25_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_18_clock = clock;
  assign ces_25_18_io_ins_0 = ces_24_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_18_io_ins_1 = ces_25_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_18_io_ins_2 = ces_26_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_18_io_ins_3 = ces_25_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_19_clock = clock;
  assign ces_25_19_io_ins_0 = ces_24_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_19_io_ins_1 = ces_25_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_19_io_ins_2 = ces_26_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_19_io_ins_3 = ces_25_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_20_clock = clock;
  assign ces_25_20_io_ins_0 = ces_24_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_20_io_ins_1 = ces_25_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_20_io_ins_2 = ces_26_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_20_io_ins_3 = ces_25_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_21_clock = clock;
  assign ces_25_21_io_ins_0 = ces_24_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_21_io_ins_1 = ces_25_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_21_io_ins_2 = ces_26_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_21_io_ins_3 = ces_25_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_22_clock = clock;
  assign ces_25_22_io_ins_0 = ces_24_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_22_io_ins_1 = ces_25_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_22_io_ins_2 = ces_26_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_22_io_ins_3 = ces_25_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_23_clock = clock;
  assign ces_25_23_io_ins_0 = ces_24_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_23_io_ins_1 = ces_25_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_23_io_ins_2 = ces_26_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_23_io_ins_3 = ces_25_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_24_clock = clock;
  assign ces_25_24_io_ins_0 = ces_24_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_24_io_ins_1 = ces_25_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_24_io_ins_2 = ces_26_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_24_io_ins_3 = ces_25_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_25_clock = clock;
  assign ces_25_25_io_ins_0 = ces_24_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_25_io_ins_1 = ces_25_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_25_io_ins_2 = ces_26_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_25_io_ins_3 = ces_25_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_26_clock = clock;
  assign ces_25_26_io_ins_0 = ces_24_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_26_io_ins_1 = ces_25_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_26_io_ins_2 = ces_26_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_26_io_ins_3 = ces_25_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_27_clock = clock;
  assign ces_25_27_io_ins_0 = ces_24_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_27_io_ins_1 = ces_25_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_27_io_ins_2 = ces_26_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_27_io_ins_3 = ces_25_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_28_clock = clock;
  assign ces_25_28_io_ins_0 = ces_24_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_28_io_ins_1 = ces_25_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_28_io_ins_2 = ces_26_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_28_io_ins_3 = ces_25_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_29_clock = clock;
  assign ces_25_29_io_ins_0 = ces_24_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_29_io_ins_1 = ces_25_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_29_io_ins_2 = ces_26_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_29_io_ins_3 = ces_25_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_30_clock = clock;
  assign ces_25_30_io_ins_0 = ces_24_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_30_io_ins_1 = ces_25_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_25_30_io_ins_2 = ces_26_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_30_io_ins_3 = ces_25_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_25_31_clock = clock;
  assign ces_25_31_io_ins_0 = ces_24_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_31_io_ins_1 = io_insVertical_0_25; // @[MockArray.scala 45:87]
  assign ces_25_31_io_ins_2 = ces_26_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_31_io_ins_3 = ces_25_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_0_clock = clock;
  assign ces_26_0_io_ins_0 = ces_25_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_0_io_ins_1 = ces_26_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_0_io_ins_2 = ces_27_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_0_io_ins_3 = io_insVertical_1_26; // @[MockArray.scala 47:87]
  assign ces_26_1_clock = clock;
  assign ces_26_1_io_ins_0 = ces_25_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_1_io_ins_1 = ces_26_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_1_io_ins_2 = ces_27_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_1_io_ins_3 = ces_26_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_2_clock = clock;
  assign ces_26_2_io_ins_0 = ces_25_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_2_io_ins_1 = ces_26_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_2_io_ins_2 = ces_27_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_2_io_ins_3 = ces_26_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_3_clock = clock;
  assign ces_26_3_io_ins_0 = ces_25_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_3_io_ins_1 = ces_26_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_3_io_ins_2 = ces_27_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_3_io_ins_3 = ces_26_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_4_clock = clock;
  assign ces_26_4_io_ins_0 = ces_25_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_4_io_ins_1 = ces_26_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_4_io_ins_2 = ces_27_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_4_io_ins_3 = ces_26_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_5_clock = clock;
  assign ces_26_5_io_ins_0 = ces_25_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_5_io_ins_1 = ces_26_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_5_io_ins_2 = ces_27_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_5_io_ins_3 = ces_26_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_6_clock = clock;
  assign ces_26_6_io_ins_0 = ces_25_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_6_io_ins_1 = ces_26_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_6_io_ins_2 = ces_27_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_6_io_ins_3 = ces_26_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_7_clock = clock;
  assign ces_26_7_io_ins_0 = ces_25_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_7_io_ins_1 = ces_26_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_7_io_ins_2 = ces_27_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_7_io_ins_3 = ces_26_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_8_clock = clock;
  assign ces_26_8_io_ins_0 = ces_25_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_8_io_ins_1 = ces_26_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_8_io_ins_2 = ces_27_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_8_io_ins_3 = ces_26_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_9_clock = clock;
  assign ces_26_9_io_ins_0 = ces_25_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_9_io_ins_1 = ces_26_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_9_io_ins_2 = ces_27_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_9_io_ins_3 = ces_26_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_10_clock = clock;
  assign ces_26_10_io_ins_0 = ces_25_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_10_io_ins_1 = ces_26_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_10_io_ins_2 = ces_27_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_10_io_ins_3 = ces_26_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_11_clock = clock;
  assign ces_26_11_io_ins_0 = ces_25_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_11_io_ins_1 = ces_26_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_11_io_ins_2 = ces_27_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_11_io_ins_3 = ces_26_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_12_clock = clock;
  assign ces_26_12_io_ins_0 = ces_25_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_12_io_ins_1 = ces_26_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_12_io_ins_2 = ces_27_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_12_io_ins_3 = ces_26_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_13_clock = clock;
  assign ces_26_13_io_ins_0 = ces_25_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_13_io_ins_1 = ces_26_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_13_io_ins_2 = ces_27_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_13_io_ins_3 = ces_26_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_14_clock = clock;
  assign ces_26_14_io_ins_0 = ces_25_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_14_io_ins_1 = ces_26_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_14_io_ins_2 = ces_27_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_14_io_ins_3 = ces_26_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_15_clock = clock;
  assign ces_26_15_io_ins_0 = ces_25_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_15_io_ins_1 = ces_26_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_15_io_ins_2 = ces_27_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_15_io_ins_3 = ces_26_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_16_clock = clock;
  assign ces_26_16_io_ins_0 = ces_25_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_16_io_ins_1 = ces_26_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_16_io_ins_2 = ces_27_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_16_io_ins_3 = ces_26_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_17_clock = clock;
  assign ces_26_17_io_ins_0 = ces_25_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_17_io_ins_1 = ces_26_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_17_io_ins_2 = ces_27_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_17_io_ins_3 = ces_26_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_18_clock = clock;
  assign ces_26_18_io_ins_0 = ces_25_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_18_io_ins_1 = ces_26_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_18_io_ins_2 = ces_27_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_18_io_ins_3 = ces_26_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_19_clock = clock;
  assign ces_26_19_io_ins_0 = ces_25_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_19_io_ins_1 = ces_26_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_19_io_ins_2 = ces_27_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_19_io_ins_3 = ces_26_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_20_clock = clock;
  assign ces_26_20_io_ins_0 = ces_25_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_20_io_ins_1 = ces_26_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_20_io_ins_2 = ces_27_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_20_io_ins_3 = ces_26_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_21_clock = clock;
  assign ces_26_21_io_ins_0 = ces_25_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_21_io_ins_1 = ces_26_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_21_io_ins_2 = ces_27_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_21_io_ins_3 = ces_26_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_22_clock = clock;
  assign ces_26_22_io_ins_0 = ces_25_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_22_io_ins_1 = ces_26_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_22_io_ins_2 = ces_27_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_22_io_ins_3 = ces_26_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_23_clock = clock;
  assign ces_26_23_io_ins_0 = ces_25_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_23_io_ins_1 = ces_26_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_23_io_ins_2 = ces_27_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_23_io_ins_3 = ces_26_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_24_clock = clock;
  assign ces_26_24_io_ins_0 = ces_25_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_24_io_ins_1 = ces_26_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_24_io_ins_2 = ces_27_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_24_io_ins_3 = ces_26_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_25_clock = clock;
  assign ces_26_25_io_ins_0 = ces_25_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_25_io_ins_1 = ces_26_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_25_io_ins_2 = ces_27_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_25_io_ins_3 = ces_26_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_26_clock = clock;
  assign ces_26_26_io_ins_0 = ces_25_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_26_io_ins_1 = ces_26_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_26_io_ins_2 = ces_27_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_26_io_ins_3 = ces_26_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_27_clock = clock;
  assign ces_26_27_io_ins_0 = ces_25_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_27_io_ins_1 = ces_26_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_27_io_ins_2 = ces_27_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_27_io_ins_3 = ces_26_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_28_clock = clock;
  assign ces_26_28_io_ins_0 = ces_25_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_28_io_ins_1 = ces_26_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_28_io_ins_2 = ces_27_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_28_io_ins_3 = ces_26_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_29_clock = clock;
  assign ces_26_29_io_ins_0 = ces_25_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_29_io_ins_1 = ces_26_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_29_io_ins_2 = ces_27_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_29_io_ins_3 = ces_26_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_30_clock = clock;
  assign ces_26_30_io_ins_0 = ces_25_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_30_io_ins_1 = ces_26_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_26_30_io_ins_2 = ces_27_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_30_io_ins_3 = ces_26_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_26_31_clock = clock;
  assign ces_26_31_io_ins_0 = ces_25_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_31_io_ins_1 = io_insVertical_0_26; // @[MockArray.scala 45:87]
  assign ces_26_31_io_ins_2 = ces_27_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_31_io_ins_3 = ces_26_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_0_clock = clock;
  assign ces_27_0_io_ins_0 = ces_26_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_0_io_ins_1 = ces_27_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_0_io_ins_2 = ces_28_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_0_io_ins_3 = io_insVertical_1_27; // @[MockArray.scala 47:87]
  assign ces_27_1_clock = clock;
  assign ces_27_1_io_ins_0 = ces_26_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_1_io_ins_1 = ces_27_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_1_io_ins_2 = ces_28_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_1_io_ins_3 = ces_27_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_2_clock = clock;
  assign ces_27_2_io_ins_0 = ces_26_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_2_io_ins_1 = ces_27_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_2_io_ins_2 = ces_28_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_2_io_ins_3 = ces_27_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_3_clock = clock;
  assign ces_27_3_io_ins_0 = ces_26_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_3_io_ins_1 = ces_27_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_3_io_ins_2 = ces_28_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_3_io_ins_3 = ces_27_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_4_clock = clock;
  assign ces_27_4_io_ins_0 = ces_26_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_4_io_ins_1 = ces_27_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_4_io_ins_2 = ces_28_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_4_io_ins_3 = ces_27_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_5_clock = clock;
  assign ces_27_5_io_ins_0 = ces_26_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_5_io_ins_1 = ces_27_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_5_io_ins_2 = ces_28_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_5_io_ins_3 = ces_27_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_6_clock = clock;
  assign ces_27_6_io_ins_0 = ces_26_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_6_io_ins_1 = ces_27_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_6_io_ins_2 = ces_28_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_6_io_ins_3 = ces_27_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_7_clock = clock;
  assign ces_27_7_io_ins_0 = ces_26_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_7_io_ins_1 = ces_27_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_7_io_ins_2 = ces_28_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_7_io_ins_3 = ces_27_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_8_clock = clock;
  assign ces_27_8_io_ins_0 = ces_26_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_8_io_ins_1 = ces_27_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_8_io_ins_2 = ces_28_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_8_io_ins_3 = ces_27_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_9_clock = clock;
  assign ces_27_9_io_ins_0 = ces_26_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_9_io_ins_1 = ces_27_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_9_io_ins_2 = ces_28_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_9_io_ins_3 = ces_27_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_10_clock = clock;
  assign ces_27_10_io_ins_0 = ces_26_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_10_io_ins_1 = ces_27_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_10_io_ins_2 = ces_28_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_10_io_ins_3 = ces_27_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_11_clock = clock;
  assign ces_27_11_io_ins_0 = ces_26_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_11_io_ins_1 = ces_27_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_11_io_ins_2 = ces_28_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_11_io_ins_3 = ces_27_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_12_clock = clock;
  assign ces_27_12_io_ins_0 = ces_26_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_12_io_ins_1 = ces_27_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_12_io_ins_2 = ces_28_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_12_io_ins_3 = ces_27_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_13_clock = clock;
  assign ces_27_13_io_ins_0 = ces_26_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_13_io_ins_1 = ces_27_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_13_io_ins_2 = ces_28_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_13_io_ins_3 = ces_27_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_14_clock = clock;
  assign ces_27_14_io_ins_0 = ces_26_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_14_io_ins_1 = ces_27_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_14_io_ins_2 = ces_28_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_14_io_ins_3 = ces_27_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_15_clock = clock;
  assign ces_27_15_io_ins_0 = ces_26_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_15_io_ins_1 = ces_27_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_15_io_ins_2 = ces_28_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_15_io_ins_3 = ces_27_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_16_clock = clock;
  assign ces_27_16_io_ins_0 = ces_26_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_16_io_ins_1 = ces_27_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_16_io_ins_2 = ces_28_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_16_io_ins_3 = ces_27_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_17_clock = clock;
  assign ces_27_17_io_ins_0 = ces_26_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_17_io_ins_1 = ces_27_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_17_io_ins_2 = ces_28_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_17_io_ins_3 = ces_27_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_18_clock = clock;
  assign ces_27_18_io_ins_0 = ces_26_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_18_io_ins_1 = ces_27_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_18_io_ins_2 = ces_28_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_18_io_ins_3 = ces_27_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_19_clock = clock;
  assign ces_27_19_io_ins_0 = ces_26_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_19_io_ins_1 = ces_27_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_19_io_ins_2 = ces_28_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_19_io_ins_3 = ces_27_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_20_clock = clock;
  assign ces_27_20_io_ins_0 = ces_26_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_20_io_ins_1 = ces_27_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_20_io_ins_2 = ces_28_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_20_io_ins_3 = ces_27_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_21_clock = clock;
  assign ces_27_21_io_ins_0 = ces_26_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_21_io_ins_1 = ces_27_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_21_io_ins_2 = ces_28_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_21_io_ins_3 = ces_27_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_22_clock = clock;
  assign ces_27_22_io_ins_0 = ces_26_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_22_io_ins_1 = ces_27_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_22_io_ins_2 = ces_28_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_22_io_ins_3 = ces_27_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_23_clock = clock;
  assign ces_27_23_io_ins_0 = ces_26_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_23_io_ins_1 = ces_27_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_23_io_ins_2 = ces_28_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_23_io_ins_3 = ces_27_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_24_clock = clock;
  assign ces_27_24_io_ins_0 = ces_26_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_24_io_ins_1 = ces_27_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_24_io_ins_2 = ces_28_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_24_io_ins_3 = ces_27_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_25_clock = clock;
  assign ces_27_25_io_ins_0 = ces_26_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_25_io_ins_1 = ces_27_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_25_io_ins_2 = ces_28_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_25_io_ins_3 = ces_27_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_26_clock = clock;
  assign ces_27_26_io_ins_0 = ces_26_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_26_io_ins_1 = ces_27_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_26_io_ins_2 = ces_28_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_26_io_ins_3 = ces_27_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_27_clock = clock;
  assign ces_27_27_io_ins_0 = ces_26_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_27_io_ins_1 = ces_27_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_27_io_ins_2 = ces_28_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_27_io_ins_3 = ces_27_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_28_clock = clock;
  assign ces_27_28_io_ins_0 = ces_26_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_28_io_ins_1 = ces_27_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_28_io_ins_2 = ces_28_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_28_io_ins_3 = ces_27_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_29_clock = clock;
  assign ces_27_29_io_ins_0 = ces_26_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_29_io_ins_1 = ces_27_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_29_io_ins_2 = ces_28_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_29_io_ins_3 = ces_27_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_30_clock = clock;
  assign ces_27_30_io_ins_0 = ces_26_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_30_io_ins_1 = ces_27_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_27_30_io_ins_2 = ces_28_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_30_io_ins_3 = ces_27_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_27_31_clock = clock;
  assign ces_27_31_io_ins_0 = ces_26_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_31_io_ins_1 = io_insVertical_0_27; // @[MockArray.scala 45:87]
  assign ces_27_31_io_ins_2 = ces_28_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_31_io_ins_3 = ces_27_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_0_clock = clock;
  assign ces_28_0_io_ins_0 = ces_27_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_0_io_ins_1 = ces_28_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_0_io_ins_2 = ces_29_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_0_io_ins_3 = io_insVertical_1_28; // @[MockArray.scala 47:87]
  assign ces_28_1_clock = clock;
  assign ces_28_1_io_ins_0 = ces_27_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_1_io_ins_1 = ces_28_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_1_io_ins_2 = ces_29_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_1_io_ins_3 = ces_28_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_2_clock = clock;
  assign ces_28_2_io_ins_0 = ces_27_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_2_io_ins_1 = ces_28_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_2_io_ins_2 = ces_29_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_2_io_ins_3 = ces_28_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_3_clock = clock;
  assign ces_28_3_io_ins_0 = ces_27_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_3_io_ins_1 = ces_28_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_3_io_ins_2 = ces_29_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_3_io_ins_3 = ces_28_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_4_clock = clock;
  assign ces_28_4_io_ins_0 = ces_27_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_4_io_ins_1 = ces_28_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_4_io_ins_2 = ces_29_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_4_io_ins_3 = ces_28_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_5_clock = clock;
  assign ces_28_5_io_ins_0 = ces_27_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_5_io_ins_1 = ces_28_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_5_io_ins_2 = ces_29_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_5_io_ins_3 = ces_28_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_6_clock = clock;
  assign ces_28_6_io_ins_0 = ces_27_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_6_io_ins_1 = ces_28_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_6_io_ins_2 = ces_29_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_6_io_ins_3 = ces_28_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_7_clock = clock;
  assign ces_28_7_io_ins_0 = ces_27_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_7_io_ins_1 = ces_28_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_7_io_ins_2 = ces_29_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_7_io_ins_3 = ces_28_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_8_clock = clock;
  assign ces_28_8_io_ins_0 = ces_27_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_8_io_ins_1 = ces_28_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_8_io_ins_2 = ces_29_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_8_io_ins_3 = ces_28_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_9_clock = clock;
  assign ces_28_9_io_ins_0 = ces_27_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_9_io_ins_1 = ces_28_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_9_io_ins_2 = ces_29_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_9_io_ins_3 = ces_28_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_10_clock = clock;
  assign ces_28_10_io_ins_0 = ces_27_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_10_io_ins_1 = ces_28_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_10_io_ins_2 = ces_29_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_10_io_ins_3 = ces_28_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_11_clock = clock;
  assign ces_28_11_io_ins_0 = ces_27_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_11_io_ins_1 = ces_28_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_11_io_ins_2 = ces_29_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_11_io_ins_3 = ces_28_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_12_clock = clock;
  assign ces_28_12_io_ins_0 = ces_27_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_12_io_ins_1 = ces_28_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_12_io_ins_2 = ces_29_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_12_io_ins_3 = ces_28_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_13_clock = clock;
  assign ces_28_13_io_ins_0 = ces_27_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_13_io_ins_1 = ces_28_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_13_io_ins_2 = ces_29_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_13_io_ins_3 = ces_28_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_14_clock = clock;
  assign ces_28_14_io_ins_0 = ces_27_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_14_io_ins_1 = ces_28_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_14_io_ins_2 = ces_29_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_14_io_ins_3 = ces_28_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_15_clock = clock;
  assign ces_28_15_io_ins_0 = ces_27_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_15_io_ins_1 = ces_28_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_15_io_ins_2 = ces_29_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_15_io_ins_3 = ces_28_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_16_clock = clock;
  assign ces_28_16_io_ins_0 = ces_27_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_16_io_ins_1 = ces_28_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_16_io_ins_2 = ces_29_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_16_io_ins_3 = ces_28_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_17_clock = clock;
  assign ces_28_17_io_ins_0 = ces_27_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_17_io_ins_1 = ces_28_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_17_io_ins_2 = ces_29_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_17_io_ins_3 = ces_28_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_18_clock = clock;
  assign ces_28_18_io_ins_0 = ces_27_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_18_io_ins_1 = ces_28_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_18_io_ins_2 = ces_29_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_18_io_ins_3 = ces_28_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_19_clock = clock;
  assign ces_28_19_io_ins_0 = ces_27_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_19_io_ins_1 = ces_28_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_19_io_ins_2 = ces_29_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_19_io_ins_3 = ces_28_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_20_clock = clock;
  assign ces_28_20_io_ins_0 = ces_27_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_20_io_ins_1 = ces_28_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_20_io_ins_2 = ces_29_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_20_io_ins_3 = ces_28_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_21_clock = clock;
  assign ces_28_21_io_ins_0 = ces_27_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_21_io_ins_1 = ces_28_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_21_io_ins_2 = ces_29_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_21_io_ins_3 = ces_28_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_22_clock = clock;
  assign ces_28_22_io_ins_0 = ces_27_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_22_io_ins_1 = ces_28_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_22_io_ins_2 = ces_29_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_22_io_ins_3 = ces_28_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_23_clock = clock;
  assign ces_28_23_io_ins_0 = ces_27_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_23_io_ins_1 = ces_28_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_23_io_ins_2 = ces_29_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_23_io_ins_3 = ces_28_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_24_clock = clock;
  assign ces_28_24_io_ins_0 = ces_27_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_24_io_ins_1 = ces_28_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_24_io_ins_2 = ces_29_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_24_io_ins_3 = ces_28_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_25_clock = clock;
  assign ces_28_25_io_ins_0 = ces_27_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_25_io_ins_1 = ces_28_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_25_io_ins_2 = ces_29_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_25_io_ins_3 = ces_28_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_26_clock = clock;
  assign ces_28_26_io_ins_0 = ces_27_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_26_io_ins_1 = ces_28_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_26_io_ins_2 = ces_29_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_26_io_ins_3 = ces_28_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_27_clock = clock;
  assign ces_28_27_io_ins_0 = ces_27_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_27_io_ins_1 = ces_28_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_27_io_ins_2 = ces_29_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_27_io_ins_3 = ces_28_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_28_clock = clock;
  assign ces_28_28_io_ins_0 = ces_27_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_28_io_ins_1 = ces_28_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_28_io_ins_2 = ces_29_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_28_io_ins_3 = ces_28_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_29_clock = clock;
  assign ces_28_29_io_ins_0 = ces_27_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_29_io_ins_1 = ces_28_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_29_io_ins_2 = ces_29_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_29_io_ins_3 = ces_28_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_30_clock = clock;
  assign ces_28_30_io_ins_0 = ces_27_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_30_io_ins_1 = ces_28_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_28_30_io_ins_2 = ces_29_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_30_io_ins_3 = ces_28_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_28_31_clock = clock;
  assign ces_28_31_io_ins_0 = ces_27_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_31_io_ins_1 = io_insVertical_0_28; // @[MockArray.scala 45:87]
  assign ces_28_31_io_ins_2 = ces_29_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_31_io_ins_3 = ces_28_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_0_clock = clock;
  assign ces_29_0_io_ins_0 = ces_28_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_0_io_ins_1 = ces_29_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_0_io_ins_2 = ces_30_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_0_io_ins_3 = io_insVertical_1_29; // @[MockArray.scala 47:87]
  assign ces_29_1_clock = clock;
  assign ces_29_1_io_ins_0 = ces_28_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_1_io_ins_1 = ces_29_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_1_io_ins_2 = ces_30_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_1_io_ins_3 = ces_29_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_2_clock = clock;
  assign ces_29_2_io_ins_0 = ces_28_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_2_io_ins_1 = ces_29_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_2_io_ins_2 = ces_30_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_2_io_ins_3 = ces_29_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_3_clock = clock;
  assign ces_29_3_io_ins_0 = ces_28_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_3_io_ins_1 = ces_29_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_3_io_ins_2 = ces_30_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_3_io_ins_3 = ces_29_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_4_clock = clock;
  assign ces_29_4_io_ins_0 = ces_28_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_4_io_ins_1 = ces_29_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_4_io_ins_2 = ces_30_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_4_io_ins_3 = ces_29_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_5_clock = clock;
  assign ces_29_5_io_ins_0 = ces_28_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_5_io_ins_1 = ces_29_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_5_io_ins_2 = ces_30_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_5_io_ins_3 = ces_29_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_6_clock = clock;
  assign ces_29_6_io_ins_0 = ces_28_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_6_io_ins_1 = ces_29_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_6_io_ins_2 = ces_30_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_6_io_ins_3 = ces_29_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_7_clock = clock;
  assign ces_29_7_io_ins_0 = ces_28_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_7_io_ins_1 = ces_29_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_7_io_ins_2 = ces_30_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_7_io_ins_3 = ces_29_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_8_clock = clock;
  assign ces_29_8_io_ins_0 = ces_28_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_8_io_ins_1 = ces_29_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_8_io_ins_2 = ces_30_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_8_io_ins_3 = ces_29_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_9_clock = clock;
  assign ces_29_9_io_ins_0 = ces_28_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_9_io_ins_1 = ces_29_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_9_io_ins_2 = ces_30_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_9_io_ins_3 = ces_29_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_10_clock = clock;
  assign ces_29_10_io_ins_0 = ces_28_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_10_io_ins_1 = ces_29_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_10_io_ins_2 = ces_30_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_10_io_ins_3 = ces_29_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_11_clock = clock;
  assign ces_29_11_io_ins_0 = ces_28_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_11_io_ins_1 = ces_29_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_11_io_ins_2 = ces_30_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_11_io_ins_3 = ces_29_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_12_clock = clock;
  assign ces_29_12_io_ins_0 = ces_28_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_12_io_ins_1 = ces_29_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_12_io_ins_2 = ces_30_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_12_io_ins_3 = ces_29_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_13_clock = clock;
  assign ces_29_13_io_ins_0 = ces_28_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_13_io_ins_1 = ces_29_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_13_io_ins_2 = ces_30_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_13_io_ins_3 = ces_29_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_14_clock = clock;
  assign ces_29_14_io_ins_0 = ces_28_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_14_io_ins_1 = ces_29_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_14_io_ins_2 = ces_30_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_14_io_ins_3 = ces_29_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_15_clock = clock;
  assign ces_29_15_io_ins_0 = ces_28_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_15_io_ins_1 = ces_29_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_15_io_ins_2 = ces_30_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_15_io_ins_3 = ces_29_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_16_clock = clock;
  assign ces_29_16_io_ins_0 = ces_28_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_16_io_ins_1 = ces_29_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_16_io_ins_2 = ces_30_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_16_io_ins_3 = ces_29_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_17_clock = clock;
  assign ces_29_17_io_ins_0 = ces_28_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_17_io_ins_1 = ces_29_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_17_io_ins_2 = ces_30_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_17_io_ins_3 = ces_29_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_18_clock = clock;
  assign ces_29_18_io_ins_0 = ces_28_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_18_io_ins_1 = ces_29_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_18_io_ins_2 = ces_30_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_18_io_ins_3 = ces_29_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_19_clock = clock;
  assign ces_29_19_io_ins_0 = ces_28_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_19_io_ins_1 = ces_29_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_19_io_ins_2 = ces_30_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_19_io_ins_3 = ces_29_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_20_clock = clock;
  assign ces_29_20_io_ins_0 = ces_28_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_20_io_ins_1 = ces_29_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_20_io_ins_2 = ces_30_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_20_io_ins_3 = ces_29_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_21_clock = clock;
  assign ces_29_21_io_ins_0 = ces_28_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_21_io_ins_1 = ces_29_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_21_io_ins_2 = ces_30_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_21_io_ins_3 = ces_29_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_22_clock = clock;
  assign ces_29_22_io_ins_0 = ces_28_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_22_io_ins_1 = ces_29_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_22_io_ins_2 = ces_30_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_22_io_ins_3 = ces_29_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_23_clock = clock;
  assign ces_29_23_io_ins_0 = ces_28_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_23_io_ins_1 = ces_29_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_23_io_ins_2 = ces_30_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_23_io_ins_3 = ces_29_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_24_clock = clock;
  assign ces_29_24_io_ins_0 = ces_28_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_24_io_ins_1 = ces_29_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_24_io_ins_2 = ces_30_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_24_io_ins_3 = ces_29_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_25_clock = clock;
  assign ces_29_25_io_ins_0 = ces_28_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_25_io_ins_1 = ces_29_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_25_io_ins_2 = ces_30_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_25_io_ins_3 = ces_29_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_26_clock = clock;
  assign ces_29_26_io_ins_0 = ces_28_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_26_io_ins_1 = ces_29_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_26_io_ins_2 = ces_30_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_26_io_ins_3 = ces_29_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_27_clock = clock;
  assign ces_29_27_io_ins_0 = ces_28_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_27_io_ins_1 = ces_29_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_27_io_ins_2 = ces_30_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_27_io_ins_3 = ces_29_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_28_clock = clock;
  assign ces_29_28_io_ins_0 = ces_28_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_28_io_ins_1 = ces_29_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_28_io_ins_2 = ces_30_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_28_io_ins_3 = ces_29_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_29_clock = clock;
  assign ces_29_29_io_ins_0 = ces_28_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_29_io_ins_1 = ces_29_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_29_io_ins_2 = ces_30_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_29_io_ins_3 = ces_29_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_30_clock = clock;
  assign ces_29_30_io_ins_0 = ces_28_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_30_io_ins_1 = ces_29_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_29_30_io_ins_2 = ces_30_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_30_io_ins_3 = ces_29_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_29_31_clock = clock;
  assign ces_29_31_io_ins_0 = ces_28_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_31_io_ins_1 = io_insVertical_0_29; // @[MockArray.scala 45:87]
  assign ces_29_31_io_ins_2 = ces_30_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_31_io_ins_3 = ces_29_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_0_clock = clock;
  assign ces_30_0_io_ins_0 = ces_29_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_0_io_ins_1 = ces_30_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_0_io_ins_2 = ces_31_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_0_io_ins_3 = io_insVertical_1_30; // @[MockArray.scala 47:87]
  assign ces_30_1_clock = clock;
  assign ces_30_1_io_ins_0 = ces_29_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_1_io_ins_1 = ces_30_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_1_io_ins_2 = ces_31_1_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_1_io_ins_3 = ces_30_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_2_clock = clock;
  assign ces_30_2_io_ins_0 = ces_29_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_2_io_ins_1 = ces_30_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_2_io_ins_2 = ces_31_2_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_2_io_ins_3 = ces_30_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_3_clock = clock;
  assign ces_30_3_io_ins_0 = ces_29_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_3_io_ins_1 = ces_30_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_3_io_ins_2 = ces_31_3_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_3_io_ins_3 = ces_30_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_4_clock = clock;
  assign ces_30_4_io_ins_0 = ces_29_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_4_io_ins_1 = ces_30_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_4_io_ins_2 = ces_31_4_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_4_io_ins_3 = ces_30_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_5_clock = clock;
  assign ces_30_5_io_ins_0 = ces_29_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_5_io_ins_1 = ces_30_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_5_io_ins_2 = ces_31_5_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_5_io_ins_3 = ces_30_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_6_clock = clock;
  assign ces_30_6_io_ins_0 = ces_29_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_6_io_ins_1 = ces_30_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_6_io_ins_2 = ces_31_6_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_6_io_ins_3 = ces_30_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_7_clock = clock;
  assign ces_30_7_io_ins_0 = ces_29_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_7_io_ins_1 = ces_30_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_7_io_ins_2 = ces_31_7_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_7_io_ins_3 = ces_30_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_8_clock = clock;
  assign ces_30_8_io_ins_0 = ces_29_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_8_io_ins_1 = ces_30_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_8_io_ins_2 = ces_31_8_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_8_io_ins_3 = ces_30_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_9_clock = clock;
  assign ces_30_9_io_ins_0 = ces_29_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_9_io_ins_1 = ces_30_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_9_io_ins_2 = ces_31_9_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_9_io_ins_3 = ces_30_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_10_clock = clock;
  assign ces_30_10_io_ins_0 = ces_29_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_10_io_ins_1 = ces_30_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_10_io_ins_2 = ces_31_10_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_10_io_ins_3 = ces_30_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_11_clock = clock;
  assign ces_30_11_io_ins_0 = ces_29_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_11_io_ins_1 = ces_30_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_11_io_ins_2 = ces_31_11_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_11_io_ins_3 = ces_30_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_12_clock = clock;
  assign ces_30_12_io_ins_0 = ces_29_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_12_io_ins_1 = ces_30_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_12_io_ins_2 = ces_31_12_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_12_io_ins_3 = ces_30_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_13_clock = clock;
  assign ces_30_13_io_ins_0 = ces_29_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_13_io_ins_1 = ces_30_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_13_io_ins_2 = ces_31_13_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_13_io_ins_3 = ces_30_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_14_clock = clock;
  assign ces_30_14_io_ins_0 = ces_29_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_14_io_ins_1 = ces_30_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_14_io_ins_2 = ces_31_14_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_14_io_ins_3 = ces_30_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_15_clock = clock;
  assign ces_30_15_io_ins_0 = ces_29_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_15_io_ins_1 = ces_30_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_15_io_ins_2 = ces_31_15_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_15_io_ins_3 = ces_30_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_16_clock = clock;
  assign ces_30_16_io_ins_0 = ces_29_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_16_io_ins_1 = ces_30_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_16_io_ins_2 = ces_31_16_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_16_io_ins_3 = ces_30_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_17_clock = clock;
  assign ces_30_17_io_ins_0 = ces_29_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_17_io_ins_1 = ces_30_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_17_io_ins_2 = ces_31_17_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_17_io_ins_3 = ces_30_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_18_clock = clock;
  assign ces_30_18_io_ins_0 = ces_29_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_18_io_ins_1 = ces_30_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_18_io_ins_2 = ces_31_18_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_18_io_ins_3 = ces_30_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_19_clock = clock;
  assign ces_30_19_io_ins_0 = ces_29_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_19_io_ins_1 = ces_30_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_19_io_ins_2 = ces_31_19_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_19_io_ins_3 = ces_30_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_20_clock = clock;
  assign ces_30_20_io_ins_0 = ces_29_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_20_io_ins_1 = ces_30_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_20_io_ins_2 = ces_31_20_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_20_io_ins_3 = ces_30_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_21_clock = clock;
  assign ces_30_21_io_ins_0 = ces_29_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_21_io_ins_1 = ces_30_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_21_io_ins_2 = ces_31_21_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_21_io_ins_3 = ces_30_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_22_clock = clock;
  assign ces_30_22_io_ins_0 = ces_29_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_22_io_ins_1 = ces_30_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_22_io_ins_2 = ces_31_22_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_22_io_ins_3 = ces_30_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_23_clock = clock;
  assign ces_30_23_io_ins_0 = ces_29_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_23_io_ins_1 = ces_30_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_23_io_ins_2 = ces_31_23_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_23_io_ins_3 = ces_30_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_24_clock = clock;
  assign ces_30_24_io_ins_0 = ces_29_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_24_io_ins_1 = ces_30_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_24_io_ins_2 = ces_31_24_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_24_io_ins_3 = ces_30_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_25_clock = clock;
  assign ces_30_25_io_ins_0 = ces_29_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_25_io_ins_1 = ces_30_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_25_io_ins_2 = ces_31_25_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_25_io_ins_3 = ces_30_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_26_clock = clock;
  assign ces_30_26_io_ins_0 = ces_29_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_26_io_ins_1 = ces_30_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_26_io_ins_2 = ces_31_26_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_26_io_ins_3 = ces_30_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_27_clock = clock;
  assign ces_30_27_io_ins_0 = ces_29_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_27_io_ins_1 = ces_30_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_27_io_ins_2 = ces_31_27_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_27_io_ins_3 = ces_30_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_28_clock = clock;
  assign ces_30_28_io_ins_0 = ces_29_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_28_io_ins_1 = ces_30_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_28_io_ins_2 = ces_31_28_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_28_io_ins_3 = ces_30_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_29_clock = clock;
  assign ces_30_29_io_ins_0 = ces_29_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_29_io_ins_1 = ces_30_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_29_io_ins_2 = ces_31_29_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_29_io_ins_3 = ces_30_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_30_clock = clock;
  assign ces_30_30_io_ins_0 = ces_29_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_30_io_ins_1 = ces_30_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_30_30_io_ins_2 = ces_31_30_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_30_io_ins_3 = ces_30_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_30_31_clock = clock;
  assign ces_30_31_io_ins_0 = ces_29_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_31_io_ins_1 = io_insVertical_0_30; // @[MockArray.scala 45:87]
  assign ces_30_31_io_ins_2 = ces_31_31_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_31_io_ins_3 = ces_30_30_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_0_clock = clock;
  assign ces_31_0_io_ins_0 = ces_30_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_0_io_ins_1 = ces_31_1_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_0_io_ins_2 = io_insHorizontal_1_0; // @[MockArray.scala 46:87]
  assign ces_31_0_io_ins_3 = io_insVertical_1_31; // @[MockArray.scala 47:87]
  assign ces_31_1_clock = clock;
  assign ces_31_1_io_ins_0 = ces_30_1_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_1_io_ins_1 = ces_31_2_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_1_io_ins_2 = io_insHorizontal_1_1; // @[MockArray.scala 46:87]
  assign ces_31_1_io_ins_3 = ces_31_0_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_2_clock = clock;
  assign ces_31_2_io_ins_0 = ces_30_2_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_2_io_ins_1 = ces_31_3_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_2_io_ins_2 = io_insHorizontal_1_2; // @[MockArray.scala 46:87]
  assign ces_31_2_io_ins_3 = ces_31_1_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_3_clock = clock;
  assign ces_31_3_io_ins_0 = ces_30_3_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_3_io_ins_1 = ces_31_4_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_3_io_ins_2 = io_insHorizontal_1_3; // @[MockArray.scala 46:87]
  assign ces_31_3_io_ins_3 = ces_31_2_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_4_clock = clock;
  assign ces_31_4_io_ins_0 = ces_30_4_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_4_io_ins_1 = ces_31_5_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_4_io_ins_2 = io_insHorizontal_1_4; // @[MockArray.scala 46:87]
  assign ces_31_4_io_ins_3 = ces_31_3_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_5_clock = clock;
  assign ces_31_5_io_ins_0 = ces_30_5_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_5_io_ins_1 = ces_31_6_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_5_io_ins_2 = io_insHorizontal_1_5; // @[MockArray.scala 46:87]
  assign ces_31_5_io_ins_3 = ces_31_4_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_6_clock = clock;
  assign ces_31_6_io_ins_0 = ces_30_6_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_6_io_ins_1 = ces_31_7_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_6_io_ins_2 = io_insHorizontal_1_6; // @[MockArray.scala 46:87]
  assign ces_31_6_io_ins_3 = ces_31_5_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_7_clock = clock;
  assign ces_31_7_io_ins_0 = ces_30_7_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_7_io_ins_1 = ces_31_8_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_7_io_ins_2 = io_insHorizontal_1_7; // @[MockArray.scala 46:87]
  assign ces_31_7_io_ins_3 = ces_31_6_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_8_clock = clock;
  assign ces_31_8_io_ins_0 = ces_30_8_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_8_io_ins_1 = ces_31_9_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_8_io_ins_2 = io_insHorizontal_1_8; // @[MockArray.scala 46:87]
  assign ces_31_8_io_ins_3 = ces_31_7_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_9_clock = clock;
  assign ces_31_9_io_ins_0 = ces_30_9_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_9_io_ins_1 = ces_31_10_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_9_io_ins_2 = io_insHorizontal_1_9; // @[MockArray.scala 46:87]
  assign ces_31_9_io_ins_3 = ces_31_8_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_10_clock = clock;
  assign ces_31_10_io_ins_0 = ces_30_10_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_10_io_ins_1 = ces_31_11_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_10_io_ins_2 = io_insHorizontal_1_10; // @[MockArray.scala 46:87]
  assign ces_31_10_io_ins_3 = ces_31_9_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_11_clock = clock;
  assign ces_31_11_io_ins_0 = ces_30_11_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_11_io_ins_1 = ces_31_12_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_11_io_ins_2 = io_insHorizontal_1_11; // @[MockArray.scala 46:87]
  assign ces_31_11_io_ins_3 = ces_31_10_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_12_clock = clock;
  assign ces_31_12_io_ins_0 = ces_30_12_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_12_io_ins_1 = ces_31_13_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_12_io_ins_2 = io_insHorizontal_1_12; // @[MockArray.scala 46:87]
  assign ces_31_12_io_ins_3 = ces_31_11_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_13_clock = clock;
  assign ces_31_13_io_ins_0 = ces_30_13_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_13_io_ins_1 = ces_31_14_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_13_io_ins_2 = io_insHorizontal_1_13; // @[MockArray.scala 46:87]
  assign ces_31_13_io_ins_3 = ces_31_12_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_14_clock = clock;
  assign ces_31_14_io_ins_0 = ces_30_14_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_14_io_ins_1 = ces_31_15_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_14_io_ins_2 = io_insHorizontal_1_14; // @[MockArray.scala 46:87]
  assign ces_31_14_io_ins_3 = ces_31_13_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_15_clock = clock;
  assign ces_31_15_io_ins_0 = ces_30_15_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_15_io_ins_1 = ces_31_16_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_15_io_ins_2 = io_insHorizontal_1_15; // @[MockArray.scala 46:87]
  assign ces_31_15_io_ins_3 = ces_31_14_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_16_clock = clock;
  assign ces_31_16_io_ins_0 = ces_30_16_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_16_io_ins_1 = ces_31_17_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_16_io_ins_2 = io_insHorizontal_1_16; // @[MockArray.scala 46:87]
  assign ces_31_16_io_ins_3 = ces_31_15_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_17_clock = clock;
  assign ces_31_17_io_ins_0 = ces_30_17_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_17_io_ins_1 = ces_31_18_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_17_io_ins_2 = io_insHorizontal_1_17; // @[MockArray.scala 46:87]
  assign ces_31_17_io_ins_3 = ces_31_16_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_18_clock = clock;
  assign ces_31_18_io_ins_0 = ces_30_18_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_18_io_ins_1 = ces_31_19_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_18_io_ins_2 = io_insHorizontal_1_18; // @[MockArray.scala 46:87]
  assign ces_31_18_io_ins_3 = ces_31_17_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_19_clock = clock;
  assign ces_31_19_io_ins_0 = ces_30_19_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_19_io_ins_1 = ces_31_20_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_19_io_ins_2 = io_insHorizontal_1_19; // @[MockArray.scala 46:87]
  assign ces_31_19_io_ins_3 = ces_31_18_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_20_clock = clock;
  assign ces_31_20_io_ins_0 = ces_30_20_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_20_io_ins_1 = ces_31_21_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_20_io_ins_2 = io_insHorizontal_1_20; // @[MockArray.scala 46:87]
  assign ces_31_20_io_ins_3 = ces_31_19_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_21_clock = clock;
  assign ces_31_21_io_ins_0 = ces_30_21_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_21_io_ins_1 = ces_31_22_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_21_io_ins_2 = io_insHorizontal_1_21; // @[MockArray.scala 46:87]
  assign ces_31_21_io_ins_3 = ces_31_20_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_22_clock = clock;
  assign ces_31_22_io_ins_0 = ces_30_22_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_22_io_ins_1 = ces_31_23_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_22_io_ins_2 = io_insHorizontal_1_22; // @[MockArray.scala 46:87]
  assign ces_31_22_io_ins_3 = ces_31_21_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_23_clock = clock;
  assign ces_31_23_io_ins_0 = ces_30_23_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_23_io_ins_1 = ces_31_24_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_23_io_ins_2 = io_insHorizontal_1_23; // @[MockArray.scala 46:87]
  assign ces_31_23_io_ins_3 = ces_31_22_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_24_clock = clock;
  assign ces_31_24_io_ins_0 = ces_30_24_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_24_io_ins_1 = ces_31_25_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_24_io_ins_2 = io_insHorizontal_1_24; // @[MockArray.scala 46:87]
  assign ces_31_24_io_ins_3 = ces_31_23_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_25_clock = clock;
  assign ces_31_25_io_ins_0 = ces_30_25_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_25_io_ins_1 = ces_31_26_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_25_io_ins_2 = io_insHorizontal_1_25; // @[MockArray.scala 46:87]
  assign ces_31_25_io_ins_3 = ces_31_24_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_26_clock = clock;
  assign ces_31_26_io_ins_0 = ces_30_26_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_26_io_ins_1 = ces_31_27_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_26_io_ins_2 = io_insHorizontal_1_26; // @[MockArray.scala 46:87]
  assign ces_31_26_io_ins_3 = ces_31_25_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_27_clock = clock;
  assign ces_31_27_io_ins_0 = ces_30_27_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_27_io_ins_1 = ces_31_28_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_27_io_ins_2 = io_insHorizontal_1_27; // @[MockArray.scala 46:87]
  assign ces_31_27_io_ins_3 = ces_31_26_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_28_clock = clock;
  assign ces_31_28_io_ins_0 = ces_30_28_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_28_io_ins_1 = ces_31_29_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_28_io_ins_2 = io_insHorizontal_1_28; // @[MockArray.scala 46:87]
  assign ces_31_28_io_ins_3 = ces_31_27_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_29_clock = clock;
  assign ces_31_29_io_ins_0 = ces_30_29_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_29_io_ins_1 = ces_31_30_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_29_io_ins_2 = io_insHorizontal_1_29; // @[MockArray.scala 46:87]
  assign ces_31_29_io_ins_3 = ces_31_28_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_30_clock = clock;
  assign ces_31_30_io_ins_0 = ces_30_30_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_30_io_ins_1 = ces_31_31_io_outs_3; // @[MockArray.scala 62:19]
  assign ces_31_30_io_ins_2 = io_insHorizontal_1_30; // @[MockArray.scala 46:87]
  assign ces_31_30_io_ins_3 = ces_31_29_io_outs_1; // @[MockArray.scala 63:19]
  assign ces_31_31_clock = clock;
  assign ces_31_31_io_ins_0 = ces_30_31_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_31_io_ins_1 = io_insVertical_0_31; // @[MockArray.scala 45:87]
  assign ces_31_31_io_ins_2 = io_insHorizontal_1_31; // @[MockArray.scala 46:87]
  assign ces_31_31_io_ins_3 = ces_31_30_io_outs_1; // @[MockArray.scala 63:19]
endmodule
