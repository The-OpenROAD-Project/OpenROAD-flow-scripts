(* blackbox *) module AND2_X1 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AND2_X2 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AND2_X4 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AND3_X1 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AND3_X2 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AND3_X4 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AND4_X1 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AND4_X2 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AND4_X4 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module ANTENNA_X1 (A, VDD, VSS);
  input A;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI211_X1 (A, B, C1, C2, ZN, VDD, VSS);
  input A;
  input B;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI211_X2 (A, B, C1, C2, ZN, VDD, VSS);
  input A;
  input B;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI211_X4 (A, B, C1, C2, ZN, VDD, VSS);
  input A;
  input B;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI21_X1 (A, B1, B2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI21_X2 (A, B1, B2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI21_X4 (A, B1, B2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI221_X1 (A, B1, B2, C1, C2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI221_X2 (A, B1, B2, C1, C2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI221_X4 (A, B1, B2, C1, C2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI222_X1 (A1, A2, B1, B2, C1, C2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI222_X2 (A1, A2, B1, B2, C1, C2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI222_X4 (A1, A2, B1, B2, C1, C2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI22_X1 (A1, A2, B1, B2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI22_X2 (A1, A2, B1, B2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module AOI22_X4 (A1, A2, B1, B2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module BUF_X1 (A, Z, VDD, VSS);
  input A;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module BUF_X16 (A, Z, VDD, VSS);
  input A;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module BUF_X2 (A, Z, VDD, VSS);
  input A;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module BUF_X32 (A, Z, VDD, VSS);
  input A;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module BUF_X4 (A, Z, VDD, VSS);
  input A;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module BUF_X8 (A, Z, VDD, VSS);
  input A;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKBUF_X1 (A, Z, VDD, VSS);
  input A;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKBUF_X2 (A, Z, VDD, VSS);
  input A;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKBUF_X3 (A, Z, VDD, VSS);
  input A;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKGATETST_X1 (CK, E, SE, GCK, VDD, VSS);
  input CK;
  input E;
  input SE;
  output GCK;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKGATETST_X2 (CK, E, SE, GCK, VDD, VSS);
  input CK;
  input E;
  input SE;
  output GCK;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKGATETST_X4 (CK, E, SE, GCK, VDD, VSS);
  input CK;
  input E;
  input SE;
  output GCK;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKGATETST_X8 (CK, E, SE, GCK, VDD, VSS);
  input CK;
  input E;
  input SE;
  output GCK;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKGATE_X1 (CK, E, GCK, VDD, VSS);
  input CK;
  input E;
  output GCK;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKGATE_X2 (CK, E, GCK, VDD, VSS);
  input CK;
  input E;
  output GCK;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKGATE_X4 (CK, E, GCK, VDD, VSS);
  input CK;
  input E;
  output GCK;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module CLKGATE_X8 (CK, E, GCK, VDD, VSS);
  input CK;
  input E;
  output GCK;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DFFRS_X1 (D, RN, SN, CK, Q, QN, VDD, VSS);
  input D;
  input RN;
  input SN;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DFFRS_X2 (D, RN, SN, CK, Q, QN, VDD, VSS);
  input D;
  input RN;
  input SN;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DFFR_X1 (D, RN, CK, Q, QN, VDD, VSS);
  input D;
  input RN;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DFFR_X2 (D, RN, CK, Q, QN, VDD, VSS);
  input D;
  input RN;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DFFS_X1 (D, SN, CK, Q, QN, VDD, VSS);
  input D;
  input SN;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DFFS_X2 (D, SN, CK, Q, QN, VDD, VSS);
  input D;
  input SN;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DFF_X1 (D, CK, Q, QN, VDD, VSS);
  input D;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DFF_X2 (D, CK, Q, QN, VDD, VSS);
  input D;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DLH_X1 (D, G, Q, VDD, VSS);
  input D;
  input G;
  output Q;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DLH_X2 (D, G, Q, VDD, VSS);
  input D;
  input G;
  output Q;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DLL_X1 (D, GN, Q, VDD, VSS);
  input D;
  input GN;
  output Q;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module DLL_X2 (D, GN, Q, VDD, VSS);
  input D;
  input GN;
  output Q;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module FA_X1 (A, B, CI, CO, S, VDD, VSS);
  input A;
  input B;
  input CI;
  output CO;
  output S;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module FILLCELL_X1 (VDD, VSS);
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module FILLCELL_X2 (VDD, VSS);
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module FILLCELL_X4 (VDD, VSS);
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module FILLCELL_X8 (VDD, VSS);
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module FILLCELL_X16 (VDD, VSS);
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module FILLCELL_X32 (VDD, VSS);
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module HA_X1 (A, B, CO, S, VDD, VSS);
  input A;
  input B;
  output CO;
  output S;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module INV_X1 (A, ZN, VDD, VSS);
  input A;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module INV_X16 (A, ZN, VDD, VSS);
  input A;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module INV_X2 (A, ZN, VDD, VSS);
  input A;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module INV_X32 (A, ZN, VDD, VSS);
  input A;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module INV_X4 (A, ZN, VDD, VSS);
  input A;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module INV_X8 (A, ZN, VDD, VSS);
  input A;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module LOGIC0_X1 (Z, VDD, VSS);
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module LOGIC1_X1 (Z, VDD, VSS);
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module MUX2_X1 (A, B, S, Z, VDD, VSS);
  input A;
  input B;
  input S;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module MUX2_X2 (A, B, S, Z, VDD, VSS);
  input A;
  input B;
  input S;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NAND2_X1 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NAND2_X2 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NAND2_X4 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NAND3_X1 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NAND3_X2 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NAND3_X4 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NAND4_X1 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NAND4_X2 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NAND4_X4 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NOR2_X1 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NOR2_X2 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NOR2_X4 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NOR3_X1 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NOR3_X2 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NOR3_X4 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NOR4_X1 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NOR4_X2 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module NOR4_X4 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI211_X1 (A, B, C1, C2, ZN, VDD, VSS);
  input A;
  input B;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI211_X2 (A, B, C1, C2, ZN, VDD, VSS);
  input A;
  input B;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI211_X4 (A, B, C1, C2, ZN, VDD, VSS);
  input A;
  input B;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI21_X1 (A, B1, B2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI21_X2 (A, B1, B2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI21_X4 (A, B1, B2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI221_X1 (A, B1, B2, C1, C2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI221_X2 (A, B1, B2, C1, C2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI221_X4 (A, B1, B2, C1, C2, ZN, VDD, VSS);
  input A;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI222_X1 (A1, A2, B1, B2, C1, C2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI222_X2 (A1, A2, B1, B2, C1, C2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI222_X4 (A1, A2, B1, B2, C1, C2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  input C1;
  input C2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI22_X1 (A1, A2, B1, B2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI22_X2 (A1, A2, B1, B2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI22_X4 (A1, A2, B1, B2, ZN, VDD, VSS);
  input A1;
  input A2;
  input B1;
  input B2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OAI33_X1 (A1, A2, A3, B1, B2, B3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input B1;
  input B2;
  input B3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OR2_X1 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OR2_X2 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OR2_X4 (A1, A2, ZN, VDD, VSS);
  input A1;
  input A2;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OR3_X1 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OR3_X2 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OR3_X4 (A1, A2, A3, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OR4_X1 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OR4_X2 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module OR4_X4 (A1, A2, A3, A4, ZN, VDD, VSS);
  input A1;
  input A2;
  input A3;
  input A4;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module SDFFRS_X1 (D, RN, SE, SI, SN, CK, Q, QN, VDD, VSS);
  input D;
  input RN;
  input SE;
  input SI;
  input SN;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module SDFFRS_X2 (D, RN, SE, SI, SN, CK, Q, QN, VDD, VSS);
  input D;
  input RN;
  input SE;
  input SI;
  input SN;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module SDFFR_X1 (D, RN, SE, SI, CK, Q, QN, VDD, VSS);
  input D;
  input RN;
  input SE;
  input SI;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module SDFFR_X2 (D, RN, SE, SI, CK, Q, QN, VDD, VSS);
  input D;
  input RN;
  input SE;
  input SI;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module SDFFS_X1 (D, SE, SI, SN, CK, Q, QN, VDD, VSS);
  input D;
  input SE;
  input SI;
  input SN;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module SDFFS_X2 (D, SE, SI, SN, CK, Q, QN, VDD, VSS);
  input D;
  input SE;
  input SI;
  input SN;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module SDFF_X1 (D, SE, SI, CK, Q, QN, VDD, VSS);
  input D;
  input SE;
  input SI;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module SDFF_X2 (D, SE, SI, CK, Q, QN, VDD, VSS);
  input D;
  input SE;
  input SI;
  input CK;
  output Q;
  output QN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module TBUF_X1 (A, EN, Z, VDD, VSS);
  input A;
  input EN;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module TBUF_X16 (A, EN, Z, VDD, VSS);
  input A;
  input EN;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module TBUF_X2 (A, EN, Z, VDD, VSS);
  input A;
  input EN;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module TBUF_X4 (A, EN, Z, VDD, VSS);
  input A;
  input EN;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module TBUF_X8 (A, EN, Z, VDD, VSS);
  input A;
  input EN;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module TINV_X1 (EN, I, ZN, VDD, VSS);
  input EN;
  input I;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module TLAT_X1 (D, G, OE, Q, VDD, VSS);
  input D;
  input G;
  input OE;
  output Q;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module XNOR2_X1 (A, B, ZN, VDD, VSS);
  input A;
  input B;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module XNOR2_X2 (A, B, ZN, VDD, VSS);
  input A;
  input B;
  output ZN;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module XOR2_X1 (A, B, Z, VDD, VSS);
  input A;
  input B;
  output Z;
  inout VDD;
  inout VSS;
endmodule
(* blackbox *) module XOR2_X2 (A, B, Z, VDD, VSS);
  input A;
  input B;
  output Z;
  inout VDD;
  inout VSS;
endmodule
