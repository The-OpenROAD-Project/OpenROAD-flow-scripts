VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_512x64
  FOREIGN fakeram45_512x64 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 152.570 BY 113.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.785 0.070 1.855 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.205 0.070 2.275 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.625 0.070 2.695 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.465 0.070 3.535 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.305 0.070 4.375 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.145 0.070 5.215 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.985 0.070 6.055 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.825 0.070 6.895 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.665 0.070 7.735 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.505 0.070 8.575 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.925 0.070 8.995 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.345 0.070 9.415 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.185 0.070 10.255 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.025 0.070 11.095 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.865 0.070 11.935 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.285 0.070 12.355 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.705 0.070 12.775 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.545 0.070 13.615 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.385 0.070 14.455 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.805 0.070 14.875 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.225 0.070 15.295 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.645 0.070 15.715 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.065 0.070 16.135 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.485 0.070 16.555 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.905 0.070 16.975 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.745 0.070 17.815 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.585 0.070 18.655 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.425 0.070 19.495 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.845 0.070 19.915 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.265 0.070 20.335 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.685 0.070 20.755 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.105 0.070 21.175 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.525 0.070 21.595 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.945 0.070 22.015 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.785 0.070 22.855 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.625 0.070 23.695 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.045 0.070 24.115 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.465 0.070 24.535 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.305 0.070 25.375 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.725 0.070 25.795 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.145 0.070 26.215 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.985 0.070 27.055 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.405 0.070 27.475 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.825 0.070 27.895 ;
    END
  END w_mask_in[63]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.985 0.070 34.055 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.825 0.070 34.895 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.245 0.070 35.315 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.665 0.070 35.735 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.085 0.070 36.155 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.925 0.070 36.995 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.765 0.070 37.835 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.605 0.070 38.675 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.445 0.070 39.515 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.125 0.070 41.195 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.965 0.070 42.035 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.805 0.070 42.875 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.645 0.070 43.715 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.485 0.070 44.555 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.325 0.070 45.395 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.005 0.070 47.075 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.845 0.070 47.915 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.685 0.070 48.755 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.365 0.070 50.435 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.205 0.070 51.275 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.045 0.070 52.115 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.885 0.070 52.955 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.725 0.070 53.795 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.565 0.070 54.635 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.245 0.070 56.315 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.085 0.070 57.155 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.925 0.070 57.995 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.765 0.070 58.835 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.605 0.070 59.675 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.445 0.070 60.515 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 66.605 0.070 66.675 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.025 0.070 67.095 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.445 0.070 67.515 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.865 0.070 67.935 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.285 0.070 68.355 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.705 0.070 68.775 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.125 0.070 69.195 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.545 0.070 69.615 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 69.965 0.070 70.035 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.385 0.070 70.455 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.805 0.070 70.875 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.225 0.070 71.295 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.645 0.070 71.715 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.065 0.070 72.135 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.485 0.070 72.555 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.905 0.070 72.975 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.325 0.070 73.395 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.745 0.070 73.815 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.585 0.070 74.655 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.005 0.070 75.075 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.425 0.070 75.495 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.265 0.070 76.335 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.685 0.070 76.755 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.105 0.070 77.175 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.525 0.070 77.595 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.945 0.070 78.015 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.365 0.070 78.435 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.785 0.070 78.855 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.205 0.070 79.275 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.625 0.070 79.695 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.045 0.070 80.115 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.465 0.070 80.535 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.885 0.070 80.955 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.305 0.070 81.375 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.725 0.070 81.795 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.145 0.070 82.215 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.985 0.070 83.055 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.405 0.070 83.475 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.825 0.070 83.895 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.245 0.070 84.315 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.665 0.070 84.735 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.085 0.070 85.155 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.505 0.070 85.575 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.925 0.070 85.995 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.345 0.070 86.415 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.765 0.070 86.835 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.185 0.070 87.255 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.605 0.070 87.675 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.025 0.070 88.095 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.445 0.070 88.515 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.865 0.070 88.935 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.285 0.070 89.355 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.705 0.070 89.775 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.125 0.070 90.195 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.545 0.070 90.615 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.965 0.070 91.035 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.385 0.070 91.455 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.805 0.070 91.875 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.225 0.070 92.295 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.645 0.070 92.715 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.065 0.070 93.135 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.225 0.070 99.295 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.645 0.070 99.715 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.065 0.070 100.135 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.485 0.070 100.555 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 100.905 0.070 100.975 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.325 0.070 101.395 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.745 0.070 101.815 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.165 0.070 102.235 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.585 0.070 102.655 ;
    END
  END addr_in[8]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.745 0.070 108.815 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.165 0.070 109.235 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 109.585 0.070 109.655 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 112.000 ;
      RECT 3.500 1.400 3.780 112.000 ;
      RECT 5.740 1.400 6.020 112.000 ;
      RECT 7.980 1.400 8.260 112.000 ;
      RECT 10.220 1.400 10.500 112.000 ;
      RECT 12.460 1.400 12.740 112.000 ;
      RECT 14.700 1.400 14.980 112.000 ;
      RECT 16.940 1.400 17.220 112.000 ;
      RECT 19.180 1.400 19.460 112.000 ;
      RECT 21.420 1.400 21.700 112.000 ;
      RECT 23.660 1.400 23.940 112.000 ;
      RECT 25.900 1.400 26.180 112.000 ;
      RECT 28.140 1.400 28.420 112.000 ;
      RECT 30.380 1.400 30.660 112.000 ;
      RECT 32.620 1.400 32.900 112.000 ;
      RECT 34.860 1.400 35.140 112.000 ;
      RECT 37.100 1.400 37.380 112.000 ;
      RECT 39.340 1.400 39.620 112.000 ;
      RECT 41.580 1.400 41.860 112.000 ;
      RECT 43.820 1.400 44.100 112.000 ;
      RECT 46.060 1.400 46.340 112.000 ;
      RECT 48.300 1.400 48.580 112.000 ;
      RECT 50.540 1.400 50.820 112.000 ;
      RECT 52.780 1.400 53.060 112.000 ;
      RECT 55.020 1.400 55.300 112.000 ;
      RECT 57.260 1.400 57.540 112.000 ;
      RECT 59.500 1.400 59.780 112.000 ;
      RECT 61.740 1.400 62.020 112.000 ;
      RECT 63.980 1.400 64.260 112.000 ;
      RECT 66.220 1.400 66.500 112.000 ;
      RECT 68.460 1.400 68.740 112.000 ;
      RECT 70.700 1.400 70.980 112.000 ;
      RECT 72.940 1.400 73.220 112.000 ;
      RECT 75.180 1.400 75.460 112.000 ;
      RECT 77.420 1.400 77.700 112.000 ;
      RECT 79.660 1.400 79.940 112.000 ;
      RECT 81.900 1.400 82.180 112.000 ;
      RECT 84.140 1.400 84.420 112.000 ;
      RECT 86.380 1.400 86.660 112.000 ;
      RECT 88.620 1.400 88.900 112.000 ;
      RECT 90.860 1.400 91.140 112.000 ;
      RECT 93.100 1.400 93.380 112.000 ;
      RECT 95.340 1.400 95.620 112.000 ;
      RECT 97.580 1.400 97.860 112.000 ;
      RECT 99.820 1.400 100.100 112.000 ;
      RECT 102.060 1.400 102.340 112.000 ;
      RECT 104.300 1.400 104.580 112.000 ;
      RECT 106.540 1.400 106.820 112.000 ;
      RECT 108.780 1.400 109.060 112.000 ;
      RECT 111.020 1.400 111.300 112.000 ;
      RECT 113.260 1.400 113.540 112.000 ;
      RECT 115.500 1.400 115.780 112.000 ;
      RECT 117.740 1.400 118.020 112.000 ;
      RECT 119.980 1.400 120.260 112.000 ;
      RECT 122.220 1.400 122.500 112.000 ;
      RECT 124.460 1.400 124.740 112.000 ;
      RECT 126.700 1.400 126.980 112.000 ;
      RECT 128.940 1.400 129.220 112.000 ;
      RECT 131.180 1.400 131.460 112.000 ;
      RECT 133.420 1.400 133.700 112.000 ;
      RECT 135.660 1.400 135.940 112.000 ;
      RECT 137.900 1.400 138.180 112.000 ;
      RECT 140.140 1.400 140.420 112.000 ;
      RECT 142.380 1.400 142.660 112.000 ;
      RECT 144.620 1.400 144.900 112.000 ;
      RECT 146.860 1.400 147.140 112.000 ;
      RECT 149.100 1.400 149.380 112.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 112.000 ;
      RECT 4.620 1.400 4.900 112.000 ;
      RECT 6.860 1.400 7.140 112.000 ;
      RECT 9.100 1.400 9.380 112.000 ;
      RECT 11.340 1.400 11.620 112.000 ;
      RECT 13.580 1.400 13.860 112.000 ;
      RECT 15.820 1.400 16.100 112.000 ;
      RECT 18.060 1.400 18.340 112.000 ;
      RECT 20.300 1.400 20.580 112.000 ;
      RECT 22.540 1.400 22.820 112.000 ;
      RECT 24.780 1.400 25.060 112.000 ;
      RECT 27.020 1.400 27.300 112.000 ;
      RECT 29.260 1.400 29.540 112.000 ;
      RECT 31.500 1.400 31.780 112.000 ;
      RECT 33.740 1.400 34.020 112.000 ;
      RECT 35.980 1.400 36.260 112.000 ;
      RECT 38.220 1.400 38.500 112.000 ;
      RECT 40.460 1.400 40.740 112.000 ;
      RECT 42.700 1.400 42.980 112.000 ;
      RECT 44.940 1.400 45.220 112.000 ;
      RECT 47.180 1.400 47.460 112.000 ;
      RECT 49.420 1.400 49.700 112.000 ;
      RECT 51.660 1.400 51.940 112.000 ;
      RECT 53.900 1.400 54.180 112.000 ;
      RECT 56.140 1.400 56.420 112.000 ;
      RECT 58.380 1.400 58.660 112.000 ;
      RECT 60.620 1.400 60.900 112.000 ;
      RECT 62.860 1.400 63.140 112.000 ;
      RECT 65.100 1.400 65.380 112.000 ;
      RECT 67.340 1.400 67.620 112.000 ;
      RECT 69.580 1.400 69.860 112.000 ;
      RECT 71.820 1.400 72.100 112.000 ;
      RECT 74.060 1.400 74.340 112.000 ;
      RECT 76.300 1.400 76.580 112.000 ;
      RECT 78.540 1.400 78.820 112.000 ;
      RECT 80.780 1.400 81.060 112.000 ;
      RECT 83.020 1.400 83.300 112.000 ;
      RECT 85.260 1.400 85.540 112.000 ;
      RECT 87.500 1.400 87.780 112.000 ;
      RECT 89.740 1.400 90.020 112.000 ;
      RECT 91.980 1.400 92.260 112.000 ;
      RECT 94.220 1.400 94.500 112.000 ;
      RECT 96.460 1.400 96.740 112.000 ;
      RECT 98.700 1.400 98.980 112.000 ;
      RECT 100.940 1.400 101.220 112.000 ;
      RECT 103.180 1.400 103.460 112.000 ;
      RECT 105.420 1.400 105.700 112.000 ;
      RECT 107.660 1.400 107.940 112.000 ;
      RECT 109.900 1.400 110.180 112.000 ;
      RECT 112.140 1.400 112.420 112.000 ;
      RECT 114.380 1.400 114.660 112.000 ;
      RECT 116.620 1.400 116.900 112.000 ;
      RECT 118.860 1.400 119.140 112.000 ;
      RECT 121.100 1.400 121.380 112.000 ;
      RECT 123.340 1.400 123.620 112.000 ;
      RECT 125.580 1.400 125.860 112.000 ;
      RECT 127.820 1.400 128.100 112.000 ;
      RECT 130.060 1.400 130.340 112.000 ;
      RECT 132.300 1.400 132.580 112.000 ;
      RECT 134.540 1.400 134.820 112.000 ;
      RECT 136.780 1.400 137.060 112.000 ;
      RECT 139.020 1.400 139.300 112.000 ;
      RECT 141.260 1.400 141.540 112.000 ;
      RECT 143.500 1.400 143.780 112.000 ;
      RECT 145.740 1.400 146.020 112.000 ;
      RECT 147.980 1.400 148.260 112.000 ;
      RECT 150.220 1.400 150.500 112.000 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 152.570 113.400 ;
    LAYER metal2 ;
    RECT 0 0 152.570 113.400 ;
    LAYER metal3 ;
    RECT 0.070 0 152.570 113.400 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.785 ;
    RECT 0 1.855 0.070 2.205 ;
    RECT 0 2.275 0.070 2.625 ;
    RECT 0 2.695 0.070 3.045 ;
    RECT 0 3.115 0.070 3.465 ;
    RECT 0 3.535 0.070 3.885 ;
    RECT 0 3.955 0.070 4.305 ;
    RECT 0 4.375 0.070 4.725 ;
    RECT 0 4.795 0.070 5.145 ;
    RECT 0 5.215 0.070 5.565 ;
    RECT 0 5.635 0.070 5.985 ;
    RECT 0 6.055 0.070 6.405 ;
    RECT 0 6.475 0.070 6.825 ;
    RECT 0 6.895 0.070 7.245 ;
    RECT 0 7.315 0.070 7.665 ;
    RECT 0 7.735 0.070 8.085 ;
    RECT 0 8.155 0.070 8.505 ;
    RECT 0 8.575 0.070 8.925 ;
    RECT 0 8.995 0.070 9.345 ;
    RECT 0 9.415 0.070 9.765 ;
    RECT 0 9.835 0.070 10.185 ;
    RECT 0 10.255 0.070 10.605 ;
    RECT 0 10.675 0.070 11.025 ;
    RECT 0 11.095 0.070 11.445 ;
    RECT 0 11.515 0.070 11.865 ;
    RECT 0 11.935 0.070 12.285 ;
    RECT 0 12.355 0.070 12.705 ;
    RECT 0 12.775 0.070 13.125 ;
    RECT 0 13.195 0.070 13.545 ;
    RECT 0 13.615 0.070 13.965 ;
    RECT 0 14.035 0.070 14.385 ;
    RECT 0 14.455 0.070 14.805 ;
    RECT 0 14.875 0.070 15.225 ;
    RECT 0 15.295 0.070 15.645 ;
    RECT 0 15.715 0.070 16.065 ;
    RECT 0 16.135 0.070 16.485 ;
    RECT 0 16.555 0.070 16.905 ;
    RECT 0 16.975 0.070 17.325 ;
    RECT 0 17.395 0.070 17.745 ;
    RECT 0 17.815 0.070 18.165 ;
    RECT 0 18.235 0.070 18.585 ;
    RECT 0 18.655 0.070 19.005 ;
    RECT 0 19.075 0.070 19.425 ;
    RECT 0 19.495 0.070 19.845 ;
    RECT 0 19.915 0.070 20.265 ;
    RECT 0 20.335 0.070 20.685 ;
    RECT 0 20.755 0.070 21.105 ;
    RECT 0 21.175 0.070 21.525 ;
    RECT 0 21.595 0.070 21.945 ;
    RECT 0 22.015 0.070 22.365 ;
    RECT 0 22.435 0.070 22.785 ;
    RECT 0 22.855 0.070 23.205 ;
    RECT 0 23.275 0.070 23.625 ;
    RECT 0 23.695 0.070 24.045 ;
    RECT 0 24.115 0.070 24.465 ;
    RECT 0 24.535 0.070 24.885 ;
    RECT 0 24.955 0.070 25.305 ;
    RECT 0 25.375 0.070 25.725 ;
    RECT 0 25.795 0.070 26.145 ;
    RECT 0 26.215 0.070 26.565 ;
    RECT 0 26.635 0.070 26.985 ;
    RECT 0 27.055 0.070 27.405 ;
    RECT 0 27.475 0.070 27.825 ;
    RECT 0 27.895 0.070 33.985 ;
    RECT 0 34.055 0.070 34.405 ;
    RECT 0 34.475 0.070 34.825 ;
    RECT 0 34.895 0.070 35.245 ;
    RECT 0 35.315 0.070 35.665 ;
    RECT 0 35.735 0.070 36.085 ;
    RECT 0 36.155 0.070 36.505 ;
    RECT 0 36.575 0.070 36.925 ;
    RECT 0 36.995 0.070 37.345 ;
    RECT 0 37.415 0.070 37.765 ;
    RECT 0 37.835 0.070 38.185 ;
    RECT 0 38.255 0.070 38.605 ;
    RECT 0 38.675 0.070 39.025 ;
    RECT 0 39.095 0.070 39.445 ;
    RECT 0 39.515 0.070 39.865 ;
    RECT 0 39.935 0.070 40.285 ;
    RECT 0 40.355 0.070 40.705 ;
    RECT 0 40.775 0.070 41.125 ;
    RECT 0 41.195 0.070 41.545 ;
    RECT 0 41.615 0.070 41.965 ;
    RECT 0 42.035 0.070 42.385 ;
    RECT 0 42.455 0.070 42.805 ;
    RECT 0 42.875 0.070 43.225 ;
    RECT 0 43.295 0.070 43.645 ;
    RECT 0 43.715 0.070 44.065 ;
    RECT 0 44.135 0.070 44.485 ;
    RECT 0 44.555 0.070 44.905 ;
    RECT 0 44.975 0.070 45.325 ;
    RECT 0 45.395 0.070 45.745 ;
    RECT 0 45.815 0.070 46.165 ;
    RECT 0 46.235 0.070 46.585 ;
    RECT 0 46.655 0.070 47.005 ;
    RECT 0 47.075 0.070 47.425 ;
    RECT 0 47.495 0.070 47.845 ;
    RECT 0 47.915 0.070 48.265 ;
    RECT 0 48.335 0.070 48.685 ;
    RECT 0 48.755 0.070 49.105 ;
    RECT 0 49.175 0.070 49.525 ;
    RECT 0 49.595 0.070 49.945 ;
    RECT 0 50.015 0.070 50.365 ;
    RECT 0 50.435 0.070 50.785 ;
    RECT 0 50.855 0.070 51.205 ;
    RECT 0 51.275 0.070 51.625 ;
    RECT 0 51.695 0.070 52.045 ;
    RECT 0 52.115 0.070 52.465 ;
    RECT 0 52.535 0.070 52.885 ;
    RECT 0 52.955 0.070 53.305 ;
    RECT 0 53.375 0.070 53.725 ;
    RECT 0 53.795 0.070 54.145 ;
    RECT 0 54.215 0.070 54.565 ;
    RECT 0 54.635 0.070 54.985 ;
    RECT 0 55.055 0.070 55.405 ;
    RECT 0 55.475 0.070 55.825 ;
    RECT 0 55.895 0.070 56.245 ;
    RECT 0 56.315 0.070 56.665 ;
    RECT 0 56.735 0.070 57.085 ;
    RECT 0 57.155 0.070 57.505 ;
    RECT 0 57.575 0.070 57.925 ;
    RECT 0 57.995 0.070 58.345 ;
    RECT 0 58.415 0.070 58.765 ;
    RECT 0 58.835 0.070 59.185 ;
    RECT 0 59.255 0.070 59.605 ;
    RECT 0 59.675 0.070 60.025 ;
    RECT 0 60.095 0.070 60.445 ;
    RECT 0 60.515 0.070 66.605 ;
    RECT 0 66.675 0.070 67.025 ;
    RECT 0 67.095 0.070 67.445 ;
    RECT 0 67.515 0.070 67.865 ;
    RECT 0 67.935 0.070 68.285 ;
    RECT 0 68.355 0.070 68.705 ;
    RECT 0 68.775 0.070 69.125 ;
    RECT 0 69.195 0.070 69.545 ;
    RECT 0 69.615 0.070 69.965 ;
    RECT 0 70.035 0.070 70.385 ;
    RECT 0 70.455 0.070 70.805 ;
    RECT 0 70.875 0.070 71.225 ;
    RECT 0 71.295 0.070 71.645 ;
    RECT 0 71.715 0.070 72.065 ;
    RECT 0 72.135 0.070 72.485 ;
    RECT 0 72.555 0.070 72.905 ;
    RECT 0 72.975 0.070 73.325 ;
    RECT 0 73.395 0.070 73.745 ;
    RECT 0 73.815 0.070 74.165 ;
    RECT 0 74.235 0.070 74.585 ;
    RECT 0 74.655 0.070 75.005 ;
    RECT 0 75.075 0.070 75.425 ;
    RECT 0 75.495 0.070 75.845 ;
    RECT 0 75.915 0.070 76.265 ;
    RECT 0 76.335 0.070 76.685 ;
    RECT 0 76.755 0.070 77.105 ;
    RECT 0 77.175 0.070 77.525 ;
    RECT 0 77.595 0.070 77.945 ;
    RECT 0 78.015 0.070 78.365 ;
    RECT 0 78.435 0.070 78.785 ;
    RECT 0 78.855 0.070 79.205 ;
    RECT 0 79.275 0.070 79.625 ;
    RECT 0 79.695 0.070 80.045 ;
    RECT 0 80.115 0.070 80.465 ;
    RECT 0 80.535 0.070 80.885 ;
    RECT 0 80.955 0.070 81.305 ;
    RECT 0 81.375 0.070 81.725 ;
    RECT 0 81.795 0.070 82.145 ;
    RECT 0 82.215 0.070 82.565 ;
    RECT 0 82.635 0.070 82.985 ;
    RECT 0 83.055 0.070 83.405 ;
    RECT 0 83.475 0.070 83.825 ;
    RECT 0 83.895 0.070 84.245 ;
    RECT 0 84.315 0.070 84.665 ;
    RECT 0 84.735 0.070 85.085 ;
    RECT 0 85.155 0.070 85.505 ;
    RECT 0 85.575 0.070 85.925 ;
    RECT 0 85.995 0.070 86.345 ;
    RECT 0 86.415 0.070 86.765 ;
    RECT 0 86.835 0.070 87.185 ;
    RECT 0 87.255 0.070 87.605 ;
    RECT 0 87.675 0.070 88.025 ;
    RECT 0 88.095 0.070 88.445 ;
    RECT 0 88.515 0.070 88.865 ;
    RECT 0 88.935 0.070 89.285 ;
    RECT 0 89.355 0.070 89.705 ;
    RECT 0 89.775 0.070 90.125 ;
    RECT 0 90.195 0.070 90.545 ;
    RECT 0 90.615 0.070 90.965 ;
    RECT 0 91.035 0.070 91.385 ;
    RECT 0 91.455 0.070 91.805 ;
    RECT 0 91.875 0.070 92.225 ;
    RECT 0 92.295 0.070 92.645 ;
    RECT 0 92.715 0.070 93.065 ;
    RECT 0 93.135 0.070 99.225 ;
    RECT 0 99.295 0.070 99.645 ;
    RECT 0 99.715 0.070 100.065 ;
    RECT 0 100.135 0.070 100.485 ;
    RECT 0 100.555 0.070 100.905 ;
    RECT 0 100.975 0.070 101.325 ;
    RECT 0 101.395 0.070 101.745 ;
    RECT 0 101.815 0.070 102.165 ;
    RECT 0 102.235 0.070 102.585 ;
    RECT 0 102.655 0.070 108.745 ;
    RECT 0 108.815 0.070 109.165 ;
    RECT 0 109.235 0.070 109.585 ;
    RECT 0 109.655 0.070 113.400 ;
    LAYER metal4 ;
    RECT 0 0 152.570 1.400 ;
    RECT 0 112.000 152.570 113.400 ;
    RECT 0.000 1.400 1.260 112.000 ;
    RECT 1.540 1.400 2.380 112.000 ;
    RECT 2.660 1.400 3.500 112.000 ;
    RECT 3.780 1.400 4.620 112.000 ;
    RECT 4.900 1.400 5.740 112.000 ;
    RECT 6.020 1.400 6.860 112.000 ;
    RECT 7.140 1.400 7.980 112.000 ;
    RECT 8.260 1.400 9.100 112.000 ;
    RECT 9.380 1.400 10.220 112.000 ;
    RECT 10.500 1.400 11.340 112.000 ;
    RECT 11.620 1.400 12.460 112.000 ;
    RECT 12.740 1.400 13.580 112.000 ;
    RECT 13.860 1.400 14.700 112.000 ;
    RECT 14.980 1.400 15.820 112.000 ;
    RECT 16.100 1.400 16.940 112.000 ;
    RECT 17.220 1.400 18.060 112.000 ;
    RECT 18.340 1.400 19.180 112.000 ;
    RECT 19.460 1.400 20.300 112.000 ;
    RECT 20.580 1.400 21.420 112.000 ;
    RECT 21.700 1.400 22.540 112.000 ;
    RECT 22.820 1.400 23.660 112.000 ;
    RECT 23.940 1.400 24.780 112.000 ;
    RECT 25.060 1.400 25.900 112.000 ;
    RECT 26.180 1.400 27.020 112.000 ;
    RECT 27.300 1.400 28.140 112.000 ;
    RECT 28.420 1.400 29.260 112.000 ;
    RECT 29.540 1.400 30.380 112.000 ;
    RECT 30.660 1.400 31.500 112.000 ;
    RECT 31.780 1.400 32.620 112.000 ;
    RECT 32.900 1.400 33.740 112.000 ;
    RECT 34.020 1.400 34.860 112.000 ;
    RECT 35.140 1.400 35.980 112.000 ;
    RECT 36.260 1.400 37.100 112.000 ;
    RECT 37.380 1.400 38.220 112.000 ;
    RECT 38.500 1.400 39.340 112.000 ;
    RECT 39.620 1.400 40.460 112.000 ;
    RECT 40.740 1.400 41.580 112.000 ;
    RECT 41.860 1.400 42.700 112.000 ;
    RECT 42.980 1.400 43.820 112.000 ;
    RECT 44.100 1.400 44.940 112.000 ;
    RECT 45.220 1.400 46.060 112.000 ;
    RECT 46.340 1.400 47.180 112.000 ;
    RECT 47.460 1.400 48.300 112.000 ;
    RECT 48.580 1.400 49.420 112.000 ;
    RECT 49.700 1.400 50.540 112.000 ;
    RECT 50.820 1.400 51.660 112.000 ;
    RECT 51.940 1.400 52.780 112.000 ;
    RECT 53.060 1.400 53.900 112.000 ;
    RECT 54.180 1.400 55.020 112.000 ;
    RECT 55.300 1.400 56.140 112.000 ;
    RECT 56.420 1.400 57.260 112.000 ;
    RECT 57.540 1.400 58.380 112.000 ;
    RECT 58.660 1.400 59.500 112.000 ;
    RECT 59.780 1.400 60.620 112.000 ;
    RECT 60.900 1.400 61.740 112.000 ;
    RECT 62.020 1.400 62.860 112.000 ;
    RECT 63.140 1.400 63.980 112.000 ;
    RECT 64.260 1.400 65.100 112.000 ;
    RECT 65.380 1.400 66.220 112.000 ;
    RECT 66.500 1.400 67.340 112.000 ;
    RECT 67.620 1.400 68.460 112.000 ;
    RECT 68.740 1.400 69.580 112.000 ;
    RECT 69.860 1.400 70.700 112.000 ;
    RECT 70.980 1.400 71.820 112.000 ;
    RECT 72.100 1.400 72.940 112.000 ;
    RECT 73.220 1.400 74.060 112.000 ;
    RECT 74.340 1.400 75.180 112.000 ;
    RECT 75.460 1.400 76.300 112.000 ;
    RECT 76.580 1.400 77.420 112.000 ;
    RECT 77.700 1.400 78.540 112.000 ;
    RECT 78.820 1.400 79.660 112.000 ;
    RECT 79.940 1.400 80.780 112.000 ;
    RECT 81.060 1.400 81.900 112.000 ;
    RECT 82.180 1.400 83.020 112.000 ;
    RECT 83.300 1.400 84.140 112.000 ;
    RECT 84.420 1.400 85.260 112.000 ;
    RECT 85.540 1.400 86.380 112.000 ;
    RECT 86.660 1.400 87.500 112.000 ;
    RECT 87.780 1.400 88.620 112.000 ;
    RECT 88.900 1.400 89.740 112.000 ;
    RECT 90.020 1.400 90.860 112.000 ;
    RECT 91.140 1.400 91.980 112.000 ;
    RECT 92.260 1.400 93.100 112.000 ;
    RECT 93.380 1.400 94.220 112.000 ;
    RECT 94.500 1.400 95.340 112.000 ;
    RECT 95.620 1.400 96.460 112.000 ;
    RECT 96.740 1.400 97.580 112.000 ;
    RECT 97.860 1.400 98.700 112.000 ;
    RECT 98.980 1.400 99.820 112.000 ;
    RECT 100.100 1.400 100.940 112.000 ;
    RECT 101.220 1.400 102.060 112.000 ;
    RECT 102.340 1.400 103.180 112.000 ;
    RECT 103.460 1.400 104.300 112.000 ;
    RECT 104.580 1.400 105.420 112.000 ;
    RECT 105.700 1.400 106.540 112.000 ;
    RECT 106.820 1.400 107.660 112.000 ;
    RECT 107.940 1.400 108.780 112.000 ;
    RECT 109.060 1.400 109.900 112.000 ;
    RECT 110.180 1.400 111.020 112.000 ;
    RECT 111.300 1.400 112.140 112.000 ;
    RECT 112.420 1.400 113.260 112.000 ;
    RECT 113.540 1.400 114.380 112.000 ;
    RECT 114.660 1.400 115.500 112.000 ;
    RECT 115.780 1.400 116.620 112.000 ;
    RECT 116.900 1.400 117.740 112.000 ;
    RECT 118.020 1.400 118.860 112.000 ;
    RECT 119.140 1.400 119.980 112.000 ;
    RECT 120.260 1.400 121.100 112.000 ;
    RECT 121.380 1.400 122.220 112.000 ;
    RECT 122.500 1.400 123.340 112.000 ;
    RECT 123.620 1.400 124.460 112.000 ;
    RECT 124.740 1.400 125.580 112.000 ;
    RECT 125.860 1.400 126.700 112.000 ;
    RECT 126.980 1.400 127.820 112.000 ;
    RECT 128.100 1.400 128.940 112.000 ;
    RECT 129.220 1.400 130.060 112.000 ;
    RECT 130.340 1.400 131.180 112.000 ;
    RECT 131.460 1.400 132.300 112.000 ;
    RECT 132.580 1.400 133.420 112.000 ;
    RECT 133.700 1.400 134.540 112.000 ;
    RECT 134.820 1.400 135.660 112.000 ;
    RECT 135.940 1.400 136.780 112.000 ;
    RECT 137.060 1.400 137.900 112.000 ;
    RECT 138.180 1.400 139.020 112.000 ;
    RECT 139.300 1.400 140.140 112.000 ;
    RECT 140.420 1.400 141.260 112.000 ;
    RECT 141.540 1.400 142.380 112.000 ;
    RECT 142.660 1.400 143.500 112.000 ;
    RECT 143.780 1.400 144.620 112.000 ;
    RECT 144.900 1.400 145.740 112.000 ;
    RECT 146.020 1.400 146.860 112.000 ;
    RECT 147.140 1.400 147.980 112.000 ;
    RECT 148.260 1.400 149.100 112.000 ;
    RECT 149.380 1.400 150.220 112.000 ;
    RECT 150.500 1.400 152.570 112.000 ;
    LAYER OVERLAP ;
    RECT 0 0 152.570 113.400 ;
  END
END fakeram45_512x64

END LIBRARY
