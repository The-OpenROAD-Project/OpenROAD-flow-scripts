(* blackbox *) module BUFx10_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx12_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx12f_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx16f_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx24_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx2_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx3_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx4_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx4f_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx5_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx6f_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module BUFx8_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx10_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx11_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx12_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx14_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx16_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx20_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx5p33_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx6p67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx8_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module CKINVDCx9p33_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB1xp67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB2xp67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB3xp67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module HB4xp67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx11_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx13_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx1_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx2_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx3_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx4_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx5_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx6_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVx8_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVxp33_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
(* blackbox *) module INVxp67_ASAP7_75t_L (Y, A);
	output Y;
	input A;
endmodule
