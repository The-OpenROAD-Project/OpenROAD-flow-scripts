/*
 *  Copyright 2023 CEA*
 *  *Commissariat a l'Energie Atomique et aux Energies Alternatives (CEA)
 *
 *  SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
 *
 *  Licensed under the Solderpad Hardware License v 2.1 (the “License”); you
 *  may not use this file except in compliance with the License, or, at your
 *  option, the Apache License version 2.0. You may obtain a copy of the
 *  License at
 *
 *  https://solderpad.org/licenses/SHL-2.1/
 *
 *  Unless required by applicable law or agreed to in writing, any work
 *  distributed under the License is distributed on an “AS IS” BASIS, WITHOUT
 *  WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See the
 *  License for the specific language governing permissions and limitations
 *  under the License.
 */
/*
 *  Authors       : Cesar Fuguet
 *  Creation Date : March, 2020
 *  Description   : Wrapper for Behavioral SRAM macros
 *  History       :
 */
module hpdcache_sram
#(
    parameter int unsigned ADDR_SIZE = 0,
    parameter int unsigned DATA_SIZE = 0,
    parameter int unsigned DEPTH = 2**ADDR_SIZE
)
(
    input  logic                  clk,
    input  logic                  rst_n,
    input  logic                  cs,
    input  logic                  we,
    input  logic [ADDR_SIZE-1:0]  addr,
    input  logic [DATA_SIZE-1:0]  wdata,
    output logic [DATA_SIZE-1:0]  rdata
);

    fakeram7_256x32 ram_i (
        .clk(clk),
        .ce_in(cs),
        .we_in(we),
        .addr_in(addr),
        .wd_in(wdata),
        .rd_out(rdata)
    );
    // hpdcache_sram_1rw #(
    //     .ADDR_SIZE(ADDR_SIZE),
    //     .DATA_SIZE(DATA_SIZE),
    //     .DEPTH(DEPTH)
    // ) ram_i (
    //     .clk,
    //     .rst_n,
    //     .cs,
    //     .we,
    //     .addr,
    //     .wdata,
    //     .rdata
    // );

endmodule : hpdcache_sram
