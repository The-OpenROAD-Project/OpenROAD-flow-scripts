module MuxTest_width_1_inputs_4_outputs_8_pipeline_0( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [1:0] io_selects_0_0, // @[:@6.4]
  input  [1:0] io_selects_0_1, // @[:@6.4]
  input  [1:0] io_selects_1_0, // @[:@6.4]
  input  [1:0] io_selects_1_1, // @[:@6.4]
  input  [1:0] io_selects_2_0, // @[:@6.4]
  input  [1:0] io_selects_2_1, // @[:@6.4]
  input  [1:0] io_selects_3_0, // @[:@6.4]
  input  [1:0] io_selects_3_1, // @[:@6.4]
  input  [1:0] io_selects_4_0, // @[:@6.4]
  input  [1:0] io_selects_4_1, // @[:@6.4]
  input  [1:0] io_selects_5_0, // @[:@6.4]
  input  [1:0] io_selects_5_1, // @[:@6.4]
  input  [1:0] io_selects_6_0, // @[:@6.4]
  input  [1:0] io_selects_6_1, // @[:@6.4]
  input  [1:0] io_selects_7_0, // @[:@6.4]
  input  [1:0] io_selects_7_1, // @[:@6.4]
  input  [2:0] io_operation_0, // @[:@6.4]
  input  [2:0] io_operation_1, // @[:@6.4]
  input  [2:0] io_operation_2, // @[:@6.4]
  input  [2:0] io_operation_3, // @[:@6.4]
  input  [2:0] io_operation_4, // @[:@6.4]
  input  [2:0] io_operation_5, // @[:@6.4]
  input  [2:0] io_operation_6, // @[:@6.4]
  input  [2:0] io_operation_7, // @[:@6.4]
  input        io_inputs_0, // @[:@6.4]
  input        io_inputs_1, // @[:@6.4]
  input        io_inputs_2, // @[:@6.4]
  input        io_inputs_3, // @[:@6.4]
  output       io_outputs_0, // @[:@6.4]
  output       io_outputs_1, // @[:@6.4]
  output       io_outputs_2, // @[:@6.4]
  output       io_outputs_3, // @[:@6.4]
  output       io_outputs_4, // @[:@6.4]
  output       io_outputs_5, // @[:@6.4]
  output       io_outputs_6, // @[:@6.4]
  output       io_outputs_7 // @[:@6.4]
);
  wire  _GEN_1; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_2; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_3; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_5; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_6; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_7; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [1:0] _T_394; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire  _T_395; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@9.4]
  wire [1:0] _T_397; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@10.4]
  wire  _T_399; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@11.4]
  wire  _T_400; // @[Mux.scala 46:19:@12.4]
  wire  _T_401; // @[Mux.scala 46:16:@13.4]
  wire  _T_402; // @[Mux.scala 46:19:@14.4]
  wire [1:0] _T_403; // @[Mux.scala 46:16:@15.4]
  wire  _T_404; // @[Mux.scala 46:19:@16.4]
  wire [1:0] _T_405; // @[Mux.scala 46:16:@17.4]
  wire  _T_406; // @[Mux.scala 46:19:@18.4]
  wire [1:0] _T_407; // @[Mux.scala 46:16:@19.4]
  wire  _GEN_9; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_10; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_11; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_13; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_14; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_15; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [1:0] _T_411; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire  _T_412; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@21.4]
  wire [1:0] _T_414; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@22.4]
  wire  _T_416; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@23.4]
  wire  _T_417; // @[Mux.scala 46:19:@24.4]
  wire  _T_418; // @[Mux.scala 46:16:@25.4]
  wire  _T_419; // @[Mux.scala 46:19:@26.4]
  wire [1:0] _T_420; // @[Mux.scala 46:16:@27.4]
  wire  _T_421; // @[Mux.scala 46:19:@28.4]
  wire [1:0] _T_422; // @[Mux.scala 46:16:@29.4]
  wire  _T_423; // @[Mux.scala 46:19:@30.4]
  wire [1:0] _T_424; // @[Mux.scala 46:16:@31.4]
  wire  _GEN_17; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_18; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_19; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_21; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_22; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_23; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [1:0] _T_428; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire  _T_429; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@33.4]
  wire [1:0] _T_431; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@34.4]
  wire  _T_433; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@35.4]
  wire  _T_434; // @[Mux.scala 46:19:@36.4]
  wire  _T_435; // @[Mux.scala 46:16:@37.4]
  wire  _T_436; // @[Mux.scala 46:19:@38.4]
  wire [1:0] _T_437; // @[Mux.scala 46:16:@39.4]
  wire  _T_438; // @[Mux.scala 46:19:@40.4]
  wire [1:0] _T_439; // @[Mux.scala 46:16:@41.4]
  wire  _T_440; // @[Mux.scala 46:19:@42.4]
  wire [1:0] _T_441; // @[Mux.scala 46:16:@43.4]
  wire  _GEN_25; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_26; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_27; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_29; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_30; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_31; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [1:0] _T_445; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire  _T_446; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@45.4]
  wire [1:0] _T_448; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@46.4]
  wire  _T_450; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@47.4]
  wire  _T_451; // @[Mux.scala 46:19:@48.4]
  wire  _T_452; // @[Mux.scala 46:16:@49.4]
  wire  _T_453; // @[Mux.scala 46:19:@50.4]
  wire [1:0] _T_454; // @[Mux.scala 46:16:@51.4]
  wire  _T_455; // @[Mux.scala 46:19:@52.4]
  wire [1:0] _T_456; // @[Mux.scala 46:16:@53.4]
  wire  _T_457; // @[Mux.scala 46:19:@54.4]
  wire [1:0] _T_458; // @[Mux.scala 46:16:@55.4]
  wire  _GEN_33; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_34; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_35; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_37; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_38; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_39; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [1:0] _T_462; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire  _T_463; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@57.4]
  wire [1:0] _T_465; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@58.4]
  wire  _T_467; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@59.4]
  wire  _T_468; // @[Mux.scala 46:19:@60.4]
  wire  _T_469; // @[Mux.scala 46:16:@61.4]
  wire  _T_470; // @[Mux.scala 46:19:@62.4]
  wire [1:0] _T_471; // @[Mux.scala 46:16:@63.4]
  wire  _T_472; // @[Mux.scala 46:19:@64.4]
  wire [1:0] _T_473; // @[Mux.scala 46:16:@65.4]
  wire  _T_474; // @[Mux.scala 46:19:@66.4]
  wire [1:0] _T_475; // @[Mux.scala 46:16:@67.4]
  wire  _GEN_41; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_42; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_43; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_45; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_46; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_47; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [1:0] _T_479; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire  _T_480; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@69.4]
  wire [1:0] _T_482; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@70.4]
  wire  _T_484; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@71.4]
  wire  _T_485; // @[Mux.scala 46:19:@72.4]
  wire  _T_486; // @[Mux.scala 46:16:@73.4]
  wire  _T_487; // @[Mux.scala 46:19:@74.4]
  wire [1:0] _T_488; // @[Mux.scala 46:16:@75.4]
  wire  _T_489; // @[Mux.scala 46:19:@76.4]
  wire [1:0] _T_490; // @[Mux.scala 46:16:@77.4]
  wire  _T_491; // @[Mux.scala 46:19:@78.4]
  wire [1:0] _T_492; // @[Mux.scala 46:16:@79.4]
  wire  _GEN_49; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_50; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_51; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_53; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_54; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_55; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [1:0] _T_496; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire  _T_497; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@81.4]
  wire [1:0] _T_499; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@82.4]
  wire  _T_501; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@83.4]
  wire  _T_502; // @[Mux.scala 46:19:@84.4]
  wire  _T_503; // @[Mux.scala 46:16:@85.4]
  wire  _T_504; // @[Mux.scala 46:19:@86.4]
  wire [1:0] _T_505; // @[Mux.scala 46:16:@87.4]
  wire  _T_506; // @[Mux.scala 46:19:@88.4]
  wire [1:0] _T_507; // @[Mux.scala 46:16:@89.4]
  wire  _T_508; // @[Mux.scala 46:19:@90.4]
  wire [1:0] _T_509; // @[Mux.scala 46:16:@91.4]
  wire  _GEN_57; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_58; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_59; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_61; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_62; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_63; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [1:0] _T_513; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire  _T_514; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@93.4]
  wire [1:0] _T_516; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@94.4]
  wire  _T_518; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@95.4]
  wire  _T_519; // @[Mux.scala 46:19:@96.4]
  wire  _T_520; // @[Mux.scala 46:16:@97.4]
  wire  _T_521; // @[Mux.scala 46:19:@98.4]
  wire [1:0] _T_522; // @[Mux.scala 46:16:@99.4]
  wire  _T_523; // @[Mux.scala 46:19:@100.4]
  wire [1:0] _T_524; // @[Mux.scala 46:16:@101.4]
  wire  _T_525; // @[Mux.scala 46:19:@102.4]
  wire [1:0] _T_526; // @[Mux.scala 46:16:@103.4]
  assign _GEN_1 = 2'h1 == io_selects_0_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_2 = 2'h2 == io_selects_0_0 ? io_inputs_2 : _GEN_1; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_3 = 2'h3 == io_selects_0_0 ? io_inputs_3 : _GEN_2; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_5 = 2'h1 == io_selects_0_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_6 = 2'h2 == io_selects_0_1 ? io_inputs_2 : _GEN_5; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_7 = 2'h3 == io_selects_0_1 ? io_inputs_3 : _GEN_6; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _T_394 = _GEN_3 + _GEN_7; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _T_395 = _GEN_3 + _GEN_7; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@9.4]
  assign _T_397 = _GEN_3 * _GEN_7; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@10.4]
  assign _T_399 = _GEN_3 / _GEN_7; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@11.4]
  assign _T_400 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_401 = _T_400 ? _T_399 : 1'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_402 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_403 = _T_402 ? _T_397 : {{1'd0}, _T_401}; // @[Mux.scala 46:16:@15.4]
  assign _T_404 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_405 = _T_404 ? {{1'd0}, _T_395} : _T_403; // @[Mux.scala 46:16:@17.4]
  assign _T_406 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _T_407 = _T_406 ? {{1'd0}, _GEN_3} : _T_405; // @[Mux.scala 46:16:@19.4]
  assign _GEN_9 = 2'h1 == io_selects_1_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_10 = 2'h2 == io_selects_1_0 ? io_inputs_2 : _GEN_9; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_11 = 2'h3 == io_selects_1_0 ? io_inputs_3 : _GEN_10; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_13 = 2'h1 == io_selects_1_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_14 = 2'h2 == io_selects_1_1 ? io_inputs_2 : _GEN_13; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_15 = 2'h3 == io_selects_1_1 ? io_inputs_3 : _GEN_14; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _T_411 = _GEN_11 + _GEN_15; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _T_412 = _GEN_11 + _GEN_15; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@21.4]
  assign _T_414 = _GEN_11 * _GEN_15; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@22.4]
  assign _T_416 = _GEN_11 / _GEN_15; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@23.4]
  assign _T_417 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_418 = _T_417 ? _T_416 : 1'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_419 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_420 = _T_419 ? _T_414 : {{1'd0}, _T_418}; // @[Mux.scala 46:16:@27.4]
  assign _T_421 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_422 = _T_421 ? {{1'd0}, _T_412} : _T_420; // @[Mux.scala 46:16:@29.4]
  assign _T_423 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _T_424 = _T_423 ? {{1'd0}, _GEN_11} : _T_422; // @[Mux.scala 46:16:@31.4]
  assign _GEN_17 = 2'h1 == io_selects_2_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_18 = 2'h2 == io_selects_2_0 ? io_inputs_2 : _GEN_17; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_19 = 2'h3 == io_selects_2_0 ? io_inputs_3 : _GEN_18; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_21 = 2'h1 == io_selects_2_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_22 = 2'h2 == io_selects_2_1 ? io_inputs_2 : _GEN_21; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_23 = 2'h3 == io_selects_2_1 ? io_inputs_3 : _GEN_22; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _T_428 = _GEN_19 + _GEN_23; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _T_429 = _GEN_19 + _GEN_23; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@33.4]
  assign _T_431 = _GEN_19 * _GEN_23; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@34.4]
  assign _T_433 = _GEN_19 / _GEN_23; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@35.4]
  assign _T_434 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_435 = _T_434 ? _T_433 : 1'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_436 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_437 = _T_436 ? _T_431 : {{1'd0}, _T_435}; // @[Mux.scala 46:16:@39.4]
  assign _T_438 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_439 = _T_438 ? {{1'd0}, _T_429} : _T_437; // @[Mux.scala 46:16:@41.4]
  assign _T_440 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _T_441 = _T_440 ? {{1'd0}, _GEN_19} : _T_439; // @[Mux.scala 46:16:@43.4]
  assign _GEN_25 = 2'h1 == io_selects_3_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_26 = 2'h2 == io_selects_3_0 ? io_inputs_2 : _GEN_25; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_27 = 2'h3 == io_selects_3_0 ? io_inputs_3 : _GEN_26; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_29 = 2'h1 == io_selects_3_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_30 = 2'h2 == io_selects_3_1 ? io_inputs_2 : _GEN_29; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_31 = 2'h3 == io_selects_3_1 ? io_inputs_3 : _GEN_30; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _T_445 = _GEN_27 + _GEN_31; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _T_446 = _GEN_27 + _GEN_31; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@45.4]
  assign _T_448 = _GEN_27 * _GEN_31; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@46.4]
  assign _T_450 = _GEN_27 / _GEN_31; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@47.4]
  assign _T_451 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_452 = _T_451 ? _T_450 : 1'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_453 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_454 = _T_453 ? _T_448 : {{1'd0}, _T_452}; // @[Mux.scala 46:16:@51.4]
  assign _T_455 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_456 = _T_455 ? {{1'd0}, _T_446} : _T_454; // @[Mux.scala 46:16:@53.4]
  assign _T_457 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _T_458 = _T_457 ? {{1'd0}, _GEN_27} : _T_456; // @[Mux.scala 46:16:@55.4]
  assign _GEN_33 = 2'h1 == io_selects_4_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_34 = 2'h2 == io_selects_4_0 ? io_inputs_2 : _GEN_33; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_35 = 2'h3 == io_selects_4_0 ? io_inputs_3 : _GEN_34; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_37 = 2'h1 == io_selects_4_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_38 = 2'h2 == io_selects_4_1 ? io_inputs_2 : _GEN_37; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_39 = 2'h3 == io_selects_4_1 ? io_inputs_3 : _GEN_38; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _T_462 = _GEN_35 + _GEN_39; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _T_463 = _GEN_35 + _GEN_39; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@57.4]
  assign _T_465 = _GEN_35 * _GEN_39; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@58.4]
  assign _T_467 = _GEN_35 / _GEN_39; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@59.4]
  assign _T_468 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_469 = _T_468 ? _T_467 : 1'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_470 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_471 = _T_470 ? _T_465 : {{1'd0}, _T_469}; // @[Mux.scala 46:16:@63.4]
  assign _T_472 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_473 = _T_472 ? {{1'd0}, _T_463} : _T_471; // @[Mux.scala 46:16:@65.4]
  assign _T_474 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _T_475 = _T_474 ? {{1'd0}, _GEN_35} : _T_473; // @[Mux.scala 46:16:@67.4]
  assign _GEN_41 = 2'h1 == io_selects_5_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_42 = 2'h2 == io_selects_5_0 ? io_inputs_2 : _GEN_41; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_43 = 2'h3 == io_selects_5_0 ? io_inputs_3 : _GEN_42; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_45 = 2'h1 == io_selects_5_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_46 = 2'h2 == io_selects_5_1 ? io_inputs_2 : _GEN_45; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_47 = 2'h3 == io_selects_5_1 ? io_inputs_3 : _GEN_46; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _T_479 = _GEN_43 + _GEN_47; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _T_480 = _GEN_43 + _GEN_47; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@69.4]
  assign _T_482 = _GEN_43 * _GEN_47; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@70.4]
  assign _T_484 = _GEN_43 / _GEN_47; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@71.4]
  assign _T_485 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_486 = _T_485 ? _T_484 : 1'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_487 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_488 = _T_487 ? _T_482 : {{1'd0}, _T_486}; // @[Mux.scala 46:16:@75.4]
  assign _T_489 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_490 = _T_489 ? {{1'd0}, _T_480} : _T_488; // @[Mux.scala 46:16:@77.4]
  assign _T_491 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _T_492 = _T_491 ? {{1'd0}, _GEN_43} : _T_490; // @[Mux.scala 46:16:@79.4]
  assign _GEN_49 = 2'h1 == io_selects_6_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_50 = 2'h2 == io_selects_6_0 ? io_inputs_2 : _GEN_49; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_51 = 2'h3 == io_selects_6_0 ? io_inputs_3 : _GEN_50; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_53 = 2'h1 == io_selects_6_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_54 = 2'h2 == io_selects_6_1 ? io_inputs_2 : _GEN_53; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_55 = 2'h3 == io_selects_6_1 ? io_inputs_3 : _GEN_54; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _T_496 = _GEN_51 + _GEN_55; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _T_497 = _GEN_51 + _GEN_55; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@81.4]
  assign _T_499 = _GEN_51 * _GEN_55; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@82.4]
  assign _T_501 = _GEN_51 / _GEN_55; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@83.4]
  assign _T_502 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_503 = _T_502 ? _T_501 : 1'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_504 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_505 = _T_504 ? _T_499 : {{1'd0}, _T_503}; // @[Mux.scala 46:16:@87.4]
  assign _T_506 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_507 = _T_506 ? {{1'd0}, _T_497} : _T_505; // @[Mux.scala 46:16:@89.4]
  assign _T_508 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _T_509 = _T_508 ? {{1'd0}, _GEN_51} : _T_507; // @[Mux.scala 46:16:@91.4]
  assign _GEN_57 = 2'h1 == io_selects_7_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_58 = 2'h2 == io_selects_7_0 ? io_inputs_2 : _GEN_57; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_59 = 2'h3 == io_selects_7_0 ? io_inputs_3 : _GEN_58; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_61 = 2'h1 == io_selects_7_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_62 = 2'h2 == io_selects_7_1 ? io_inputs_2 : _GEN_61; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_63 = 2'h3 == io_selects_7_1 ? io_inputs_3 : _GEN_62; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _T_513 = _GEN_59 + _GEN_63; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _T_514 = _GEN_59 + _GEN_63; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 32:53:@93.4]
  assign _T_516 = _GEN_59 * _GEN_63; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 33:58:@94.4]
  assign _T_518 = _GEN_59 / _GEN_63; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 34:56:@95.4]
  assign _T_519 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_520 = _T_519 ? _T_518 : 1'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_521 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_522 = _T_521 ? _T_516 : {{1'd0}, _T_520}; // @[Mux.scala 46:16:@99.4]
  assign _T_523 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_524 = _T_523 ? {{1'd0}, _T_514} : _T_522; // @[Mux.scala 46:16:@101.4]
  assign _T_525 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign _T_526 = _T_525 ? {{1'd0}, _GEN_59} : _T_524; // @[Mux.scala 46:16:@103.4]
  assign io_outputs_0 = _T_407[0]; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 23:14:@104.4]
  assign io_outputs_1 = _T_424[0]; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 23:14:@105.4]
  assign io_outputs_2 = _T_441[0]; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 23:14:@106.4]
  assign io_outputs_3 = _T_458[0]; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 23:14:@107.4]
  assign io_outputs_4 = _T_475[0]; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 23:14:@108.4]
  assign io_outputs_5 = _T_492[0]; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 23:14:@109.4]
  assign io_outputs_6 = _T_509[0]; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 23:14:@110.4]
  assign io_outputs_7 = _T_526[0]; // @[MuxTest_width_1_inputs_4_outputs_8_pipeline_0s.scala 23:14:@111.4]
endmodule
