VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram7_256x32
  FOREIGN fakeram7_256x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 4.180 BY 67.200 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.096 0.024 0.120 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.960 0.024 0.984 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.824 0.024 1.848 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.688 0.024 2.712 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.552 0.024 3.576 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.416 0.024 4.440 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.280 0.024 5.304 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.144 0.024 6.168 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.008 0.024 7.032 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.872 0.024 7.896 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.736 0.024 8.760 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.600 0.024 9.624 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.464 0.024 10.488 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.328 0.024 11.352 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.192 0.024 12.216 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.056 0.024 13.080 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.920 0.024 13.944 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.784 0.024 14.808 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.648 0.024 15.672 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.512 0.024 16.536 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.376 0.024 17.400 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.240 0.024 18.264 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.104 0.024 19.128 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.968 0.024 19.992 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.832 0.024 20.856 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.696 0.024 21.720 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.560 0.024 22.584 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.424 0.024 23.448 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.288 0.024 24.312 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.152 0.024 25.176 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.016 0.024 26.040 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.880 0.024 26.904 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.408 0.024 27.432 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.272 0.024 28.296 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.136 0.024 29.160 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.000 0.024 30.024 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.864 0.024 30.888 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.728 0.024 31.752 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.592 0.024 32.616 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 33.456 0.024 33.480 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 34.320 0.024 34.344 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 35.184 0.024 35.208 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.048 0.024 36.072 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.912 0.024 36.936 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.776 0.024 37.800 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 38.640 0.024 38.664 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 39.504 0.024 39.528 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 40.368 0.024 40.392 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 41.232 0.024 41.256 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 42.096 0.024 42.120 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 42.960 0.024 42.984 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 43.824 0.024 43.848 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 44.688 0.024 44.712 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 45.552 0.024 45.576 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 46.416 0.024 46.440 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 47.280 0.024 47.304 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 48.144 0.024 48.168 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.008 0.024 49.032 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.872 0.024 49.896 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 50.736 0.024 50.760 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.600 0.024 51.624 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 52.464 0.024 52.488 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 53.328 0.024 53.352 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.192 0.024 54.216 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.720 0.024 54.744 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 55.584 0.024 55.608 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 56.448 0.024 56.472 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 57.312 0.024 57.336 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 58.176 0.024 58.200 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.040 0.024 59.064 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.904 0.024 59.928 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 60.768 0.024 60.792 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 61.296 0.024 61.320 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 62.160 0.024 62.184 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 63.024 0.024 63.048 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.048 4.084 0.144 ;
      RECT 0.096 0.816 4.084 0.912 ;
      RECT 0.096 1.584 4.084 1.680 ;
      RECT 0.096 2.352 4.084 2.448 ;
      RECT 0.096 3.120 4.084 3.216 ;
      RECT 0.096 3.888 4.084 3.984 ;
      RECT 0.096 4.656 4.084 4.752 ;
      RECT 0.096 5.424 4.084 5.520 ;
      RECT 0.096 6.192 4.084 6.288 ;
      RECT 0.096 6.960 4.084 7.056 ;
      RECT 0.096 7.728 4.084 7.824 ;
      RECT 0.096 8.496 4.084 8.592 ;
      RECT 0.096 9.264 4.084 9.360 ;
      RECT 0.096 10.032 4.084 10.128 ;
      RECT 0.096 10.800 4.084 10.896 ;
      RECT 0.096 11.568 4.084 11.664 ;
      RECT 0.096 12.336 4.084 12.432 ;
      RECT 0.096 13.104 4.084 13.200 ;
      RECT 0.096 13.872 4.084 13.968 ;
      RECT 0.096 14.640 4.084 14.736 ;
      RECT 0.096 15.408 4.084 15.504 ;
      RECT 0.096 16.176 4.084 16.272 ;
      RECT 0.096 16.944 4.084 17.040 ;
      RECT 0.096 17.712 4.084 17.808 ;
      RECT 0.096 18.480 4.084 18.576 ;
      RECT 0.096 19.248 4.084 19.344 ;
      RECT 0.096 20.016 4.084 20.112 ;
      RECT 0.096 20.784 4.084 20.880 ;
      RECT 0.096 21.552 4.084 21.648 ;
      RECT 0.096 22.320 4.084 22.416 ;
      RECT 0.096 23.088 4.084 23.184 ;
      RECT 0.096 23.856 4.084 23.952 ;
      RECT 0.096 24.624 4.084 24.720 ;
      RECT 0.096 25.392 4.084 25.488 ;
      RECT 0.096 26.160 4.084 26.256 ;
      RECT 0.096 26.928 4.084 27.024 ;
      RECT 0.096 27.696 4.084 27.792 ;
      RECT 0.096 28.464 4.084 28.560 ;
      RECT 0.096 29.232 4.084 29.328 ;
      RECT 0.096 30.000 4.084 30.096 ;
      RECT 0.096 30.768 4.084 30.864 ;
      RECT 0.096 31.536 4.084 31.632 ;
      RECT 0.096 32.304 4.084 32.400 ;
      RECT 0.096 33.072 4.084 33.168 ;
      RECT 0.096 33.840 4.084 33.936 ;
      RECT 0.096 34.608 4.084 34.704 ;
      RECT 0.096 35.376 4.084 35.472 ;
      RECT 0.096 36.144 4.084 36.240 ;
      RECT 0.096 36.912 4.084 37.008 ;
      RECT 0.096 37.680 4.084 37.776 ;
      RECT 0.096 38.448 4.084 38.544 ;
      RECT 0.096 39.216 4.084 39.312 ;
      RECT 0.096 39.984 4.084 40.080 ;
      RECT 0.096 40.752 4.084 40.848 ;
      RECT 0.096 41.520 4.084 41.616 ;
      RECT 0.096 42.288 4.084 42.384 ;
      RECT 0.096 43.056 4.084 43.152 ;
      RECT 0.096 43.824 4.084 43.920 ;
      RECT 0.096 44.592 4.084 44.688 ;
      RECT 0.096 45.360 4.084 45.456 ;
      RECT 0.096 46.128 4.084 46.224 ;
      RECT 0.096 46.896 4.084 46.992 ;
      RECT 0.096 47.664 4.084 47.760 ;
      RECT 0.096 48.432 4.084 48.528 ;
      RECT 0.096 49.200 4.084 49.296 ;
      RECT 0.096 49.968 4.084 50.064 ;
      RECT 0.096 50.736 4.084 50.832 ;
      RECT 0.096 51.504 4.084 51.600 ;
      RECT 0.096 52.272 4.084 52.368 ;
      RECT 0.096 53.040 4.084 53.136 ;
      RECT 0.096 53.808 4.084 53.904 ;
      RECT 0.096 54.576 4.084 54.672 ;
      RECT 0.096 55.344 4.084 55.440 ;
      RECT 0.096 56.112 4.084 56.208 ;
      RECT 0.096 56.880 4.084 56.976 ;
      RECT 0.096 57.648 4.084 57.744 ;
      RECT 0.096 58.416 4.084 58.512 ;
      RECT 0.096 59.184 4.084 59.280 ;
      RECT 0.096 59.952 4.084 60.048 ;
      RECT 0.096 60.720 4.084 60.816 ;
      RECT 0.096 61.488 4.084 61.584 ;
      RECT 0.096 62.256 4.084 62.352 ;
      RECT 0.096 63.024 4.084 63.120 ;
      RECT 0.096 63.792 4.084 63.888 ;
      RECT 0.096 64.560 4.084 64.656 ;
      RECT 0.096 65.328 4.084 65.424 ;
      RECT 0.096 66.096 4.084 66.192 ;
      RECT 0.096 66.864 4.084 66.960 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.096 0.432 4.084 0.528 ;
      RECT 0.096 1.200 4.084 1.296 ;
      RECT 0.096 1.968 4.084 2.064 ;
      RECT 0.096 2.736 4.084 2.832 ;
      RECT 0.096 3.504 4.084 3.600 ;
      RECT 0.096 4.272 4.084 4.368 ;
      RECT 0.096 5.040 4.084 5.136 ;
      RECT 0.096 5.808 4.084 5.904 ;
      RECT 0.096 6.576 4.084 6.672 ;
      RECT 0.096 7.344 4.084 7.440 ;
      RECT 0.096 8.112 4.084 8.208 ;
      RECT 0.096 8.880 4.084 8.976 ;
      RECT 0.096 9.648 4.084 9.744 ;
      RECT 0.096 10.416 4.084 10.512 ;
      RECT 0.096 11.184 4.084 11.280 ;
      RECT 0.096 11.952 4.084 12.048 ;
      RECT 0.096 12.720 4.084 12.816 ;
      RECT 0.096 13.488 4.084 13.584 ;
      RECT 0.096 14.256 4.084 14.352 ;
      RECT 0.096 15.024 4.084 15.120 ;
      RECT 0.096 15.792 4.084 15.888 ;
      RECT 0.096 16.560 4.084 16.656 ;
      RECT 0.096 17.328 4.084 17.424 ;
      RECT 0.096 18.096 4.084 18.192 ;
      RECT 0.096 18.864 4.084 18.960 ;
      RECT 0.096 19.632 4.084 19.728 ;
      RECT 0.096 20.400 4.084 20.496 ;
      RECT 0.096 21.168 4.084 21.264 ;
      RECT 0.096 21.936 4.084 22.032 ;
      RECT 0.096 22.704 4.084 22.800 ;
      RECT 0.096 23.472 4.084 23.568 ;
      RECT 0.096 24.240 4.084 24.336 ;
      RECT 0.096 25.008 4.084 25.104 ;
      RECT 0.096 25.776 4.084 25.872 ;
      RECT 0.096 26.544 4.084 26.640 ;
      RECT 0.096 27.312 4.084 27.408 ;
      RECT 0.096 28.080 4.084 28.176 ;
      RECT 0.096 28.848 4.084 28.944 ;
      RECT 0.096 29.616 4.084 29.712 ;
      RECT 0.096 30.384 4.084 30.480 ;
      RECT 0.096 31.152 4.084 31.248 ;
      RECT 0.096 31.920 4.084 32.016 ;
      RECT 0.096 32.688 4.084 32.784 ;
      RECT 0.096 33.456 4.084 33.552 ;
      RECT 0.096 34.224 4.084 34.320 ;
      RECT 0.096 34.992 4.084 35.088 ;
      RECT 0.096 35.760 4.084 35.856 ;
      RECT 0.096 36.528 4.084 36.624 ;
      RECT 0.096 37.296 4.084 37.392 ;
      RECT 0.096 38.064 4.084 38.160 ;
      RECT 0.096 38.832 4.084 38.928 ;
      RECT 0.096 39.600 4.084 39.696 ;
      RECT 0.096 40.368 4.084 40.464 ;
      RECT 0.096 41.136 4.084 41.232 ;
      RECT 0.096 41.904 4.084 42.000 ;
      RECT 0.096 42.672 4.084 42.768 ;
      RECT 0.096 43.440 4.084 43.536 ;
      RECT 0.096 44.208 4.084 44.304 ;
      RECT 0.096 44.976 4.084 45.072 ;
      RECT 0.096 45.744 4.084 45.840 ;
      RECT 0.096 46.512 4.084 46.608 ;
      RECT 0.096 47.280 4.084 47.376 ;
      RECT 0.096 48.048 4.084 48.144 ;
      RECT 0.096 48.816 4.084 48.912 ;
      RECT 0.096 49.584 4.084 49.680 ;
      RECT 0.096 50.352 4.084 50.448 ;
      RECT 0.096 51.120 4.084 51.216 ;
      RECT 0.096 51.888 4.084 51.984 ;
      RECT 0.096 52.656 4.084 52.752 ;
      RECT 0.096 53.424 4.084 53.520 ;
      RECT 0.096 54.192 4.084 54.288 ;
      RECT 0.096 54.960 4.084 55.056 ;
      RECT 0.096 55.728 4.084 55.824 ;
      RECT 0.096 56.496 4.084 56.592 ;
      RECT 0.096 57.264 4.084 57.360 ;
      RECT 0.096 58.032 4.084 58.128 ;
      RECT 0.096 58.800 4.084 58.896 ;
      RECT 0.096 59.568 4.084 59.664 ;
      RECT 0.096 60.336 4.084 60.432 ;
      RECT 0.096 61.104 4.084 61.200 ;
      RECT 0.096 61.872 4.084 61.968 ;
      RECT 0.096 62.640 4.084 62.736 ;
      RECT 0.096 63.408 4.084 63.504 ;
      RECT 0.096 64.176 4.084 64.272 ;
      RECT 0.096 64.944 4.084 65.040 ;
      RECT 0.096 65.712 4.084 65.808 ;
      RECT 0.096 66.480 4.084 66.576 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 4.180 67.200 ;
    LAYER M2 ;
    RECT 0 0 4.180 67.200 ;
    LAYER M3 ;
    RECT 0 0 4.180 67.200 ;
    LAYER M4 ;
    RECT 0.024 0 0.096 67.200 ;
    RECT 4.084 0 4.180 67.200 ;
    RECT 0.096 0.000 4.084 0.048 ;
    RECT 0.096 0.144 4.084 0.432 ;
    RECT 0.096 0.528 4.084 0.816 ;
    RECT 0.096 0.912 4.084 1.200 ;
    RECT 0.096 1.296 4.084 1.584 ;
    RECT 0.096 1.680 4.084 1.968 ;
    RECT 0.096 2.064 4.084 2.352 ;
    RECT 0.096 2.448 4.084 2.736 ;
    RECT 0.096 2.832 4.084 3.120 ;
    RECT 0.096 3.216 4.084 3.504 ;
    RECT 0.096 3.600 4.084 3.888 ;
    RECT 0.096 3.984 4.084 4.272 ;
    RECT 0.096 4.368 4.084 4.656 ;
    RECT 0.096 4.752 4.084 5.040 ;
    RECT 0.096 5.136 4.084 5.424 ;
    RECT 0.096 5.520 4.084 5.808 ;
    RECT 0.096 5.904 4.084 6.192 ;
    RECT 0.096 6.288 4.084 6.576 ;
    RECT 0.096 6.672 4.084 6.960 ;
    RECT 0.096 7.056 4.084 7.344 ;
    RECT 0.096 7.440 4.084 7.728 ;
    RECT 0.096 7.824 4.084 8.112 ;
    RECT 0.096 8.208 4.084 8.496 ;
    RECT 0.096 8.592 4.084 8.880 ;
    RECT 0.096 8.976 4.084 9.264 ;
    RECT 0.096 9.360 4.084 9.648 ;
    RECT 0.096 9.744 4.084 10.032 ;
    RECT 0.096 10.128 4.084 10.416 ;
    RECT 0.096 10.512 4.084 10.800 ;
    RECT 0.096 10.896 4.084 11.184 ;
    RECT 0.096 11.280 4.084 11.568 ;
    RECT 0.096 11.664 4.084 11.952 ;
    RECT 0.096 12.048 4.084 12.336 ;
    RECT 0.096 12.432 4.084 12.720 ;
    RECT 0.096 12.816 4.084 13.104 ;
    RECT 0.096 13.200 4.084 13.488 ;
    RECT 0.096 13.584 4.084 13.872 ;
    RECT 0.096 13.968 4.084 14.256 ;
    RECT 0.096 14.352 4.084 14.640 ;
    RECT 0.096 14.736 4.084 15.024 ;
    RECT 0.096 15.120 4.084 15.408 ;
    RECT 0.096 15.504 4.084 15.792 ;
    RECT 0.096 15.888 4.084 16.176 ;
    RECT 0.096 16.272 4.084 16.560 ;
    RECT 0.096 16.656 4.084 16.944 ;
    RECT 0.096 17.040 4.084 17.328 ;
    RECT 0.096 17.424 4.084 17.712 ;
    RECT 0.096 17.808 4.084 18.096 ;
    RECT 0.096 18.192 4.084 18.480 ;
    RECT 0.096 18.576 4.084 18.864 ;
    RECT 0.096 18.960 4.084 19.248 ;
    RECT 0.096 19.344 4.084 19.632 ;
    RECT 0.096 19.728 4.084 20.016 ;
    RECT 0.096 20.112 4.084 20.400 ;
    RECT 0.096 20.496 4.084 20.784 ;
    RECT 0.096 20.880 4.084 21.168 ;
    RECT 0.096 21.264 4.084 21.552 ;
    RECT 0.096 21.648 4.084 21.936 ;
    RECT 0.096 22.032 4.084 22.320 ;
    RECT 0.096 22.416 4.084 22.704 ;
    RECT 0.096 22.800 4.084 23.088 ;
    RECT 0.096 23.184 4.084 23.472 ;
    RECT 0.096 23.568 4.084 23.856 ;
    RECT 0.096 23.952 4.084 24.240 ;
    RECT 0.096 24.336 4.084 24.624 ;
    RECT 0.096 24.720 4.084 25.008 ;
    RECT 0.096 25.104 4.084 25.392 ;
    RECT 0.096 25.488 4.084 25.776 ;
    RECT 0.096 25.872 4.084 26.160 ;
    RECT 0.096 26.256 4.084 26.544 ;
    RECT 0.096 26.640 4.084 26.928 ;
    RECT 0.096 27.024 4.084 27.312 ;
    RECT 0.096 27.408 4.084 27.696 ;
    RECT 0.096 27.792 4.084 28.080 ;
    RECT 0.096 28.176 4.084 28.464 ;
    RECT 0.096 28.560 4.084 28.848 ;
    RECT 0.096 28.944 4.084 29.232 ;
    RECT 0.096 29.328 4.084 29.616 ;
    RECT 0.096 29.712 4.084 30.000 ;
    RECT 0.096 30.096 4.084 30.384 ;
    RECT 0.096 30.480 4.084 30.768 ;
    RECT 0.096 30.864 4.084 31.152 ;
    RECT 0.096 31.248 4.084 31.536 ;
    RECT 0.096 31.632 4.084 31.920 ;
    RECT 0.096 32.016 4.084 32.304 ;
    RECT 0.096 32.400 4.084 32.688 ;
    RECT 0.096 32.784 4.084 33.072 ;
    RECT 0.096 33.168 4.084 33.456 ;
    RECT 0.096 33.552 4.084 33.840 ;
    RECT 0.096 33.936 4.084 34.224 ;
    RECT 0.096 34.320 4.084 34.608 ;
    RECT 0.096 34.704 4.084 34.992 ;
    RECT 0.096 35.088 4.084 35.376 ;
    RECT 0.096 35.472 4.084 35.760 ;
    RECT 0.096 35.856 4.084 36.144 ;
    RECT 0.096 36.240 4.084 36.528 ;
    RECT 0.096 36.624 4.084 36.912 ;
    RECT 0.096 37.008 4.084 37.296 ;
    RECT 0.096 37.392 4.084 37.680 ;
    RECT 0.096 37.776 4.084 38.064 ;
    RECT 0.096 38.160 4.084 38.448 ;
    RECT 0.096 38.544 4.084 38.832 ;
    RECT 0.096 38.928 4.084 39.216 ;
    RECT 0.096 39.312 4.084 39.600 ;
    RECT 0.096 39.696 4.084 39.984 ;
    RECT 0.096 40.080 4.084 40.368 ;
    RECT 0.096 40.464 4.084 40.752 ;
    RECT 0.096 40.848 4.084 41.136 ;
    RECT 0.096 41.232 4.084 41.520 ;
    RECT 0.096 41.616 4.084 41.904 ;
    RECT 0.096 42.000 4.084 42.288 ;
    RECT 0.096 42.384 4.084 42.672 ;
    RECT 0.096 42.768 4.084 43.056 ;
    RECT 0.096 43.152 4.084 43.440 ;
    RECT 0.096 43.536 4.084 43.824 ;
    RECT 0.096 43.920 4.084 44.208 ;
    RECT 0.096 44.304 4.084 44.592 ;
    RECT 0.096 44.688 4.084 44.976 ;
    RECT 0.096 45.072 4.084 45.360 ;
    RECT 0.096 45.456 4.084 45.744 ;
    RECT 0.096 45.840 4.084 46.128 ;
    RECT 0.096 46.224 4.084 46.512 ;
    RECT 0.096 46.608 4.084 46.896 ;
    RECT 0.096 46.992 4.084 47.280 ;
    RECT 0.096 47.376 4.084 47.664 ;
    RECT 0.096 47.760 4.084 48.048 ;
    RECT 0.096 48.144 4.084 48.432 ;
    RECT 0.096 48.528 4.084 48.816 ;
    RECT 0.096 48.912 4.084 49.200 ;
    RECT 0.096 49.296 4.084 49.584 ;
    RECT 0.096 49.680 4.084 49.968 ;
    RECT 0.096 50.064 4.084 50.352 ;
    RECT 0.096 50.448 4.084 50.736 ;
    RECT 0.096 50.832 4.084 51.120 ;
    RECT 0.096 51.216 4.084 51.504 ;
    RECT 0.096 51.600 4.084 51.888 ;
    RECT 0.096 51.984 4.084 52.272 ;
    RECT 0.096 52.368 4.084 52.656 ;
    RECT 0.096 52.752 4.084 53.040 ;
    RECT 0.096 53.136 4.084 53.424 ;
    RECT 0.096 53.520 4.084 53.808 ;
    RECT 0.096 53.904 4.084 54.192 ;
    RECT 0.096 54.288 4.084 54.576 ;
    RECT 0.096 54.672 4.084 54.960 ;
    RECT 0.096 55.056 4.084 55.344 ;
    RECT 0.096 55.440 4.084 55.728 ;
    RECT 0.096 55.824 4.084 56.112 ;
    RECT 0.096 56.208 4.084 56.496 ;
    RECT 0.096 56.592 4.084 56.880 ;
    RECT 0.096 56.976 4.084 57.264 ;
    RECT 0.096 57.360 4.084 57.648 ;
    RECT 0.096 57.744 4.084 58.032 ;
    RECT 0.096 58.128 4.084 58.416 ;
    RECT 0.096 58.512 4.084 58.800 ;
    RECT 0.096 58.896 4.084 59.184 ;
    RECT 0.096 59.280 4.084 59.568 ;
    RECT 0.096 59.664 4.084 59.952 ;
    RECT 0.096 60.048 4.084 60.336 ;
    RECT 0.096 60.432 4.084 60.720 ;
    RECT 0.096 60.816 4.084 61.104 ;
    RECT 0.096 61.200 4.084 61.488 ;
    RECT 0.096 61.584 4.084 61.872 ;
    RECT 0.096 61.968 4.084 62.256 ;
    RECT 0.096 62.352 4.084 62.640 ;
    RECT 0.096 62.736 4.084 63.024 ;
    RECT 0.096 63.120 4.084 63.408 ;
    RECT 0.096 63.504 4.084 63.792 ;
    RECT 0.096 63.888 4.084 64.176 ;
    RECT 0.096 64.272 4.084 64.560 ;
    RECT 0.096 64.656 4.084 64.944 ;
    RECT 0.096 65.040 4.084 65.328 ;
    RECT 0.096 65.424 4.084 65.712 ;
    RECT 0.096 65.808 4.084 66.096 ;
    RECT 0.096 66.192 4.084 66.480 ;
    RECT 0.096 66.576 4.084 66.864 ;
    RECT 0.096 66.960 4.084 67.200 ;
    RECT 0 0.000 0.024 0.096 ;
    RECT 0 0.120 0.024 0.960 ;
    RECT 0 0.984 0.024 1.824 ;
    RECT 0 1.848 0.024 2.688 ;
    RECT 0 2.712 0.024 3.552 ;
    RECT 0 3.576 0.024 4.416 ;
    RECT 0 4.440 0.024 5.280 ;
    RECT 0 5.304 0.024 6.144 ;
    RECT 0 6.168 0.024 7.008 ;
    RECT 0 7.032 0.024 7.872 ;
    RECT 0 7.896 0.024 8.736 ;
    RECT 0 8.760 0.024 9.600 ;
    RECT 0 9.624 0.024 10.464 ;
    RECT 0 10.488 0.024 11.328 ;
    RECT 0 11.352 0.024 12.192 ;
    RECT 0 12.216 0.024 13.056 ;
    RECT 0 13.080 0.024 13.920 ;
    RECT 0 13.944 0.024 14.784 ;
    RECT 0 14.808 0.024 15.648 ;
    RECT 0 15.672 0.024 16.512 ;
    RECT 0 16.536 0.024 17.376 ;
    RECT 0 17.400 0.024 18.240 ;
    RECT 0 18.264 0.024 19.104 ;
    RECT 0 19.128 0.024 19.968 ;
    RECT 0 19.992 0.024 20.832 ;
    RECT 0 20.856 0.024 21.696 ;
    RECT 0 21.720 0.024 22.560 ;
    RECT 0 22.584 0.024 23.424 ;
    RECT 0 23.448 0.024 24.288 ;
    RECT 0 24.312 0.024 25.152 ;
    RECT 0 25.176 0.024 26.016 ;
    RECT 0 26.040 0.024 26.880 ;
    RECT 0 26.904 0.024 27.408 ;
    RECT 0 27.432 0.024 28.272 ;
    RECT 0 28.296 0.024 29.136 ;
    RECT 0 29.160 0.024 30.000 ;
    RECT 0 30.024 0.024 30.864 ;
    RECT 0 30.888 0.024 31.728 ;
    RECT 0 31.752 0.024 32.592 ;
    RECT 0 32.616 0.024 33.456 ;
    RECT 0 33.480 0.024 34.320 ;
    RECT 0 34.344 0.024 35.184 ;
    RECT 0 35.208 0.024 36.048 ;
    RECT 0 36.072 0.024 36.912 ;
    RECT 0 36.936 0.024 37.776 ;
    RECT 0 37.800 0.024 38.640 ;
    RECT 0 38.664 0.024 39.504 ;
    RECT 0 39.528 0.024 40.368 ;
    RECT 0 40.392 0.024 41.232 ;
    RECT 0 41.256 0.024 42.096 ;
    RECT 0 42.120 0.024 42.960 ;
    RECT 0 42.984 0.024 43.824 ;
    RECT 0 43.848 0.024 44.688 ;
    RECT 0 44.712 0.024 45.552 ;
    RECT 0 45.576 0.024 46.416 ;
    RECT 0 46.440 0.024 47.280 ;
    RECT 0 47.304 0.024 48.144 ;
    RECT 0 48.168 0.024 49.008 ;
    RECT 0 49.032 0.024 49.872 ;
    RECT 0 49.896 0.024 50.736 ;
    RECT 0 50.760 0.024 51.600 ;
    RECT 0 51.624 0.024 52.464 ;
    RECT 0 52.488 0.024 53.328 ;
    RECT 0 53.352 0.024 54.192 ;
    RECT 0 54.216 0.024 54.720 ;
    RECT 0 54.744 0.024 55.584 ;
    RECT 0 55.608 0.024 56.448 ;
    RECT 0 56.472 0.024 57.312 ;
    RECT 0 57.336 0.024 58.176 ;
    RECT 0 58.200 0.024 59.040 ;
    RECT 0 59.064 0.024 59.904 ;
    RECT 0 59.928 0.024 60.768 ;
    RECT 0 60.792 0.024 61.632 ;
    RECT 0 61.656 0.024 62.496 ;
    RECT 0 62.520 0.024 63.360 ;
    RECT 0 63.384 0.024 64.224 ;
    RECT 0 64.248 0.024 65.088 ;
    RECT 0 65.112 0.024 65.952 ;
    RECT 0 65.976 0.024 66.816 ;
    RECT 0 66.840 0.024 67.680 ;
    RECT 0 67.704 0.024 68.544 ;
    RECT 0 68.568 0.024 69.408 ;
    RECT 0 69.432 0.024 70.272 ;
    RECT 0 70.296 0.024 71.136 ;
    RECT 0 71.160 0.024 72.000 ;
    RECT 0 72.024 0.024 72.864 ;
    RECT 0 72.888 0.024 73.728 ;
    RECT 0 73.752 0.024 74.592 ;
    RECT 0 74.616 0.024 75.456 ;
    RECT 0 75.480 0.024 76.320 ;
    RECT 0 76.344 0.024 77.184 ;
    RECT 0 77.208 0.024 78.048 ;
    RECT 0 78.072 0.024 78.912 ;
    RECT 0 78.936 0.024 79.776 ;
    RECT 0 79.800 0.024 80.640 ;
    RECT 0 80.664 0.024 81.504 ;
    RECT 0 81.528 0.024 82.032 ;
    RECT 0 82.056 0.024 82.896 ;
    RECT 0 82.920 0.024 83.760 ;
    RECT 0 83.784 0.024 84.624 ;
    RECT 0 84.648 0.024 85.488 ;
    RECT 0 85.512 0.024 86.352 ;
    RECT 0 86.376 0.024 87.216 ;
    RECT 0 87.240 0.024 88.080 ;
    RECT 0 88.104 0.024 88.608 ;
    RECT 0 88.632 0.024 89.472 ;
    RECT 0 89.496 0.024 90.336 ;
    RECT 0 90.360 0.024 67.200 ;
    LAYER OVERLAP ;
    RECT 0 0 4.180 67.200 ;
  END
END fakeram7_256x32

END LIBRARY
