# BSD 3-Clause License
# 
# Copyright 2020 Lawrence T. Clark, Vinay Vashishtha, or Arizona State
# University
# 
# Redistribution and use in source and binary forms, with or without
# modification, are permitted provided that the following conditions are met:
# 
# 1. Redistributions of source code must retain the above copyright notice,
# this list of conditions and the following disclaimer.
# 
# 2. Redistributions in binary form must reproduce the above copyright
# notice, this list of conditions and the following disclaimer in the
# documentation and/or other materials provided with the distribution.
# 
# 3. Neither the name of the copyright holder nor the names of its
# contributors may be used to endorse or promote products derived from this
# software without specific prior written permission.
# 
# THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
# AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
# IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
# ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
# LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
# CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
# SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
# INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
# CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
# ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
# POSSIBILITY OF SUCH DAMAGE.

VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
CLEARANCEMEASURE EUCLIDEAN ; 

UNITS 
DATABASE MICRONS 4000 ; 
END UNITS 
MANUFACTURINGGRID 0.001 ; 

PROPERTYDEFINITIONS 
LAYER LEF58_TYPE STRING ; 
LAYER LEF58_PITCH STRING ; 
LAYER LEF58_GAP STRING ; 
LAYER LEF58_EOLKEEPOUT STRING ; 
# LAYER LEF58_SPACING STRING ; 
LAYER LEF58_CORNERSPACING STRING ; 
LAYER LEF58_WIDTHTABLE STRING ; 
LAYER LEF58_CUTCLASS STRING ; 
LAYER LEF58_SPACINGTABLE STRING ; 
LAYER LEF58_ENCLOSURE STRING ; 
LAYER LEF58_RIGHTWAYONGRIDONLY STRING ; 
LAYER LEF58_RECTONLY STRING ; 
END PROPERTYDEFINITIONS 

LAYER OVERLAP 
TYPE OVERLAP ; 
END OVERLAP 

LAYER nwell 
TYPE MASTERSLICE ; 
PROPERTY LEF58_TYPE "TYPE NWELL ;" ; 
END nwell 

LAYER pwell 
TYPE MASTERSLICE ; 
PROPERTY LEF58_TYPE "TYPE PWELL ;" ; 
END pwell 

LAYER Gate 
TYPE MASTERSLICE ; 
END Gate 

LAYER Active 
TYPE MASTERSLICE ; 
END Active 

LAYER V0 
TYPE CUT ; 
SPACING 0.018 ; 
WIDTH 0.018 ; 
END V0 

LAYER M1 
TYPE ROUTING ; 
DIRECTION VERTICAL ; 
PITCH 0.036 ; 
WIDTH 0.018 ; 
SPACING 0.018 ; 
AREA 0.000666 ; # Min Area # This should ideally be 16x not 4x as each dimension is scaled up by 1 
# we only allow landing on pins (set in router) so area should not matter 
SPACING 0.018 RANGE 0.036 1 ; # This rule is redundant with the SPACING rule 

PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.01825 EXTENSION 0 0 0.031 ;" ; # Tip to Tip Spacing 

PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERONLY 0.01 WIDTH 0.018 SPACING 0.018 ;" ; 
OFFSET 0 ; 

END M1 

LAYER V1 
TYPE CUT ; 
SPACING 0.018 ; # unlike generate, this is really spacing, not center to center. 
WIDTH 0.018 ; 
END V1 

LAYER M2 
TYPE ROUTING ; 
DIRECTION HORIZONTAL ; 
WIDTH 0.018 ; # Min Width 
SPACING 0.018 ; # Min Spacing 

OFFSET -0.27 ; 

# MINSIZE is set so that the minimum lenght of a segment is 36nm. At the proper rule size of 
# 31nm, the lines can't be minimum space. This causes DRCs (like crazy). Same for M3 
# MINSIZE 0.028 0.018 ; 
# area is adjusted to match this (Nanoroute requires both AREA and MINSIZE) 

AREA 0.000666 ; 
MINSIZE 0.037 0.018 ; 

PITCH 0.045 0.036 ; 

# this enforces the correct routing tracks on M2 with wide M2 power rails 

PROPERTY LEF58_PITCH " 
PITCH 0.036 FIRSTLASTPITCH 0.045 
; 
" ; 

# this checks for distance in any direction so is not correct 
# 0.0175 is to avoid conflicts with the adjacent lines. This should be caught by CORNERSPACING below 
# SPACING 0.031 ENDOFLINE 0.025 WITHIN 0.0175 ; 

# SWK
# PROPERTY LEF58_SPACING 
# " SPACING 0.018 ENDOFLINE 0.025 WITHIN 0.02 ENDTOEND 0.031 
# PARALLELEDGE 0.025 WITHIN 0.02 ; " ; 
SPACING 0.031 ENDOFLINE 0.025 WITHIN 0.02 PARALLELEDGE 0.025 WITHIN 0.02 ;

PROPERTY LEF58_EOLKEEPOUT " 
EOLKEEPOUT 0.025 EXTENSION 0 0.0125 0.031 CORNERONLY ; 
" ; 

PROPERTY LEF58_CORNERSPACING " 
CORNERSPACING CONVEXCORNER WIDTH 0 SPACING 0.02 ; 
" ; # CORNER to CORNER SPACING Rule 

# Originally no width table for M2 since it is the follow rails. 
# They can be 1x or 2x (2x causes DRCs on SAV V1). However, this seems to allow a double width M2 
# on vias, which violates. Thus, this is added. Note that wide power follow rails will violate. 

PROPERTY LEF58_WIDTHTABLE " 
WIDTHTABLE 0.018 0.09 0.162 0.234 0.306 0.378 ; 
" ; 

PROPERTY LEF58_RIGHTWAYONGRIDONLY " 
RIGHTWAYONGRIDONLY ; 
" ; 

PROPERTY LEF58_RECTONLY " 
RECTONLY ; 
" ; 

END M2 

LAYER V2 
TYPE CUT ; 
SPACING 0.018 ; 
WIDTH 0.018 ; 
END V2 

LAYER M3 
TYPE ROUTING ; 
DIRECTION VERTICAL ; 
PITCH 0.036 ; 
OFFSET 0 ; 
WIDTH 0.018 ; # Min Width 
SPACING 0.018 ; # Min Spacing 

# MINSIZE is set so that the minimum lenght of a segment is 36nm. At the proper rule size of 
# 31nm, the lines can't be minimum space. This causes DRCs (like crazy). Same for M2 
# MINSIZE 0.028 0.018 ; 
# area is adjusted to match this (Nanoroute requires both AREA and MINSIZE) 

AREA 0.000666 ; 
MINSIZE 0.037 0.018 ; 

# SWK
# PROPERTY LEF58_SPACING 
# " SPACING 0.018 ENDOFLINE 0.025 WITHIN 0.0125 ENDTOEND 0.031 
# PARALLELEDGE 0.025 WITHIN 0.02 ; " ; 
SPACING 0.031 ENDOFLINE 0.025 WITHIN 0.0125 PARALLELEDGE 0.025 WITHIN 0.02 ;

PROPERTY LEF58_EOLKEEPOUT " 
EOLKEEPOUT 0.025 EXTENSION 0 0.0125 0.031 CORNERONLY ; 
" ; 

PROPERTY LEF58_CORNERSPACING " 
CORNERSPACING CONVEXCORNER WIDTH 0 SPACING 0.02 
; 
" ; # CORNER to CORNER SPACING Rule 

# to make the special route widths integer values of the tracks, i.e., 0.25, 1.25, 2.25, 3.25 min widths 
# the widths should be calculated in the APR tool, since viaGen does not seem to respect these 

PROPERTY LEF58_WIDTHTABLE 
" WIDTHTABLE 0.018 0.09 0.162 0.234 0.306 0.378 ; " ; 

PROPERTY LEF58_RIGHTWAYONGRIDONLY " 
RIGHTWAYONGRIDONLY ; 
" ; 

PROPERTY LEF58_RECTONLY " 
RECTONLY ; 
" ; 

END M3 

LAYER V3 
TYPE CUT ; 
#SPACING 0.018 ; 
WIDTH 0.018 ; 

# different format to allow long vias for SAV power connections 

PROPERTY LEF58_CUTCLASS " 
CUTCLASS V3       WIDTH 0.018 LENGTH 0.024 CUTS 0.25 ; 
CUTCLASS V3_0p480 WIDTH 0.018 LENGTH 0.12 CUTS 1 ; 
CUTCLASS V3_0p864 WIDTH 0.018 LENGTH 0.216 CUTS 2 ; 
" ; 

#PROPERTY LEF58_SPACINGTABLE " 
#SPACINGTABLE 
#DEFAULT 0.034 
#CUTCLASS V3 V3_0p480 V3_0p864 
#V3 0 0 0 0 0 0 
#V3_0p480 0 0 0 0 0 0 
#V3_0p864 0 0 0 0 0 0 
#; 
#" ; 
SPACING 0.034 ;

# ENCLOSURE CUTCLASS V3 END 0.005 SIDE 0 ; 
# covered below? 
# ENCLOSURE CUTCLASS V3 END 0.005 SIDE 0 ; 

# SWK
#PROPERTY LEF58_ENCLOSURE " 
#ENCLOSURE CUTCLASS V3 BELOW EOL 0 0.005 0 ; 
#ENCLOSURE CUTCLASS V3 ABOVE EOL 0 0.011 0 ; 
#ENCLOSURE CUTCLASS V3_0p480 END 0 SIDE 0 ; 
#ENCLOSURE CUTCLASS V3_0p864 END 0 SIDE 0 ; 
#" ; 

END V3 

LAYER M4 
TYPE ROUTING ; 
DIRECTION HORIZONTAL ; 
PITCH 0.048 ; 
WIDTH 0.024 ; 
SPACING 0.024 ; 

OFFSET 0.003 ; 

AREA 0.002 ; 

# SWK
# PROPERTY LEF58_SPACING " 
# SPACING 0.024 ENDOFLINE 0.025 WITHIN 0.04 ENDTOEND 0.04 ; " ; 
SPACING 0.04 ENDOFLINE 0.025 WITHIN 0.04 ;

PROPERTY LEF58_WIDTHTABLE 
" WIDTHTABLE 0.024 0.12 0.216 0.312 0.408 ; " ; 

PROPERTY LEF58_CORNERSPACING " 
CORNERSPACING CONVEXCORNER CORNERONLY 0.048 
WIDTH 0 SPACING 0.04 ; 
" ; 

PROPERTY LEF58_EOLKEEPOUT " 
EOLKEEPOUT 0.025 EXTENSION 0.048 0.02425 0.048 CORNERONLY ; 
" ; 

# spacing table is required for the rule that has wide metal requires a 72nm (288 scaled) 
# spacing between wide and minimum metals 

SPACINGTABLE 
PARALLELRUNLENGTH 0 
WIDTH 0 0.024 
WIDTH 0.025 0.072 ; 

PROPERTY LEF58_RIGHTWAYONGRIDONLY " 
RIGHTWAYONGRIDONLY ; 
" ; 

PROPERTY LEF58_RECTONLY " 
RECTONLY ; 
" ; 

END M4 

LAYER V4 
TYPE CUT ; 

# spacing is 1 * 8.5 = 34 
# SPACING 0.034 ; 
# WIDTH 0.018 ; 
# ENCLOSURE 0.011 0 ; 

# SWK
PROPERTY LEF58_CUTCLASS " 
CUTCLASS Vx WIDTH 0.024 LENGTH 0.024 ; 
CUTCLASS Vx_0p480 WIDTH 0.024 LENGTH 0.12 CUTS 1 ; 
CUTCLASS Vx_0p864 WIDTH 0.024 LENGTH 0.216 CUTS 2 ; 
CUTCLASS Vx_1p248 WIDTH 0.024 LENGTH 0.312 CUTS 3 ; 
CUTCLASS Vx_1p632 WIDTH 0.024 LENGTH 0.408 CUTS 4 ; 
" ; 
WIDTH 0.024 ;

#PROPERTY LEF58_SPACINGTABLE " 
#SPACINGTABLE 
#DEFAULT 0.034 
#CUTCLASS Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632 
#Vx 0 0 0 0 0 0 0 0 0 0 
#Vx_0p480 0 0 0 0 0 0 0 0 0 0 
#Vx_0p864 0 0 0 0 0 0 0 0 0 0 
#Vx_1p248 0 0 0 0 0 0 0 0 0 0 
#Vx_1p632 0 0 0 0 0 0 0 0 0 0 
#; 
#" ; 
SPACING 0.034 ;

# SWK
#PROPERTY LEF58_ENCLOSURE " 
#ENCLOSURE CUTCLASS Vx 0.011 0 ; 
#ENCLOSURE CUTCLASS Vx EOL 0 0.011 0.011 ; 
#ENCLOSURE CUTCLASS Vx_0p480 END 0 SIDE 0 ; 
#ENCLOSURE CUTCLASS Vx_0p864 END 0 SIDE 0 ; 
#ENCLOSURE CUTCLASS Vx_1p248 END 0 SIDE 0 ; 
#ENCLOSURE CUTCLASS Vx_1p632 END 0 SIDE 0 ; 
#" ; 

END V4 

LAYER M5 
TYPE ROUTING ; 
DIRECTION VERTICAL ; 
PITCH 0.048 ; 
WIDTH 0.024 ; 
SPACING 0.024 ; 
OFFSET 0 ; 

AREA 0.002 ; 

# SWK
# PROPERTY LEF58_SPACING " 
# SPACING 0.024 ENDOFLINE 0.025 WITHIN 0.04 ENDTOEND 0.04 ; " ; 
SPACING 0.04 ENDOFLINE 0.025 WITHIN 0.04 ;

MINIMUMDENSITY 15 ; 
MAXIMUMDENSITY 90 ; 
DENSITYCHECKWINDOW 20 20 ; 
DENSITYCHECKSTEP 10 ; 

PROPERTY LEF58_WIDTHTABLE 
" WIDTHTABLE 0.024 0.12 0.216 0.312 0.408 0.504 0.6 0.696 0.792 0.888 0.984 ; " ; 

PROPERTY LEF58_CORNERSPACING " 
CORNERSPACING CONVEXCORNER CORNERONLY 0.048 
WIDTH 0 SPACING 0.04 ; 
" ; 

PROPERTY LEF58_EOLKEEPOUT " 
EOLKEEPOUT 0.025 EXTENSION 0.048 0.02425 0.048 
CORNERONLY ; 
" ; 

SPACINGTABLE 
PARALLELRUNLENGTH 0 
WIDTH 0 0.024 
WIDTH 0.025 0.072 ; 

PROPERTY LEF58_RIGHTWAYONGRIDONLY " 
RIGHTWAYONGRIDONLY ; 
" ; 

PROPERTY LEF58_RECTONLY " 
RECTONLY ; 
" ; 

END M5 

LAYER V5 
TYPE CUT ; 

# SWK
PROPERTY LEF58_CUTCLASS " 
CUTCLASS Vx WIDTH 0.024 LENGTH 0.032 ; 
CUTCLASS Vx_0p480 WIDTH 0.024 LENGTH 0.16 CUTS 1 ; 
CUTCLASS Vx_0p864 WIDTH 0.024 LENGTH 0.288 CUTS 2 ; 
CUTCLASS Vx_1p248 WIDTH 0.024 LENGTH 0.416 CUTS 3 ; 
CUTCLASS Vx_1p632 WIDTH 0.024 LENGTH 0.544 CUTS 4 ; 
" ; 
WIDTH 0.024 ;

#PROPERTY LEF58_SPACINGTABLE " 
#SPACINGTABLE 
#DEFAULT 0.034 
#CUTCLASS Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632 
#Vx 0 0 0 0 0 0 0 0 0 0 
#Vx_0p480 0 0 0 0 0 0 0 0 0 0 
#Vx_0p864 0 0 0 0 0 0 0 0 0 0 
#Vx_1p248 0 0 0 0 0 0 0 0 0 0 
#Vx_1p632 0 0 0 0 0 0 0 0 0 0 
#; 
#" ; 
SPACING 0.034 ;

# end refers to the end of the VIA! Thus, since it is rectangular the proper 
# enclosure is on the side not the end... 
# ENCLOSURE CUTCLASS Vx END 0 SIDE 0.011 ; But--this refers to top and bottom 
# actually passing the rule is done by having the correct vias below. 

# SWK
#PROPERTY LEF58_ENCLOSURE " 
#ENCLOSURE CUTCLASS Vx EOL 0 0.011 0.011 ; 
#ENCLOSURE CUTCLASS Vx_0p480 END 0 SIDE 0 ; 
#ENCLOSURE CUTCLASS Vx_0p864 END 0 SIDE 0 ; 
#ENCLOSURE CUTCLASS Vx_1p248 END 0 SIDE 0 ; 
#ENCLOSURE CUTCLASS Vx_1p632 END 0 SIDE 0 ; 
#" ; 

# PROPERTY LEF58_ENCLOSURE " 
# ENCLOSURE CUTCLASS Vx EOL 0 0.011 0 ; 
# " ; 

END V5 

LAYER M6 
TYPE ROUTING ; 
DIRECTION HORIZONTAL ; 
PITCH 0.064 ; 
WIDTH 0.032 ; 
SPACING 0.032 ; 

AREA 0.0021875 ; # Areas still need tweaking 

# SWK
# PROPERTY LEF58_SPACING 
# " SPACING 0.032 ENDOFLINE 0.0375 WITHIN 0.04 ENDTOEND 0.04 ; " ; 
SPACING 0.04 ENDOFLINE 0.0375 WITHIN 0.04 ;

PROPERTY LEF58_WIDTHTABLE 
" WIDTHTABLE 0.032 0.16 0.288 0.416 0.544 ; " ; 

PROPERTY LEF58_CORNERSPACING " 
CORNERSPACING CONVEXCORNER CORNERONLY 0.048 
WIDTH 0 SPACING 0.04 ; 
" ; 

PROPERTY LEF58_EOLKEEPOUT " 
EOLKEEPOUT 0.05 EXTENSION 0.048 0.03225 0.048 CORNERONLY ; 
" ; 

SPACINGTABLE 
PARALLELRUNLENGTH 0 
WIDTH 0 0.024 
WIDTH 0.025 0.072 ; 

PROPERTY LEF58_RIGHTWAYONGRIDONLY " 
RIGHTWAYONGRIDONLY ; 
" ; 

PROPERTY LEF58_RECTONLY " 
RECTONLY ; 
" ; 

END M6 

LAYER V6 
TYPE CUT ; 

# SWK
PROPERTY LEF58_CUTCLASS " 
CUTCLASS Vx WIDTH 0.032 LENGTH 0.032 ; 
CUTCLASS Vx_0p640 WIDTH 0.032 LENGTH 0.16 CUTS 1 ; 
CUTCLASS Vx_1p152 WIDTH 0.032 LENGTH 0.288 CUTS 2 ; 
CUTCLASS Vx_1p664 WIDTH 0.032 LENGTH 0.416 CUTS 3 ; 
CUTCLASS Vx_2p176 WIDTH 0.032 LENGTH 0.544 CUTS 4 ; 
" ; 
WIDTH 0.032 ;

#PROPERTY LEF58_SPACINGTABLE " 
#SPACINGTABLE 
#DEFAULT 0.034 
#CUTCLASS Vx Vx_0p640 Vx_1p152 Vx_1p664 Vx_2p176 
#Vx 0 0 0 0 0 0 0 0 0 0 
#Vx_0p640 0 0 0 0 0 0 0 0 0 0 
#Vx_1p152 0 0 0 0 0 0 0 0 0 0 
#Vx_1p664 0 0 0 0 0 0 0 0 0 0 
#Vx_2p176 0 0 0 0 0 0 0 0 0 0 
#; 
#" ; 
SPACING 0.034 ;

# SWK
#PROPERTY LEF58_ENCLOSURE " 
#ENCLOSURE CUTCLASS Vx 0.011 0 ; 
#ENCLOSURE CUTCLASS Vx EOL 0 0.011 0.011 ; 
#ENCLOSURE CUTCLASS Vx_0p640 END 0 SIDE 0 ; 
#ENCLOSURE CUTCLASS Vx_1p152 END 0 SIDE 0 ; 
#ENCLOSURE CUTCLASS Vx_1p664 END 0 SIDE 0 ; 
#ENCLOSURE CUTCLASS Vx_2p176 END 0 SIDE 0 ; 
#" ; 

END V6 

LAYER M7 
TYPE ROUTING ; 
DIRECTION VERTICAL ; 
PITCH 0.064 ; 
WIDTH 0.032 ; 
SPACING 0.032 ; 

AREA 0.0021875 ; # Areas still need tweaking 

# SWK
# PROPERTY LEF58_SPACING 
# " SPACING 0.03 ENDOFLINE 0.0375 WITHIN 0.04 ENDTOEND 0.04 ; " ; 
SPACING 0.04 ENDOFLINE 0.0375 WITHIN 0.04 ;

PROPERTY LEF58_WIDTHTABLE 
" WIDTHTABLE 0.032 0.16 0.288 0.416 0.544 ; " ; 
TYPE ROUTING ; 
DIRECTION VERTICAL ; 

PROPERTY LEF58_CORNERSPACING " 
CORNERSPACING CONVEXCORNER CORNERONLY 0.075 
WIDTH 0 SPACING 0.04 ; 
" ; 

PROPERTY LEF58_EOLKEEPOUT " 
EOLKEEPOUT 0.05 EXTENSION 0.048 0.03225 0.048 
CORNERONLY ; 
" ; 

SPACINGTABLE 
PARALLELRUNLENGTH 0 
WIDTH 0 0.024 
WIDTH 0.025 0.072 ; 

PROPERTY LEF58_RIGHTWAYONGRIDONLY " 
RIGHTWAYONGRIDONLY ; 
" ; 

PROPERTY LEF58_RECTONLY " 
RECTONLY ; 
" ; 

END M7 

LAYER V7 
TYPE CUT ; 
SPACING 0.046 ; 
WIDTH 0.032 ; 
END V7 

LAYER M8 
TYPE ROUTING ; 
DIRECTION HORIZONTAL ; 
PITCH 0.08 0.08 ; 
WIDTH 0.04 ; 
AREA 1.88 ; 

SPACINGTABLE 
PARALLELRUNLENGTH 0 0.39975 1.19975 1.79975 
WIDTH 0 0.04 0.04 0.04 0.04 
WIDTH 0.05975 0.04 0.04 0.04 0.04 
WIDTH 0.07975 0.04 0.04 0.04 0.04 
WIDTH 0.11975 0.04 0.04 0.04 0.04 
WIDTH 0.49975 0.04 0.04 0.04 0.5 
WIDTH 0.99975 0.04 0.04 0.04 1 ; 

MINIMUMCUT 0.5 WIDTH 1.805 WITHIN 1.705 FROMBELOW ; 
MINIMUMCUT 0.5 WIDTH 1.805 WITHIN 1.705 FROMABOVE ; 
MAXWIDTH 2 ; 
MINSTEP 0.04 STEP ; 
END M8 

LAYER V8 
TYPE CUT ; 
SPACING 0.057 ; 
WIDTH 0.04 ; 
END V8 


LAYER M9 
TYPE ROUTING ; 
DIRECTION VERTICAL ; 
PITCH 0.08 0.08 ; 
WIDTH 0.04 ; 
AREA 1.88 ; 

SPACINGTABLE 
PARALLELRUNLENGTH 0 0.39975 1.19975 1.79975 
WIDTH 0 0.04 0.04 0.04 0.04 
WIDTH 0.05975 0.04 0.04 0.04 0.04 
WIDTH 0.07975 0.04 0.04 0.04 0.04 
WIDTH 0.11975 0.04 0.04 0.04 0.04 
WIDTH 0.49975 0.04 0.04 0.04 0.5 
WIDTH 0.99975 0.04 0.04 0.04 1 ; 

MINIMUMCUT 0.5 WIDTH 1.805 WITHIN 1.705 FROMABOVE ; 
MINSTEP 0.04 STEP ; 
END M9 

LAYER V9 
TYPE CUT ; 
SPACING 0.057 ; 
WIDTH 0.04 ; 
END V9 

LAYER Pad 
TYPE ROUTING ; 
DIRECTION HORIZONTAL ; 
PITCH 0.08 0.08 ; 
WIDTH 0.04 ; 
SPACINGTABLE 
PARALLELRUNLENGTH 0 11.99975 
WIDTH 0 2 2 
WIDTH 11.99975 2 3 ; 
MINIMUMCUT 0.25 WIDTH 0.04 WITHIN 1.705 FROMBELOW ; 
MINIMUMCUT 0.25 WIDTH 0.36 WITHIN 1.705 FROMBELOW ; 
MINIMUMCUT 0.5 WIDTH 1.805 WITHIN 1.705 FROMBELOW ; 
MINIMUMDENSITY 20 ; 
MAXIMUMDENSITY 80 ; 
DENSITYCHECKWINDOW 100 100 ; 
DENSITYCHECKSTEP 50 ; 
END Pad 

# vias 

VIA VIA9Pad Default 
LAYER M9 ; 
RECT -0.05 -0.05 0.05 0.05 ; 
LAYER Pad ; 
RECT -0.05 -0.05 0.05 0.05 ; 
LAYER V9 ; 
RECT -0.05 -0.05 0.05 0.05 ; 
END VIA9Pad 

VIA VIA89 Default 
LAYER M8 ; 
RECT -0.02 -0.02 0.02 0.02 ; 
LAYER M9 ; 
RECT -0.02 -0.02 0.02 0.02 ; 
LAYER V8 ; 
RECT -0.02 -0.02 0.02 0.02 ; 
END VIA89 

VIA VIA78 Default 
LAYER M7 ; 
RECT -0.016 -0.027 0.016 0.027 ; 
LAYER M8 ; 
RECT -0.027 -0.016 0.027 0.016 ; 
LAYER V7 ; 
RECT -0.016 -0.016 0.016 0.016 ; 
END VIA78 

VIA VIA67 Default 
LAYER M6 ; 
RECT -0.027 -0.016 0.027 0.016 ; 
LAYER M7 ; 
RECT -0.016 -0.027 0.016 0.027 ; 
LAYER V6 ; 
RECT -0.016 -0.016 0.016 0.016 ; 
END VIA67 

VIA VIA56 Default 
LAYER M5 ; 
RECT -0.012 -0.027 0.012 0.027 ; 
LAYER M6 ; 
RECT -0.023 -0.016 0.023 0.016 ; 
LAYER V5 ; 
RECT -0.012 -0.016 0.012 0.016 ; 
END VIA56 

VIA VIA45 Default 
LAYER M4 ; 
RECT -0.023 -0.012 0.023 0.012 ; 
LAYER M5 ; 
RECT -0.012 -0.023 0.012 0.023 ; 
LAYER V4 ; 
RECT -0.012 -0.012 0.012 0.012 ; 
END VIA45 

VIA VIA34 Default 
LAYER M3 ; 
RECT -0.009 -0.017 0.009 0.017 ; 
LAYER M4 ; 
RECT -0.02 -0.012 0.02 0.012 ; 
LAYER V3 ; 
RECT -0.009 -0.012 0.009 0.012 ; 
END VIA34 

VIA VIA23 Default 
LAYER M2 ; 
RECT -0.014 -0.009 0.014 0.009 ; 
LAYER M3 ; 
RECT -0.009 -0.014 0.009 0.014 ; 
LAYER V2 ; 
RECT -0.009 -0.009 0.009 0.009 ; 
END VIA23 

VIA VIA12 Default 
LAYER M1 ; 
RECT -0.009 -0.011 0.009 0.011 ; 
LAYER M2 ; 
RECT -0.014 -0.009 0.014 0.009 ; 
LAYER V1 ; 
RECT -0.009 -0.009 0.009 0.009 ; 
END VIA12 

################################# 
### VIARULE GENERATE DEFAULTS ### 
################################# 

VIARULE Pad_M9 GENERATE DEFAULT 
LAYER M9 ; 
ENCLOSURE 0 0 ; 
LAYER Pad ; 
ENCLOSURE 0.011 0 ; 
LAYER V9 ; 
RECT -0.016 -0.016 0.016 0.016 ; 
SPACING 0.078 BY 0.078 ; 
END Pad_M9 

VIARULE M9_M8 GENERATE DEFAULT 
LAYER M8 ; 
ENCLOSURE 0 0 ; 
LAYER M9 ; 
ENCLOSURE 0 0.02 ; 
LAYER V8 ; 
RECT -0.02 -0.02 0.02 0.02 ; 
SPACING 0.097 BY 0.097 ; 
END M9_M8 

VIARULE M8_M7 GENERATE DEFAULT 
LAYER M7 ; 
ENCLOSURE 0 0 ; 
LAYER M8 ; 
ENCLOSURE 0.011 0 ; 
LAYER V7 ; 
RECT -0.016 -0.016 0.016 0.016 ; 
SPACING 0.078 BY 0.078 ; 
END M8_M7 

VIARULE M7_M6 GENERATE DEFAULT 
LAYER M6 ; 
ENCLOSURE 0.011 0 ; 
LAYER M7 ; 
ENCLOSURE 0 0.011 ; 
LAYER V6 ; 
RECT -0.016 -0.016 0.016 0.016 ; 
SPACING 0.078 BY 0.078 ; 
END M7_M6 

VIARULE M6_M5 GENERATE DEFAULT 
LAYER M5 ; 
ENCLOSURE 0.011 0 ; 
WIDTH 0.024 TO 0.024 ; 
LAYER M6 ; 
ENCLOSURE 0.011 0 ; 
WIDTH 0.032 TO 0.032 ; 
LAYER V5 ; 
RECT -0.012 -0.016 0.012 0.016 ; 
SPACING 0.058 BY 0.308 ; # purposely crazy to avoid dual cut on routing 
END M6_M5 


# to make the wide vias for power stripes (still SAV) 

VIARULE M3_M2widePWR0p936 GENERATE 
LAYER M2 ; 
ENCLOSURE 0 0 ; 
LAYER M3 ; 
ENCLOSURE 0 0 ; 
WIDTH 0.234 TO 0.234 ; 
LAYER V2 ; 
RECT -0.117 -0.009 0.117 0.009 ; 
SPACING 0.277 BY 0.036 ; 
END M3_M2widePWR0p936 

# to make the wide vias for powers (still SAV) 

VIARULE M4_M3widePWR0p864 GENERATE 
LAYER M3 ; 
ENCLOSURE 0 0 ; 
WIDTH 0.2335 TO 0.2345 ; 
LAYER M4 ; 
ENCLOSURE 0 0 ; 
WIDTH 0.2155 TO 0.2165 ; 
LAYER V3 ; 
RECT -0.009 -0.108 0.009 0.108 ; 
SPACING 0.036 BY 0.277 ; 
END M4_M3widePWR0p864 

# to make the wide vias for powers (still SAV) 

VIARULE M5_M4widePWR0p864 GENERATE 
LAYER M4 ; 
ENCLOSURE 0 0 ; 
LAYER M5 ; 
ENCLOSURE 0 0 ; 
WIDTH 0.216 TO 0.216 ; 
LAYER V4 ; 
RECT -0.108 -0.012 0.108 0.012 ; 
SPACING 0.532 BY 0.096 ; 
END M5_M4widePWR0p864 

# to make the wide vias for powers (still SAV) 

VIARULE M6_M5widePWR1p152 GENERATE 
LAYER M5 ; 
ENCLOSURE 0 0 ; 
LAYER M6 ; 
ENCLOSURE 0 0 ; 
WIDTH 0.288 TO 0.288 ; 
LAYER V5 ; 
RECT -0.012 -0.144 0.012 0.144 ; 
SPACING 0.096 BY 0.382 ; 
END M6_M5widePWR1p152 

# to make the wide vias for powers (still SAV) 

VIARULE M7_M6widePWR1p152 GENERATE 
LAYER M6 ; 
ENCLOSURE 0 0 ; 
LAYER M7 ; 
ENCLOSURE 0 0 ; 
WIDTH 0.288 TO 0.288 ; 
LAYER V6 ; 
RECT -0.144 -0.016 0.144 0.016 ; 
SPACING 0.532 BY 0.096 ; 
END M7_M6widePWR1p152 

VIARULE M2_M1 GENERATE DEFAULT 
LAYER M1 ; 
ENCLOSURE 0 0 ; 
LAYER M2 ; 
ENCLOSURE 0.002 0 ; 
LAYER V1 ; 
RECT -0.009 -0.009 0.009 0.009 ; 
SPACING 0.036 BY 0.036 ; 
END M2_M1 

END LIBRARY 
