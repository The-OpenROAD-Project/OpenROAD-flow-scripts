../../nangate45/lef/fakeram45_64x96.lef