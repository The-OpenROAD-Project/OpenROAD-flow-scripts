VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_1024x8
  FOREIGN fakeram130_1024x8 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 532.190 BY 308.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 16.600 0.800 17.400 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.400 0.800 24.200 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 30.200 0.800 31.000 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.000 0.800 37.800 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.800 0.800 44.600 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 50.600 0.800 51.400 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 57.400 0.800 58.200 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 64.200 0.800 65.000 ;
    END
  END w_mask_in[7]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 69.300 0.800 70.100 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 76.100 0.800 76.900 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 82.900 0.800 83.700 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 89.700 0.800 90.500 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 96.500 0.800 97.300 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 103.300 0.800 104.100 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 110.100 0.800 110.900 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 116.900 0.800 117.700 ;
    END
  END rd_out[7]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 122.000 0.800 122.800 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 128.800 0.800 129.600 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 135.600 0.800 136.400 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 142.400 0.800 143.200 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 149.200 0.800 150.000 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.000 0.800 156.800 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 162.800 0.800 163.600 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 169.600 0.800 170.400 ;
    END
  END wd_in[7]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 174.700 0.800 175.500 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 181.500 0.800 182.300 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 188.300 0.800 189.100 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 195.100 0.800 195.900 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 201.900 0.800 202.700 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 208.700 0.800 209.500 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 215.500 0.800 216.300 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 222.300 0.800 223.100 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 229.100 0.800 229.900 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 235.900 0.800 236.700 ;
    END
  END addr_in[9]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 241.000 0.800 241.800 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 247.800 0.800 248.600 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 254.600 0.800 255.400 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 15.400 17.000 18.600 291.000 ;
      RECT 42.600 17.000 45.800 291.000 ;
      RECT 69.800 17.000 73.000 291.000 ;
      RECT 97.000 17.000 100.200 291.000 ;
      RECT 124.200 17.000 127.400 291.000 ;
      RECT 151.400 17.000 154.600 291.000 ;
      RECT 178.600 17.000 181.800 291.000 ;
      RECT 205.800 17.000 209.000 291.000 ;
      RECT 233.000 17.000 236.200 291.000 ;
      RECT 260.200 17.000 263.400 291.000 ;
      RECT 287.400 17.000 290.600 291.000 ;
      RECT 314.600 17.000 317.800 291.000 ;
      RECT 341.800 17.000 345.000 291.000 ;
      RECT 369.000 17.000 372.200 291.000 ;
      RECT 396.200 17.000 399.400 291.000 ;
      RECT 423.400 17.000 426.600 291.000 ;
      RECT 450.600 17.000 453.800 291.000 ;
      RECT 477.800 17.000 481.000 291.000 ;
      RECT 505.000 17.000 508.200 291.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 29.000 17.000 32.200 291.000 ;
      RECT 56.200 17.000 59.400 291.000 ;
      RECT 83.400 17.000 86.600 291.000 ;
      RECT 110.600 17.000 113.800 291.000 ;
      RECT 137.800 17.000 141.000 291.000 ;
      RECT 165.000 17.000 168.200 291.000 ;
      RECT 192.200 17.000 195.400 291.000 ;
      RECT 219.400 17.000 222.600 291.000 ;
      RECT 246.600 17.000 249.800 291.000 ;
      RECT 273.800 17.000 277.000 291.000 ;
      RECT 301.000 17.000 304.200 291.000 ;
      RECT 328.200 17.000 331.400 291.000 ;
      RECT 355.400 17.000 358.600 291.000 ;
      RECT 382.600 17.000 385.800 291.000 ;
      RECT 409.800 17.000 413.000 291.000 ;
      RECT 437.000 17.000 440.200 291.000 ;
      RECT 464.200 17.000 467.400 291.000 ;
      RECT 491.400 17.000 494.600 291.000 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 532.190 308.000 ;
    LAYER met2 ;
    RECT 0 0 532.190 308.000 ;
    LAYER met3 ;
    RECT 0.800 0 532.190 308.000 ;
    RECT 0 0.000 0.800 16.600 ;
    RECT 0 17.400 0.800 23.400 ;
    RECT 0 24.200 0.800 30.200 ;
    RECT 0 31.000 0.800 37.000 ;
    RECT 0 37.800 0.800 43.800 ;
    RECT 0 44.600 0.800 50.600 ;
    RECT 0 51.400 0.800 57.400 ;
    RECT 0 58.200 0.800 64.200 ;
    RECT 0 65.000 0.800 69.300 ;
    RECT 0 70.100 0.800 76.100 ;
    RECT 0 76.900 0.800 82.900 ;
    RECT 0 83.700 0.800 89.700 ;
    RECT 0 90.500 0.800 96.500 ;
    RECT 0 97.300 0.800 103.300 ;
    RECT 0 104.100 0.800 110.100 ;
    RECT 0 110.900 0.800 116.900 ;
    RECT 0 117.700 0.800 122.000 ;
    RECT 0 122.800 0.800 128.800 ;
    RECT 0 129.600 0.800 135.600 ;
    RECT 0 136.400 0.800 142.400 ;
    RECT 0 143.200 0.800 149.200 ;
    RECT 0 150.000 0.800 156.000 ;
    RECT 0 156.800 0.800 162.800 ;
    RECT 0 163.600 0.800 169.600 ;
    RECT 0 170.400 0.800 174.700 ;
    RECT 0 175.500 0.800 181.500 ;
    RECT 0 182.300 0.800 188.300 ;
    RECT 0 189.100 0.800 195.100 ;
    RECT 0 195.900 0.800 201.900 ;
    RECT 0 202.700 0.800 208.700 ;
    RECT 0 209.500 0.800 215.500 ;
    RECT 0 216.300 0.800 222.300 ;
    RECT 0 223.100 0.800 229.100 ;
    RECT 0 229.900 0.800 235.900 ;
    RECT 0 236.700 0.800 241.000 ;
    RECT 0 241.800 0.800 247.800 ;
    RECT 0 248.600 0.800 254.600 ;
    RECT 0 255.400 0.800 308.000 ;
    LAYER met4 ;
    RECT 0 0 532.190 17.000 ;
    RECT 0 291.000 532.190 308.000 ;
    RECT 0.000 17.000 15.400 291.000 ;
    RECT 18.600 17.000 29.000 291.000 ;
    RECT 32.200 17.000 42.600 291.000 ;
    RECT 45.800 17.000 56.200 291.000 ;
    RECT 59.400 17.000 69.800 291.000 ;
    RECT 73.000 17.000 83.400 291.000 ;
    RECT 86.600 17.000 97.000 291.000 ;
    RECT 100.200 17.000 110.600 291.000 ;
    RECT 113.800 17.000 124.200 291.000 ;
    RECT 127.400 17.000 137.800 291.000 ;
    RECT 141.000 17.000 151.400 291.000 ;
    RECT 154.600 17.000 165.000 291.000 ;
    RECT 168.200 17.000 178.600 291.000 ;
    RECT 181.800 17.000 192.200 291.000 ;
    RECT 195.400 17.000 205.800 291.000 ;
    RECT 209.000 17.000 219.400 291.000 ;
    RECT 222.600 17.000 233.000 291.000 ;
    RECT 236.200 17.000 246.600 291.000 ;
    RECT 249.800 17.000 260.200 291.000 ;
    RECT 263.400 17.000 273.800 291.000 ;
    RECT 277.000 17.000 287.400 291.000 ;
    RECT 290.600 17.000 301.000 291.000 ;
    RECT 304.200 17.000 314.600 291.000 ;
    RECT 317.800 17.000 328.200 291.000 ;
    RECT 331.400 17.000 341.800 291.000 ;
    RECT 345.000 17.000 355.400 291.000 ;
    RECT 358.600 17.000 369.000 291.000 ;
    RECT 372.200 17.000 382.600 291.000 ;
    RECT 385.800 17.000 396.200 291.000 ;
    RECT 399.400 17.000 409.800 291.000 ;
    RECT 413.000 17.000 423.400 291.000 ;
    RECT 426.600 17.000 437.000 291.000 ;
    RECT 440.200 17.000 450.600 291.000 ;
    RECT 453.800 17.000 464.200 291.000 ;
    RECT 467.400 17.000 477.800 291.000 ;
    RECT 481.000 17.000 491.400 291.000 ;
    RECT 494.600 17.000 505.000 291.000 ;
    RECT 508.200 17.000 532.190 291.000 ;
    LAYER OVERLAP ;
    RECT 0 0 532.190 308.000 ;
  END
END fakeram130_1024x8

END LIBRARY
