VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addf_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 18.48 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.272 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.615 1.77 3.47 1.77 3.47 2.15 1.615 2.15  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.272 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.64 1.795 17.07 1.795 17.07 2.15 14.64 2.15  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.694 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.89 1.62 8.415 1.62 12.34 1.62 12.34 1.2 13.21 1.2 13.54 1.2 13.54 0.55 13.91 0.55 13.91 1.85 13.21 1.85 8.415 1.85 3.89 1.85  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8932 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.45 0.79 17.83 0.79 17.83 3.37 17.45 3.37  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.847 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 0.61 0.575 0.61 0.575 3.37 0.14 3.37  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3.04 1.595 3.04 1.595 3.62 4.71 3.62 6.79 3.62 6.79 3.005 7.13 3.005 7.13 3.62 8.37 3.62 9.105 3.62 9.105 2.705 9.335 2.705 9.335 3.62 11.31 3.62 11.31 3.005 11.65 3.005 11.65 3.62 13.43 3.62 16.445 3.62 16.445 2.48 16.675 2.48 16.675 3.62 17.2 3.62 18.48 3.62 18.48 4.22 17.2 4.22 13.43 4.22 8.37 4.22 4.71 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 18.48 -0.3 18.48 0.3 16.675 0.3 16.675 0.765 16.445 0.765 16.445 0.3 11.65 0.3 11.65 0.915 11.31 0.915 11.31 0.3 9.59 0.3 9.59 1.09 9.25 1.09 9.25 0.3 7.13 0.3 7.13 0.915 6.79 0.915 6.79 0.3 1.595 0.3 1.595 0.87 1.365 0.87 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.155 2.56 4.71 2.56 4.71 2.79 0.925 2.79 0.925 1.16 4.385 1.16 4.385 0.81 4.615 0.81 4.615 1.39 1.155 1.39  ;
        POLYGON 5.55 2.545 8.37 2.545 8.37 2.845 8.03 2.845 8.03 2.775 5.89 2.775 5.89 2.845 5.55 2.845  ;
        POLYGON 5.505 0.81 5.735 0.81 5.735 1.145 8.185 1.145 8.185 0.81 8.415 0.81 8.415 1.375 5.505 1.375  ;
        POLYGON 10.025 0.77 10.255 0.77 10.255 1.145 11.88 1.145 11.88 0.68 13.21 0.68 13.21 0.915 12.11 0.915 12.11 1.375 10.025 1.375  ;
        POLYGON 10.07 2.545 13.43 2.545 13.43 2.775 10.07 2.775  ;
        POLYGON 5.01 2.08 14.17 2.08 14.17 0.75 14.495 0.75 14.495 1.335 17.2 1.335 17.2 1.565 14.4 1.565 14.4 2.765 14.165 2.765 14.165 2.315 5.01 2.315  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addf_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.372 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.605 1.76 4.13 1.76 4.13 2.16 2.605 2.16  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.372 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.58 1.76 17.335 1.76 17.335 2.16 16.7 2.16 16.7 3.37 16.34 3.37 16.34 2.16 15.58 2.16  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.754 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.49 1.605 9.695 1.605 14.215 1.605 14.525 1.605 14.525 1.345 14.755 1.345 14.755 1.835 14.215 1.835 9.695 1.835 5.66 1.835 5.66 2.16 4.49 2.16  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0452 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.37 0.55 18.96 0.55 18.96 3.37 18.37 3.37  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.22 0.55 1.68 0.55 1.68 3.37 1.22 3.37  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.385 3.62 0.385 2.46 0.615 2.46 0.615 3.62 2.37 3.62 2.37 3.285 2.71 3.285 2.71 3.62 5.83 3.62 7.95 3.62 7.95 3.005 8.29 3.005 8.29 3.62 9.79 3.62 10.53 3.62 10.53 2.845 10.87 2.845 10.87 3.62 12.49 3.62 12.49 3.005 12.83 3.005 12.83 3.62 14.31 3.62 17.405 3.62 17.405 2.48 17.635 2.48 17.635 3.62 18.12 3.62 19.445 3.62 19.445 2.48 19.675 2.48 19.675 3.62 20.16 3.62 20.16 4.22 18.12 4.22 14.31 4.22 9.79 4.22 5.83 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 19.775 0.3 19.775 0.905 19.545 0.905 19.545 0.3 17.57 0.3 17.57 0.73 17.23 0.73 17.23 0.3 12.93 0.3 12.93 0.915 12.59 0.915 12.59 0.3 10.87 0.3 10.87 1.075 10.53 1.075 10.53 0.3 8.29 0.3 8.29 0.915 7.95 0.915 7.95 0.3 2.755 0.3 2.755 0.695 2.525 0.695 2.525 0.3 0.515 0.3 0.515 0.905 0.285 0.905 0.285 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.17 2.61 5.83 2.61 5.83 2.845 1.94 2.845 1.94 0.925 5.545 0.925 5.545 0.78 5.775 0.78 5.775 1.155 2.17 1.155  ;
        POLYGON 6.665 0.79 6.895 0.79 6.895 1.145 9.465 1.145 9.465 0.79 9.695 0.79 9.695 1.375 6.665 1.375  ;
        POLYGON 6.71 2.54 9.79 2.54 9.79 2.775 6.71 2.775  ;
        POLYGON 11.305 0.79 11.535 0.79 11.535 1.145 13.985 1.145 13.985 0.79 14.215 0.79 14.215 1.375 11.305 1.375  ;
        POLYGON 11.24 2.545 14.31 2.545 14.31 2.775 11.24 2.775  ;
        POLYGON 6.07 2.065 15.105 2.065 15.105 0.78 15.335 0.78 15.335 1.085 18.12 1.085 18.12 2.23 17.89 2.23 17.89 1.315 15.335 1.315 15.335 3.14 15.105 3.14 15.105 2.295 6.07 2.295  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addf_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 24.64 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.352 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.095 1.77 6.785 1.77 6.785 2.15 5.095 2.15  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.352 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.45 1.77 19.65 1.77 19.65 2.16 17.45 2.16  ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.734 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.33 1.625 11.86 1.625 12.325 1.625 12.325 0.65 12.755 0.65 12.755 1.625 16.615 1.625 17.11 1.625 17.11 1.855 16.615 1.855 11.86 1.855 7.33 1.855  ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.5972 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.79 1.92 22.785 1.92 23.03 1.92 23.03 1.135 20.805 1.135 20.805 0.53 21.035 0.53 21.035 0.905 23.03 0.905 23.03 0.53 23.41 0.53 23.41 3.37 23.03 3.37 23.03 2.24 22.785 2.24 21.26 2.24 21.26 3.37 20.79 3.37  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.4244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.675 1.92 3.915 1.92 3.915 3.37 3.46 3.37 3.46 2.24 1.675 2.24 1.675 3.37 1.215 3.37 1.215 0.53 1.675 0.53 1.675 0.905 3.685 0.905 3.685 0.53 3.915 0.53 3.915 1.135 1.675 1.135  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.325 3.62 0.325 2.65 0.555 2.65 0.555 3.62 2.565 3.62 2.565 2.65 2.795 2.65 2.795 3.62 4.805 3.62 4.805 3.16 5.035 3.16 5.035 3.62 8.11 3.62 10.23 3.62 10.23 3.005 10.57 3.005 10.57 3.62 11.93 3.62 12.765 3.62 12.765 2.67 12.995 2.67 12.995 3.62 14.99 3.62 14.99 3.005 15.33 3.005 15.33 3.62 16.57 3.62 19.585 3.62 19.585 3.16 19.815 3.16 19.815 3.62 21.925 3.62 21.925 2.56 22.155 2.56 22.155 3.62 22.785 3.62 24.165 3.62 24.165 2.56 24.395 2.56 24.395 3.62 24.64 3.62 24.64 4.22 22.785 4.22 16.57 4.22 11.93 4.22 8.11 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 24.64 -0.3 24.64 0.3 24.395 0.3 24.395 0.765 24.165 0.765 24.165 0.3 22.21 0.3 22.21 0.67 21.87 0.67 21.87 0.3 19.915 0.3 19.915 0.765 19.685 0.765 19.685 0.3 15.33 0.3 15.33 0.915 14.99 0.915 14.99 0.3 13.215 0.3 13.215 1.135 12.985 1.135 12.985 0.3 10.57 0.3 10.57 0.915 10.23 0.915 10.23 0.3 5.09 0.3 5.09 0.675 4.75 0.675 4.75 0.3 2.85 0.3 2.85 0.675 2.505 0.675 2.505 0.3 0.555 0.3 0.555 0.87 0.325 0.87 0.325 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 4.79 2.545 8.11 2.545 8.11 2.775 4.56 2.775 4.56 1.67 1.915 1.67 1.915 1.44 4.56 1.44 4.56 0.905 7.77 0.905 7.77 0.78 8.11 0.78 8.11 1.14 4.79 1.14  ;
        POLYGON 8.945 0.795 9.175 0.795 9.175 1.145 11.63 1.145 11.63 0.795 11.86 0.795 11.86 1.375 8.945 1.375  ;
        POLYGON 8.99 2.545 11.93 2.545 11.93 2.83 11.59 2.83 11.59 2.775 9.33 2.775 9.33 2.83 8.99 2.83  ;
        POLYGON 13.74 2.545 16.57 2.545 16.57 2.775 13.74 2.775  ;
        POLYGON 13.705 0.81 13.935 0.81 13.935 1.145 16.385 1.145 16.385 0.81 16.615 0.81 16.615 1.375 13.705 1.375  ;
        POLYGON 8.38 2.085 17.165 2.085 17.165 2.55 20.125 2.55 20.125 1.365 17.505 1.365 17.505 0.81 17.735 0.81 17.735 1.135 20.355 1.135 20.355 1.44 22.785 1.44 22.785 1.67 20.355 1.67 20.355 2.785 16.935 2.785 16.935 2.315 8.38 2.315  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addf_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addh_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addh_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.175 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.505 1.77 3.27 1.77 3.27 2.365 5.865 2.365 5.865 1.87 6.095 1.87 6.095 2.595 2.775 2.595 2.775 2.15 1.505 2.15  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.175 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.725 1.79 5.51 1.79 5.51 2.135 3.725 2.135  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8954 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 0.65 0.575 0.65 0.575 3.37 0.14 3.37  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8954 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.975 0.65 9.735 0.65 9.735 3.37 9.405 3.37 9.405 1.68 8.975 1.68  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3.23 1.595 3.23 1.595 3.62 3.59 3.62 3.59 3.285 3.93 3.285 3.93 3.62 4.33 3.62 4.33 3.285 4.67 3.285 4.67 3.62 8.205 3.62 8.205 3.075 8.435 3.075 8.435 3.62 9.055 3.62 10.08 3.62 10.08 4.22 9.055 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 8.49 0.3 8.49 1.035 8.15 1.035 8.15 0.3 1.65 0.3 1.65 0.64 1.31 0.64 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 4.23 0.53 7.25 0.53 7.25 1.035 6.91 1.035 6.91 0.76 4.57 0.76 4.57 1.035 4.23 1.035  ;
        POLYGON 1.155 2.77 2.37 2.77 2.37 3.1 3.11 3.1 3.11 2.825 6.415 2.825 6.415 1.74 7.91 1.74 7.91 1.97 6.645 1.97 6.645 3.055 3.34 3.055 3.34 3.33 2.14 3.33 2.14 3 0.925 3 0.925 0.87 3.475 0.87 3.475 0.81 3.85 0.81 3.85 1.1 1.155 1.1  ;
        POLYGON 7.01 3.01 7.12 3.01 7.12 2.375 8.14 2.375 8.14 1.495 5.57 1.495 5.57 0.99 5.91 0.99 5.91 1.265 8.37 1.265 8.37 1.91 9.055 1.91 9.055 2.25 8.37 2.25 8.37 2.61 7.35 2.61 7.35 3.24 7.01 3.24  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addh_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addh_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addh_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.073 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.715 1.74 3.78 1.74 3.78 2.35 7.38 2.35 7.38 2.205 7.77 2.205 7.77 2.71 3.435 2.71 3.435 2.15 2.715 2.15  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.073 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.01 1.21 4.39 1.21 4.39 1.72 5.62 1.72 5.62 2.12 4.01 2.12  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1771 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 0.55 1.615 0.55 1.615 3.37 1.21 3.37  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.9308 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.49 2.25 10.79 2.25 11.31 2.25 11.31 1.56 10.49 1.56 10.49 0.55 11.11 0.55 11.11 1.22 11.65 1.22 11.65 2.48 11.11 2.48 11.11 3.37 10.79 3.37 10.49 3.37  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.315 3.62 0.315 2.48 0.545 2.48 0.545 3.62 2.4 3.62 2.4 3.215 2.74 3.215 2.74 3.62 4.49 3.62 4.49 3.215 4.83 3.215 4.83 3.62 5.43 3.62 5.43 3.215 5.77 3.215 5.77 3.62 9.37 3.62 9.37 2.685 9.71 2.685 9.71 3.62 10.79 3.62 11.51 3.62 11.51 2.71 11.85 2.71 11.85 3.62 12.32 3.62 12.32 4.22 10.79 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 11.895 0.3 11.895 0.78 11.665 0.78 11.665 0.3 9.655 0.3 9.655 0.78 9.425 0.78 9.425 0.3 2.735 0.3 2.735 0.94 2.505 0.94 2.505 0.3 0.495 0.3 0.495 0.985 0.265 0.985 0.265 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 5.33 0.53 8.35 0.53 8.35 0.76 5.33 0.76  ;
        POLYGON 2.015 1.18 3.125 1.18 3.125 0.53 4.895 0.53 4.895 1.19 6.325 1.19 6.325 1.745 8.79 1.745 8.79 1.975 6.095 1.975 6.095 1.42 4.665 1.42 4.665 0.76 3.355 0.76 3.355 1.41 2.245 1.41 2.245 2.755 3.205 2.755 3.205 2.94 3.81 2.94 3.81 3.17 2.975 3.17 2.975 2.985 2.015 2.985  ;
        POLYGON 8.01 2.205 9.17 2.205 9.17 1.515 6.67 1.515 6.67 0.99 7.01 0.99 7.01 1.285 9.4 1.285 9.4 1.79 10.79 1.79 10.79 2.02 9.4 2.02 9.4 2.435 8.35 2.435 8.35 3.37 8.01 3.37  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addh_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__addh_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__addh_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.1 1.685 1.33 1.685 1.33 2.015 3.905 2.015 3.905 1.8 5.845 1.8 5.845 2.015 10.47 2.015 10.47 2.245 1.1 2.245  ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 1.2 3.965 1.2 3.965 1.305 6.585 1.305 6.585 1.555 7.62 1.555 7.62 1.785 6.355 1.785 6.355 1.57 3.47 1.57 3.47 1.775 1.64 1.775  ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2701 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.17 1.035 13.56 1.035 13.56 1.77 15.9 1.77 15.9 1.035 16.24 1.035 16.24 2.885 15.85 2.885 15.85 2.15 13.51 2.15 13.51 2.885 13.17 2.885  ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.0903 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.22 2.245 19.86 2.245 20.25 2.245 20.25 1.37 18.22 1.37 18.22 0.54 18.605 0.54 18.605 1.135 20.25 1.135 20.25 0.65 20.845 0.65 20.845 3.39 20.25 3.39 20.25 2.48 19.86 2.48 18.56 2.48 18.56 3.39 18.22 3.39  ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.145 0.475 3.145 0.475 3.62 2.335 3.62 2.335 3.105 2.565 3.105 2.565 3.62 4.425 3.62 4.425 3.105 4.655 3.105 4.655 3.62 8.3 3.62 8.3 3.445 8.64 3.445 8.64 3.62 12.045 3.62 12.045 3.285 12.385 3.285 12.385 3.62 14.51 3.62 14.51 3.285 14.85 3.285 14.85 3.62 17.125 3.62 17.125 2.73 17.355 2.73 17.355 3.62 19.395 3.62 19.395 2.73 19.625 2.73 19.625 3.62 19.86 3.62 21.605 3.62 21.605 2.73 21.835 2.73 21.835 3.62 22.4 3.62 22.4 4.22 19.86 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 21.965 0.3 21.965 0.935 21.735 0.935 21.735 0.3 19.78 0.3 19.78 0.735 19.44 0.735 19.44 0.3 17.455 0.3 17.455 0.935 17.225 0.935 17.225 0.3 14.9 0.3 14.9 0.635 14.56 0.635 14.56 0.3 12.44 0.3 12.44 1.12 12.09 1.12 12.09 0.3 4.71 0.3 4.71 1.075 4.37 1.075 4.37 0.3 0.475 0.3 0.475 0.69 0.245 0.69 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 5.72 0.63 11.1 0.63 11.1 1.075 10.76 1.075 10.76 0.86 8.64 0.86 8.64 0.915 8.3 0.915 8.3 0.86 6.06 0.86 6.06 1.075 5.72 1.075  ;
        POLYGON 0.87 2.525 10.7 2.525 10.7 1.815 12.88 1.815 12.88 2.045 10.93 2.045 10.93 2.755 3.69 2.755 3.69 3.39 3.35 3.39 3.35 2.815 1.6 2.815 1.6 3.39 1.255 3.39 1.255 2.815 0.64 2.815 0.64 1.09 1.025 1.09 1.025 0.54 2.67 0.54 2.67 0.77 1.255 0.77 1.255 1.32 0.87 1.32  ;
        POLYGON 5.72 2.985 11.385 2.985 11.385 2.825 12.89 2.825 12.89 3.115 13.825 3.115 13.825 2.75 15.545 2.75 15.545 3.115 16.47 3.115 16.47 0.76 15.565 0.76 15.565 1.235 14.03 1.235 14.03 0.76 12.92 0.76 12.92 1.585 9.64 1.585 9.64 1.38 7.885 1.38 7.885 1.325 6.84 1.325 6.84 1.09 8.115 1.09 8.115 1.145 9.64 1.145 9.64 1.09 9.98 1.09 9.98 1.35 12.69 1.35 12.69 0.53 14.26 0.53 14.26 1.005 15.335 1.005 15.335 0.53 16.7 0.53 16.7 1.74 19.86 1.74 19.86 1.97 16.7 1.97 16.7 3.345 15.315 3.345 15.315 2.98 14.055 2.98 14.055 3.345 12.66 3.345 12.66 3.055 11.615 3.055 11.615 3.215 5.72 3.215  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__addh_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.519 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.54 1.02 1.54 1.02 2.81 0.66 2.81  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.519 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 1.54 2.14 1.54 2.14 3.37 1.78 3.37  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8932 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 0.555 3.87 0.555 3.87 3.38 3.45 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.225 0.475 3.225 0.475 3.62 2.605 3.62 2.605 2.53 2.835 2.53 2.835 3.62 3.175 3.62 4.48 3.62 4.48 4.22 3.175 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 2.735 0.3 2.735 0.765 2.505 0.765 2.505 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.805 0.475 0.805 0.475 1.055 3.175 1.055 3.175 1.985 2.945 1.985 2.945 1.29 1.495 1.29 1.495 3.325 1.265 3.325 1.265 1.29 0.245 1.29  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and2_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.04 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.024 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.065 1.02 1.065 1.02 2.24 0.66 2.24  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.024 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.77 1.515 2.13 1.515 2.13 3.37 1.77 3.37  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0719 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.42 0.55 3.83 0.55 3.83 3.355 3.42 3.355  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.26 3.62 0.26 2.545 0.49 2.545 0.49 3.62 2.52 3.62 2.52 2.53 2.75 2.53 2.75 3.62 3.19 3.62 4.56 3.62 4.56 2.53 4.79 2.53 4.79 3.62 5.04 3.62 5.04 4.22 3.19 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.04 -0.3 5.04 0.3 4.79 0.3 4.79 0.765 4.56 0.765 4.56 0.3 2.53 0.3 2.53 0.69 2.3 0.69 2.3 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.195 0.55 1.51 0.55 1.51 0.93 3.19 0.93 3.19 1.755 2.96 1.755 2.96 1.165 1.51 1.165 1.51 3.355 1.28 3.355 1.28 0.78 0.195 0.78  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and2_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 9.52 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.055 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.03 1.21 3.515 1.21 3.515 1.56 1.03 1.56  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.055 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.8 4.125 1.8 4.125 2.15 0.54 2.15  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.0696 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.47 2.33 7.005 2.33 7.37 2.33 7.37 1.245 5.39 1.245 5.39 0.825 5.73 0.825 5.73 0.92 7.37 0.92 7.37 0.55 7.93 0.55 7.93 3.38 7.51 3.38 7.51 2.71 7.005 2.71 5.81 2.71 5.81 3.38 5.47 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.285 3.62 2.285 3.04 2.515 3.04 2.515 3.62 4.325 3.62 4.325 3.04 4.555 3.04 4.555 3.62 6.545 3.62 6.545 3.04 6.775 3.04 6.775 3.62 7.005 3.62 8.585 3.62 8.585 2.53 8.815 2.53 8.815 3.62 9.52 3.62 9.52 4.22 7.005 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 9.52 -0.3 9.52 0.3 9.035 0.3 9.035 0.905 8.805 0.905 8.805 0.3 6.85 0.3 6.85 0.64 6.51 0.64 6.51 0.3 4.555 0.3 4.555 0.765 4.325 0.765 4.325 0.3 0.475 0.3 0.475 0.905 0.245 0.905 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.21 2.53 4.765 2.53 4.765 1.23 3.865 1.23 3.865 0.825 2.265 0.825 2.265 0.595 4.095 0.595 4.095 0.995 4.995 0.995 4.995 1.585 7.005 1.585 7.005 1.815 4.995 1.815 4.995 2.76 3.59 2.76 3.59 3.38 3.25 3.38 3.25 2.76 1.55 2.76 1.55 3.38 1.21 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and2_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4955 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.77 1.25 1.77 1.25 1.12 1.57 1.12 1.57 2.15 0.54 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4955 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.12 2.12 1.12 2.12 2.415 1.8 2.415  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4955 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.36 1.12 2.91 1.12 2.91 2.415 2.36 2.415  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8756 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.57 0.65 5.01 0.65 5.01 3.38 4.57 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.21 3.62 1.21 3.285 1.55 3.285 1.55 3.62 3.745 3.62 3.745 2.53 3.975 2.53 3.975 3.62 4.315 3.62 5.6 3.62 5.6 4.22 4.315 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 3.875 0.3 3.875 1.09 3.645 1.09 3.645 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 2.825 3.185 2.825 3.185 0.805 0.53 0.805 0.53 1.035 0.19 1.035 0.19 0.575 3.415 0.575 3.415 1.46 4.315 1.46 4.315 1.8 3.415 1.8 3.415 3.055 2.57 3.055 2.57 3.34 2.23 3.34 2.23 3.055 0.53 3.055 0.53 3.34 0.19 3.34  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and3_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.16 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9815 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.16 1.02 1.16 1.02 2.29 0.66 2.29  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9815 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 1.16 2.14 1.16 2.14 2.29 1.78 2.29  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9815 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.865 1.16 3.26 1.16 3.26 2.29 2.865 2.29  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.48 0.65 4.95 0.65 4.95 3.38 4.48 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.32 3.62 1.32 3.16 1.55 3.16 1.55 3.62 3.36 3.62 3.36 3.16 3.59 3.16 3.59 3.62 4.25 3.62 5.58 3.62 5.58 2.53 5.81 2.53 5.81 3.62 6.16 3.62 6.16 4.22 4.25 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.16 -0.3 6.16 0.3 5.83 0.3 5.83 0.765 5.6 0.765 5.6 0.3 3.59 0.3 3.59 0.765 3.36 0.765 3.36 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.655 1.285 2.655 1.285 0.865 0.235 0.865 0.235 0.635 1.515 0.635 1.515 2.655 4.02 2.655 4.02 1.445 4.25 1.445 4.25 2.91 0.585 2.91 0.585 3.355 0.245 3.355  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and3_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 11.2 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.132 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.165 1.24 5.025 1.24 5.025 1.56 2.165 1.56  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.132 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.79 1.8 5.38 1.8 5.38 2.125 1.79 2.125  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.132 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.465 1.8 1.22 1.8 1.22 1.025 1.56 1.025 1.56 2.355 5.695 2.355 5.695 1.62 6.11 1.62 6.11 2.585 1.22 2.585 1.22 2.125 0.465 2.125  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.0592 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.55 2.385 9.26 2.385 9.61 2.385 9.61 1.1 7.25 1.1 7.25 0.81 7.59 0.81 7.59 0.87 9.545 0.87 9.545 0.55 9.99 0.55 9.99 3.34 9.59 3.34 9.59 2.725 9.26 2.725 7.89 2.725 7.89 3.34 7.55 3.34  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.23 3.62 2.23 3.285 2.57 3.285 2.57 3.62 4.27 3.62 4.27 3.285 4.61 3.285 4.61 3.62 6.53 3.62 6.53 3.285 6.87 3.285 6.87 3.62 8.57 3.62 8.57 3.285 8.91 3.285 8.91 3.62 9.26 3.62 10.665 3.62 10.665 2.53 10.895 2.53 10.895 3.62 11.2 3.62 11.2 4.22 9.26 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 11.2 -0.3 11.2 0.3 10.895 0.3 10.895 0.905 10.665 0.905 10.665 0.3 8.71 0.3 8.71 0.64 8.37 0.64 8.37 0.3 6.415 0.3 6.415 0.765 6.185 0.765 6.185 0.3 0.555 0.3 0.555 0.695 0.325 0.695 0.325 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.21 2.825 6.625 2.825 6.625 1.285 5.5 1.285 5.5 0.76 3.25 0.76 3.25 0.53 5.755 0.53 5.755 1.055 6.855 1.055 6.855 1.5 9.26 1.5 9.26 1.84 6.855 1.84 6.855 3.055 1.21 3.055  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and3_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.16 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.77 1.56 1.77 1.56 2.19 1 2.19 1 3 0.66 3  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.015 1.21 2.13 1.21 2.13 2.41 1.79 2.41 1.79 1.54 1.015 1.54  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.36 1.21 3.43 1.21 3.43 1.57 2.7 1.57 2.7 2.41 2.36 2.41  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.215 1.8 4.78 1.8 4.78 2.12 3.215 2.12  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8954 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.66 0.61 6.03 0.61 6.03 3.35 5.66 3.35  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.25 3.62 0.25 3.285 0.59 3.285 0.59 3.62 2.29 3.62 2.29 3.285 2.63 3.285 2.63 3.62 4.55 3.62 4.55 3.285 4.89 3.285 4.89 3.62 5.385 3.62 6.16 3.62 6.16 4.22 5.385 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.16 -0.3 6.16 0.3 4.845 0.3 4.845 1.035 4.505 1.035 4.505 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.27 2.825 5.155 2.825 5.155 1.505 3.77 1.505 3.77 0.76 0.535 0.76 0.535 1.09 0.305 1.09 0.305 0.53 4 0.53 4 1.265 5.385 1.265 5.385 3.055 3.65 3.055 3.65 3.39 3.31 3.39 3.31 3.055 1.61 3.055 1.61 3.39 1.27 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and4_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.28 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9195 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.12 1.77 0.63 1.77 0.63 1.03 1 1.03 1 2.15 0.12 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9195 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.23 1.77 1.75 1.77 1.75 1.03 2.12 1.03 2.12 2.15 1.23 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9195 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.35 1.77 2.87 1.77 2.87 1.03 3.24 1.03 3.24 2.15 2.35 2.15  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9195 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.47 1.77 4.595 1.77 4.595 2.15 3.47 2.15  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.495 0.805 6.07 0.805 6.07 3.235 5.495 3.235  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.3 3.62 0.3 3.16 0.53 3.16 0.53 3.62 2.285 3.62 2.285 3.28 2.625 3.28 2.625 3.62 4.325 3.62 4.325 3.285 4.665 3.285 4.665 3.62 5.23 3.62 6.6 3.62 6.6 2.65 6.83 2.65 6.83 3.62 7.28 3.62 7.28 4.22 5.23 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.28 -0.3 7.28 0.3 6.85 0.3 6.85 0.765 6.62 0.765 6.62 0.3 4.665 0.3 4.665 0.635 4.325 0.635 4.325 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.26 2.79 5 2.79 5 1.095 3.845 1.095 3.845 0.78 0.235 0.78 0.235 0.55 4.075 0.55 4.075 0.865 5.23 0.865 5.23 3.02 1.26 3.02  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and4_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__and4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__and4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.215 1.77 2.34 1.77 2.34 1.445 3.87 1.445 3.87 1.675 2.57 1.675 2.57 2.135 1.215 2.135  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.825 1.905 5.42 1.905 5.42 1.8 7.545 1.8 7.545 2.135 2.825 2.135  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 0.68 3.89 0.68 3.89 0.985 4.235 0.985 4.235 0.99 7.17 0.99 7.17 1.38 6.83 1.38 6.83 1.22 4.005 1.22 4.005 1.215 2.05 1.215 2.05 1.385 0.96 1.385  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.884 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 1.77 0.985 1.77 0.985 2.365 7.96 2.365 7.96 1.645 8.28 1.645 8.28 2.595 0.14 2.595  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.54 2.38 11.55 2.38 11.85 2.38 11.85 1.1 9.485 1.1 9.485 0.53 9.825 0.53 9.825 0.87 11.725 0.87 11.725 0.53 12.23 0.53 12.23 2.725 11.945 2.725 11.945 3.195 11.58 3.195 11.58 2.725 11.55 2.725 9.905 2.725 9.905 3.195 9.54 3.195  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.26 3.62 0.26 3.005 0.49 3.005 0.49 3.62 2.245 3.62 2.245 3.285 2.585 3.285 2.585 3.62 4.285 3.62 4.285 3.285 4.625 3.285 4.625 3.62 6.325 3.62 6.325 3.285 6.665 3.285 6.665 3.62 8.365 3.62 8.365 3.285 8.705 3.285 8.705 3.62 10.585 3.62 10.585 3.215 10.925 3.215 10.925 3.62 11.55 3.62 12.68 3.62 12.68 2.69 12.91 2.69 12.91 3.62 13.44 3.62 13.44 4.22 11.55 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 13.13 0.3 13.13 0.905 12.9 0.905 12.9 0.3 10.945 0.3 10.945 0.64 10.605 0.64 10.605 0.3 8.65 0.3 8.65 0.695 8.42 0.695 8.42 0.3 0.49 0.3 0.49 0.765 0.26 0.765 0.26 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.185 2.825 8.86 2.825 8.86 1.155 7.96 1.155 7.96 0.76 4.285 0.76 4.285 0.53 8.19 0.53 8.19 0.925 9.09 0.925 9.09 1.525 11.55 1.525 11.55 1.755 9.09 1.755 9.09 3.055 1.185 3.055  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__and4_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__antenna
  CLASS core ANTENNACELL ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__antenna 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 1.12 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNADIFFAREA 0.4104 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 0.81 0.475 0.81 0.475 2.71 0.14 2.71  ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.12 3.62 1.12 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 1.12 -0.3 1.12 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__antenna

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi21_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.775 1.77 2.34 1.77 2.34 1.16 2.68 1.16 2.68 2.15 1.775 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.115 1.77 0.66 1.77 0.66 1.16 1.01 1.16 1.01 2.15 0.115 2.15  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9135 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.91 1.77 3.475 1.77 3.475 1.16 3.815 1.16 3.815 2.15 2.91 2.15  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1456 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.24 0.55 2.58 0.55 2.58 0.87 1.545 0.87 1.545 2.725 1.24 2.725  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.57 3.62 3.525 3.62 3.525 2.69 3.755 2.69 3.755 3.62 4.48 3.62 4.48 4.22 2.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 3.855 0.3 3.855 0.765 3.625 0.765 3.625 0.3 0.475 0.3 0.475 0.765 0.245 0.765 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 2.495 0.53 2.495 0.53 3.16 2.23 3.16 2.23 2.495 2.57 2.495 2.57 3.39 0.19 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi21_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi21_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.28 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.24 6.725 1.24 6.725 1.56 4 1.56  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.29 1.4 3.63 1.4 3.63 1.8 6.725 1.8 6.725 2.12 3.29 2.12  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.893 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.58 1.8 2.28 1.8 2.28 2.125 0.58 2.125  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.0819 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.97 2.36 5.955 2.36 5.955 2.7 2.65 2.7 2.65 1.1 0.97 1.1 0.97 0.56 2.245 0.56 2.245 0.87 3.095 0.87 3.095 0.575 4.975 0.575 4.975 0.805 3.325 0.805 3.325 1.1 2.97 1.1  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.33 3.62 1.33 3.04 1.56 3.04 1.56 3.62 6.88 3.62 7.28 3.62 7.28 4.22 6.88 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.28 -0.3 7.28 0.3 6.88 0.3 6.88 0.765 6.65 0.765 6.65 0.3 2.835 0.3 2.835 0.64 2.495 0.64 2.495 0.3 0.54 0.3 0.54 0.765 0.31 0.765 0.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.31 2.53 2.035 2.53 2.035 3.095 6.65 3.095 6.65 2.435 6.88 2.435 6.88 3.325 1.8 3.325 1.8 2.76 0.54 2.76 0.54 3.38 0.31 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi21_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi21_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.368 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.8 6.42 1.8 6.42 2.12 0.6 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.368 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.21 3.465 1.21 3.465 1.325 7.065 1.325 7.065 1.805 8.35 1.805 8.35 2.12 6.835 2.12 6.835 1.57 0.6 1.57  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.624 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.295 1.79 12.79 1.79 12.79 2.15 9.295 2.15  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.8792 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.41 2.38 8.58 2.38 8.58 1.475 7.765 1.475 7.765 1.095 3.87 1.095 3.87 0.825 2.37 0.825 2.37 0.595 4.1 0.595 4.1 0.865 7.995 0.865 7.995 1.245 9.605 1.245 9.605 0.655 9.835 0.655 9.835 1.245 11.845 1.245 11.845 0.655 12.075 0.655 12.075 1.56 8.87 1.56 8.87 2.765 1.41 2.765  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 9.85 3.62 9.85 3.04 10.19 3.04 10.19 3.62 11.89 3.62 11.89 3.04 12.23 3.04 12.23 3.62 13.25 3.62 13.44 3.62 13.44 4.22 13.25 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 13.195 0.3 13.195 1.215 12.965 1.215 12.965 0.3 11.01 0.3 11.01 1.015 10.67 1.015 10.67 0.3 8.59 0.3 8.59 0.98 8.25 0.98 8.25 0.3 4.67 0.3 4.67 0.635 4.33 0.635 4.33 0.3 0.695 0.3 0.695 0.69 0.465 0.69 0.465 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.445 2.54 0.675 2.54 0.675 3.16 9.235 3.16 9.235 2.53 13.25 2.53 13.25 3.38 12.91 3.38 12.91 2.76 11.21 2.76 11.21 3.38 10.87 3.38 10.87 2.76 9.565 2.76 9.565 3.39 0.445 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi21_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi211_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0335 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.77 1.23 2.15 1.23 2.15 1.77 2.69 1.77 2.69 2.15 1.77 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0335 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.16 1 1.16 1 2.19 0.65 2.19  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8865 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 1.73 3.22 1.73 3.22 2.85 4.01 2.85 4.01 3.31 2.92 3.31  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8865 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 1.77 4.95 1.77 4.95 2.15 3.45 2.15  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.2599 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.24 0.56 3.28 0.56 3.28 1.045 4.63 1.045 4.63 0.565 4.86 0.565 4.86 1.275 3.05 1.275 3.05 1 1.54 1 1.54 2.725 1.24 2.725  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.52 3.62 4.53 3.62 4.53 2.53 4.76 2.53 4.76 3.62 5.6 3.62 5.6 4.22 2.52 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 3.74 0.3 3.74 0.815 3.51 0.815 3.51 0.3 0.48 0.3 0.48 0.87 0.25 0.87 0.25 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 2.53 0.48 2.53 0.48 3.15 2.29 3.15 2.29 2.53 2.52 2.53 2.52 3.38 0.25 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi211_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi211_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 9.52 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.076 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.16 1.24 3.31 1.24 3.31 1.56 1.16 1.56  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.076 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.42 1.8 3.77 1.8 3.77 2.12 0.42 2.12  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.758 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.8 5.22 1.8 5.22 2.36 7.885 2.36 7.885 1.8 9.025 1.8 9.025 2.12 8.43 2.12 8.43 2.595 5.665 2.595 5.665 2.71 4.6 2.71  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.758 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.65 1.8 7.395 1.8 7.395 2.12 5.65 2.12  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1268 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.17 2.36 4.04 2.36 4.04 1.56 3.655 1.56 3.655 1 2.15 1 2.15 0.68 3.915 0.68 3.915 1.24 4.915 1.24 4.915 0.87 5.41 0.87 5.41 0.56 5.75 0.56 5.75 0.87 7.65 0.87 7.65 0.56 7.99 0.56 7.99 1.1 5.145 1.1 5.145 1.56 4.36 1.56 4.36 2.78 1.17 2.78  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 6.45 3.62 6.45 3.285 6.79 3.285 6.79 3.62 8.955 3.62 9.52 3.62 9.52 4.22 8.955 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 9.52 -0.3 9.52 0.3 9.055 0.3 9.055 0.695 8.825 0.695 8.825 0.3 6.87 0.3 6.87 0.64 6.53 0.64 6.53 0.3 4.395 0.3 4.395 0.69 4.165 0.69 4.165 0.3 0.475 0.3 0.475 0.91 0.245 0.91 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.5 0.475 2.5 0.475 3.16 5.91 3.16 5.91 2.825 8.725 2.825 8.725 2.5 8.955 2.5 8.955 3.39 8.725 3.39 8.725 3.055 6.14 3.055 6.14 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi211_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi211_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.288 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.71 1.21 3.83 1.21 3.83 1.34 7.935 1.34 7.935 1.57 1.71 1.57  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.288 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.44 1.8 9.035 1.8 9.035 2.12 1.44 2.12  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.544 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.55 1.8 10.57 1.8 10.57 2.36 13.53 2.36 13.53 1.965 13.87 1.965 13.87 2.36 15.205 2.36 15.205 1.965 15.545 1.965 15.545 2.36 18.57 2.36 18.57 1.8 19.59 1.8 19.59 2.12 18.8 2.12 18.8 2.595 10.34 2.595 10.34 2.12 9.55 2.12  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.544 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.84 1.505 18.25 1.505 18.25 2.13 16.08 2.13 16.08 1.735 10.84 1.735  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.2952 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.98 0.955 1.19 0.955 1.19 0.7 2.9 0.7 2.9 0.53 3.24 0.53 3.24 0.7 4.71 0.7 4.71 0.87 6.98 0.87 6.98 0.575 7.32 0.575 7.32 0.87 8.735 0.87 8.735 1.045 10.36 1.045 10.36 0.775 10.7 0.775 10.7 1.045 13.04 1.045 13.04 0.775 13.38 0.775 13.38 1.045 15.72 1.045 15.72 0.775 16.06 0.775 16.06 1.045 18.4 1.045 18.4 0.775 18.74 0.775 18.74 1.275 8.505 1.275 8.505 1.1 4.48 1.1 4.48 0.93 1.42 0.93 1.42 1.185 1.21 1.185 1.21 2.36 8.34 2.36 8.34 2.68 0.98 2.68  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 11.7 3.62 11.7 3.285 12.04 3.285 12.04 3.62 16.975 3.62 16.975 3.285 17.315 3.285 17.315 3.62 19.755 3.62 20.16 3.62 20.16 4.22 19.755 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 19.805 0.3 19.805 1.06 19.575 1.06 19.575 0.3 17.4 0.3 17.4 0.765 17.06 0.765 17.06 0.3 14.72 0.3 14.72 0.765 14.38 0.765 14.38 0.3 12.04 0.3 12.04 0.71 11.7 0.71 11.7 0.3 9.36 0.3 9.36 0.765 9.02 0.765 9.02 0.3 5.28 0.3 5.28 0.64 4.94 0.64 4.94 0.3 0.96 0.3 0.96 0.71 0.62 0.71 0.62 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.86 3.16 9.07 3.16 9.07 2.53 9.41 2.53 9.41 2.825 19.525 2.825 19.525 2.53 19.755 2.53 19.755 3.38 19.525 3.38 19.525 3.055 9.41 3.055 9.41 3.39 0.86 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi211_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi22_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.04 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 0.55 3.24 0.55 3.24 2.15 2.92 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.48 0.55 3.8 0.55 3.8 1.8 4.545 1.8 4.545 2.15 3.48 2.15  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.55 2.12 0.55 2.12 2.15 1.8 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0965 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.61 1.085 1.005 1.085 1.005 1.77 1.57 1.77 1.57 2.15 0.61 2.15  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.35 0.585 2.68 0.585 2.68 2.38 3.89 2.38 3.89 2.71 2.35 2.71  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.33 3.62 1.33 3.04 1.56 3.04 1.56 3.62 4.675 3.62 5.04 3.62 5.04 4.22 4.675 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.04 -0.3 5.04 0.3 4.62 0.3 4.62 0.905 4.39 0.905 4.39 0.3 0.54 0.3 0.54 0.725 0.31 0.725 0.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.255 2.53 2.05 2.53 2.05 3.145 4.335 3.145 4.335 2.53 4.675 2.53 4.675 3.38 1.82 3.38 1.82 2.76 0.595 2.76 0.595 3.38 0.255 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi22_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi22_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.96 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.193 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.69 1.21 8.38 1.21 8.38 1.57 5.69 1.57  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.193 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.95 1.4 5.235 1.4 5.235 1.8 8.38 1.8 8.38 2.12 4.95 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.193 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.61 2.09 0.61 2.09 1.59 1.65 1.59 1.65 1.03 0.94 1.03  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.193 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.82 4.03 1.82 4.03 2.12 0.62 2.12  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.139725 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.72 2.36 7.67 2.36 7.67 2.78 4.345 2.78 4.345 1.15 2.32 1.15 2.32 0.715 2.555 0.715 2.555 0.87 4.925 0.87 4.925 0.64 6.65 0.64 6.65 0.87 5.155 0.87 5.155 1.1 4.72 1.1  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 3.16 1.495 3.16 1.495 3.62 3.305 3.62 3.305 3.16 3.535 3.16 3.535 3.62 8.69 3.62 8.96 3.62 8.96 4.22 8.69 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.96 -0.3 8.96 0.3 8.635 0.3 8.635 0.905 8.405 0.905 8.405 0.3 4.61 0.3 4.61 0.64 4.27 0.64 4.27 0.3 0.475 0.3 0.475 0.905 0.245 0.905 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 2.53 4.025 2.53 4.025 3.13 8.35 3.13 8.35 2.475 8.69 2.475 8.69 3.365 3.795 3.365 3.795 2.76 2.57 2.76 2.57 3.38 2.23 3.38 2.23 2.76 0.53 2.76 0.53 3.38 0.19 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi22_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi22_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.92 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.18 1.8 14.73 1.8 14.73 2.12 11.18 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.445 1.71 10.16 1.71 10.16 1.24 13.78 1.24 13.78 0.53 17.05 0.53 17.05 2.235 16.82 2.235 16.82 0.76 14.01 0.76 14.01 1.56 10.52 1.56 10.52 2.14 9.445 2.14  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 1.8 7.24 1.8 7.24 2.13 1.64 2.13  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.23 3.375 1.23 3.375 1.325 8.12 1.325 8.12 1.56 1.02 1.56 1.02 2.225 0.62 2.225  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.389 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.215 2.67 15.05 2.67 15.05 0.99 15.58 0.99 15.58 2.67 16.67 2.67 16.67 2.91 8.985 2.91 8.985 1.095 3.765 1.095 3.765 0.8 2.225 0.8 2.225 0.57 3.995 0.57 3.995 0.865 6.365 0.865 6.365 0.57 6.595 0.57 6.595 0.865 8.985 0.865 8.985 0.53 11.18 0.53 11.18 1 9.215 1  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.21 3.62 1.21 3.01 1.55 3.01 1.55 3.62 3.25 3.62 3.25 3.01 3.59 3.01 3.59 3.62 5.29 3.62 5.29 3.01 5.63 3.01 5.63 3.62 7.33 3.62 7.33 3.01 7.67 3.01 7.67 3.62 17.65 3.62 17.92 3.62 17.92 4.22 17.65 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.92 -0.3 17.92 0.3 17.595 0.3 17.595 0.73 17.365 0.73 17.365 0.3 13.075 0.3 13.075 0.73 12.845 0.73 12.845 0.3 8.69 0.3 8.69 0.635 8.35 0.635 8.35 0.3 4.61 0.3 4.61 0.635 4.27 0.635 4.27 0.3 0.475 0.3 0.475 0.695 0.245 0.695 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 2.485 8.69 2.485 8.69 3.16 17.31 3.16 17.31 2.485 17.65 2.485 17.65 3.39 8.35 3.39 8.35 2.715 6.65 2.715 6.65 3.39 6.31 3.39 6.31 2.715 4.61 2.715 4.61 3.39 4.27 3.39 4.27 2.715 2.57 2.715 2.57 3.39 2.23 3.39 2.23 2.715 0.53 2.715 0.53 3.39 0.19 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi22_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi221_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.16 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0335 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.15 1.16 5.51 1.16 5.51 2.3 5.15 2.3  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0335 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.005 1.585 4.37 1.585 4.37 2.835 4.005 2.835  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0335 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.75 1.21 2.15 1.21 2.15 1.78 2.69 1.78 2.69 2.15 1.75 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0335 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.12 1.77 0.68 1.77 0.68 1.16 1.07 1.16 1.07 2.15 0.12 2.15  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8865 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 1.55 3.24 1.55 3.24 3.32 2.92 3.32  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.4892 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.15 0.675 3.18 0.675 3.18 0.975 4.6 0.975 4.6 0.675 5.98 0.675 5.98 0.905 4.92 0.905 4.92 2.865 4.6 2.865 4.6 1.205 2.95 1.205 2.95 0.905 2.15 0.905  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3.16 1.595 3.16 1.595 3.62 2.67 3.62 5.915 3.62 6.16 3.62 6.16 4.22 5.915 4.22 2.67 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.16 -0.3 6.16 0.3 4.01 0.3 4.01 0.745 3.67 0.745 3.67 0.3 0.53 0.3 0.53 0.815 0.19 0.815 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.28 2.59 2.67 2.59 2.67 3.38 2.33 3.38 2.33 2.93 0.63 2.93 0.63 3.38 0.28 3.38  ;
        POLYGON 3.545 2.53 3.775 2.53 3.775 3.15 5.685 3.15 5.685 2.53 5.915 2.53 5.915 3.38 3.545 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi221_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi221_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.88 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.08 1.55 9.31 1.55 9.31 1.79 12.05 1.79 12.05 2.12 9.08 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.57 1.225 12.05 1.225 12.05 1.56 9.57 1.56  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.125 1.91 5.65 1.91 5.65 1.8 7.815 1.8 7.815 2.14 4.125 2.14  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.978 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.525 1.785 3.04 1.785 3.04 1.45 5.39 1.45 5.39 1.68 3.27 1.68 3.27 2.15 0.525 2.15  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.708 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 1.325 2.58 1.325 2.58 0.99 6 0.99 6 1.21 8.31 1.21 8.31 1.56 5.77 1.56 5.77 1.22 2.81 1.22 2.81 1.555 0.87 1.555  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.496525 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 0.705 0.475 0.705 0.475 0.865 2.12 0.865 2.12 0.53 6.495 0.53 6.495 0.705 7.35 0.705 7.35 0.565 8.845 0.565 8.845 2.36 12.32 2.36 12.32 0.7 12.55 0.7 12.55 2.795 8.565 2.795 8.565 0.935 6.265 0.935 6.265 0.76 2.35 0.76 2.35 1.095 0.245 1.095  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.55 3.62 2.55 3.445 2.89 3.445 2.89 3.62 5.05 3.62 5.05 3.445 5.39 3.445 5.39 3.62 12.505 3.62 12.88 3.62 12.88 4.22 12.505 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.88 -0.3 12.88 0.3 10.645 0.3 10.645 0.635 10.305 0.635 10.305 0.3 7.065 0.3 7.065 0.475 6.725 0.475 6.725 0.3 1.87 0.3 1.87 0.635 1.53 0.635 1.53 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.31 2.525 7.41 2.525 7.41 2.755 1.31 2.755  ;
        POLYGON 0.345 2.46 0.575 2.46 0.575 3.12 2.075 3.12 2.075 2.985 6.195 2.985 6.195 3.135 8.105 3.135 8.105 2.46 8.335 2.46 8.335 3.135 12.505 3.135 12.505 3.365 5.855 3.365 5.855 3.215 2.29 3.215 2.29 3.35 0.345 3.35  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi221_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi221_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.278 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.12 1.335 20.72 1.335 20.72 1.22 21.865 1.22 21.865 1.57 17.39 1.57 17.39 1.675 14.55 1.675 14.55 2.245 14.12 2.245  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.278 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.98 1.91 18.01 1.91 18.01 1.8 21.865 1.8 21.865 2.14 14.98 2.14  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.918 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.2 1.59 1.2 1.59 1.33 3.38 1.33 3.38 1.24 5.63 1.24 5.63 1.555 8.31 1.555 8.31 1.79 3.38 1.79 3.38 1.56 0.62 1.56  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.918 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.465 1.8 3.125 1.8 3.125 2.04 7.29 2.04 7.29 2.27 2.71 2.27 2.71 2.12 0.465 2.12  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.582 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.82 1.8 13.16 1.8 13.16 2.12 8.82 2.12  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.3055 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.19 0.73 2.05 0.73 2.05 0.87 2.85 0.87 2.85 0.545 6.11 0.545 6.11 1.095 8.555 1.095 8.555 0.765 8.785 0.765 8.785 1.095 11.11 1.095 11.11 0.53 11.45 0.53 11.45 1.095 13.53 1.095 13.53 0.53 13.87 0.53 13.87 0.875 16.24 0.875 16.24 0.545 18.69 0.545 18.69 0.87 20.24 0.87 20.24 0.545 22.04 0.545 22.04 0.775 20.47 0.775 20.47 1.105 18.46 1.105 18.46 0.78 16.47 0.78 16.47 1.105 13.88 1.105 13.88 2.68 21.05 2.68 21.05 2.91 13.53 2.91 13.53 1.56 8.905 1.56 8.905 1.325 5.88 1.325 5.88 0.78 3.08 0.78 3.08 1.1 1.82 1.1 1.82 0.96 0.19 0.96  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.24 3.62 0.24 2.53 0.58 2.53 0.58 3.62 2.335 3.62 2.335 3.04 2.565 3.04 2.565 3.62 4.375 3.62 4.375 3.04 4.605 3.04 4.605 3.62 6.415 3.62 6.415 3.04 6.645 3.04 6.645 3.62 8.455 3.62 8.455 3.04 8.685 3.04 8.685 3.62 21.975 3.62 22.4 3.62 22.4 4.22 21.975 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 19.99 0.3 19.99 0.64 19.65 0.64 19.65 0.3 15.91 0.3 15.91 0.64 15.57 0.64 15.57 0.3 12.515 0.3 12.515 0.795 12.285 0.795 12.285 0.3 10.275 0.3 10.275 0.795 10.045 0.795 10.045 0.3 6.7 0.3 6.7 0.795 6.36 0.795 6.36 0.3 2.62 0.3 2.62 0.64 2.28 0.64 2.28 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.26 2.53 12.56 2.53 12.56 2.76 7.72 2.76 7.72 3.38 7.38 3.38 7.38 2.76 5.68 2.76 5.68 3.38 5.34 3.38 5.34 2.76 3.64 2.76 3.64 3.38 3.3 3.38 3.3 2.76 1.6 2.76 1.6 3.38 1.26 3.38  ;
        POLYGON 9.11 3.16 21.745 3.16 21.745 2.5 21.975 2.5 21.975 3.39 9.11 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi221_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi222_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.84 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.84 1.23 7.18 1.23 7.18 2.33 7.72 2.33 7.72 2.71 6.84 2.71  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.14 2.33 5.72 2.33 5.72 1.535 6.04 1.535 6.04 2.71 5.14 2.71  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.35 1.77 3.8 1.77 3.8 2.15 2.35 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.04 1.105 4.36 1.105 4.36 1.77 4.95 1.77 4.95 2.15 4.04 2.15  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.55 2.12 0.55 2.12 2.235 1.8 2.235  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.072 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.48 1.77 1.24 1.77 1.24 0.55 1.56 0.55 1.56 2.15 0.48 2.15  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7565 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.51 0.55 4.895 0.55 4.895 0.865 5.88 0.865 5.88 0.67 7.635 0.67 7.635 1 6.6 1 6.6 2.77 6.28 2.77 6.28 1.095 4.665 1.095 4.665 0.78 2.51 0.78  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.685 2.53 0.685 3.62 2.44 3.62 2.44 3.04 2.67 3.04 2.67 3.62 7.635 3.62 7.84 3.62 7.84 4.22 7.635 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.84 -0.3 7.84 0.3 5.485 0.3 5.485 0.635 5.145 0.635 5.145 0.3 0.71 0.3 0.71 0.905 0.48 0.905 0.48 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.53 4.5 2.53 4.5 2.76 1.705 2.76 1.705 3.38 1.365 3.38  ;
        POLYGON 3.095 3.095 7.635 3.095 7.635 3.325 3.095 3.325  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi222_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi222_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.7 1.96 12.44 1.96 12.44 0.55 12.96 0.55 12.96 2.195 9.7 2.195  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.87 1.21 12.005 1.21 12.005 1.63 9.87 1.63  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.605 1.325 8.71 1.325 8.71 2.15 7.37 2.15 7.37 1.555 5.605 1.555  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.57 1.77 5.46 1.77 5.46 1.785 6.825 1.785 6.825 2.195 4.57 2.195  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.655 1.965 2.225 1.965 2.225 1.8 4.155 1.8 4.155 2.195 0.655 2.195  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.18 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.21 1.79 1.21 1.79 1.34 3.485 1.34 3.485 1.57 1.79 1.57 1.79 1.59 0.65 1.59  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.1688 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.225 0.74 2.25 0.74 2.25 0.865 4.925 0.865 4.925 0.845 5.265 0.845 5.265 0.865 9.05 0.865 9.05 0.79 9.47 0.79 9.47 2.44 13.255 2.44 13.255 0.57 13.485 0.57 13.485 2.67 9.05 2.67 9.05 1.095 2.02 1.095 2.02 0.97 0.225 0.97  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.225 3.62 0.225 2.53 0.565 2.53 0.565 3.62 2.32 3.62 2.32 3.04 2.55 3.04 2.55 3.62 4.36 3.62 4.36 3.04 4.59 3.04 4.59 3.62 13.55 3.62 14 3.62 14 4.22 13.55 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14 -0.3 14 0.3 11.5 0.3 11.5 0.635 11.16 0.635 11.16 0.3 7.405 0.3 7.405 0.635 7.065 0.635 7.065 0.3 2.795 0.3 2.795 0.635 2.455 0.635 2.455 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.245 2.53 8.425 2.53 8.425 2.76 3.625 2.76 3.625 3.38 3.285 3.38 3.285 2.76 1.585 2.76 1.585 3.38 1.245 3.38  ;
        POLYGON 5.02 3.16 13.55 3.16 13.55 3.39 5.02 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi222_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__aoi222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__aoi222_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 26.32 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.78 1.965 23.61 1.965 23.61 1.77 25.67 1.77 25.67 2.195 17.78 2.195  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.535 1.16 18.43 1.16 18.43 1.325 20.405 1.325 20.405 1.22 22.49 1.22 22.49 1.325 23.11 1.325 23.11 1.615 17.535 1.615  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.945 1.335 16.835 1.335 16.835 2.025 16.605 2.025 16.605 1.565 10.16 1.565 10.16 2.15 8.945 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.415 1.8 16.255 1.8 16.255 2.12 10.415 2.12  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.335 7.62 1.335 7.62 1.76 8.515 1.76 8.515 2.15 7.32 2.15 7.32 1.565 0.71 1.565  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.585 1.8 7.09 1.8 7.09 2.12 0.585 2.12  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.9406 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.19 0.865 5.86 0.865 5.86 0.87 6.805 0.87 6.805 0.865 15.81 0.865 15.81 0.57 19.04 0.57 19.04 0.865 19.875 0.865 19.875 0.53 23.065 0.53 23.065 0.865 24.73 0.865 24.73 0.65 25.73 0.65 25.73 1.095 22.835 1.095 22.835 0.76 20.105 0.76 20.105 1.095 18.81 1.095 18.81 0.8 17.305 0.8 17.305 2.605 24.71 2.605 24.71 2.835 17.075 2.835 17.075 0.8 16.04 0.8 16.04 1.095 7.035 1.095 7.035 1.1 5.63 1.1 5.63 1.095 0.19 1.095  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.19 3.62 0.19 2.555 0.53 2.555 0.53 3.62 2.23 3.62 2.23 3.04 2.575 3.04 2.575 3.62 4.27 3.62 4.27 3.04 4.61 3.04 4.61 3.62 6.31 3.62 6.31 3.04 6.65 3.04 6.65 3.62 8.35 3.62 8.35 3.04 8.69 3.04 8.69 3.62 25.73 3.62 26.32 3.62 26.32 4.22 25.73 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 26.32 -0.3 26.32 0.3 23.69 0.3 23.69 0.635 23.35 0.635 23.35 0.3 19.61 0.3 19.61 0.635 19.27 0.635 19.27 0.3 15.53 0.3 15.53 0.635 15.19 0.635 15.19 0.3 11.45 0.3 11.45 0.635 11.11 0.635 11.11 0.3 6.65 0.3 6.65 0.64 6.31 0.64 6.31 0.3 2.57 0.3 2.57 0.635 2.23 0.635 2.23 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.21 2.53 16.55 2.53 16.55 2.76 7.67 2.76 7.67 3.38 7.33 3.38 7.33 2.76 5.63 2.76 5.63 3.38 5.29 3.38 5.29 2.76 3.59 2.76 3.59 3.38 3.25 3.38 3.25 2.76 1.55 2.76 1.55 3.38 1.21 3.38  ;
        POLYGON 9.07 3.16 25.39 3.16 25.39 2.555 25.73 2.555 25.73 3.39 9.07 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__aoi222_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 3.36 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4985 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.65 1.22 0.65 1.22 1.63 1.59 1.63 1.59 2.19 0.705 2.19  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.33 0.575 2.955 0.575 2.955 3.38 2.485 3.38 2.485 1.6 2.33 1.6  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.53 3.62 1.53 3.13 1.87 3.13 1.87 3.62 2.255 3.62 3.36 3.62 3.36 4.22 2.255 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 3.36 -0.3 3.36 0.3 1.815 0.3 1.815 0.865 1.585 0.865 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.8 0.475 0.8 0.475 2.58 1.97 2.58 1.97 1.83 2.255 1.83 2.255 2.815 0.63 2.815 0.63 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.612 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.66 5.7 1.66 5.7 2.15 0.62 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.0968 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.085 2.33 12.805 2.33 13.32 2.33 13.32 1.42 8.085 1.42 8.085 0.675 8.345 0.675 8.345 0.98 10.325 0.98 10.325 0.675 10.555 0.675 10.555 0.98 12.565 0.98 12.565 0.675 12.795 0.675 12.795 0.98 14.805 0.98 14.805 0.675 15.035 0.675 15.035 0.98 17.045 0.98 17.045 0.675 17.275 0.675 17.275 0.98 19.285 0.98 19.285 0.53 19.515 0.53 19.515 1.42 14.12 1.42 14.12 2.33 19.415 2.33 19.415 3.38 19.185 3.38 19.185 2.93 17.175 2.93 17.175 3.38 16.945 3.38 16.945 2.93 14.935 2.93 14.935 3.38 14.705 3.38 14.705 2.93 12.805 2.93 12.695 2.93 12.695 3.38 12.465 3.38 12.465 2.93 10.455 2.93 10.455 3.38 10.225 3.38 10.225 2.93 8.315 2.93 8.315 3.38 8.085 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.385 3.62 2.385 3 2.615 3 2.615 3.62 4.625 3.62 4.625 3 4.855 3 4.855 3.62 6.865 3.62 6.865 2.53 7.095 2.53 7.095 3.62 9.105 3.62 9.105 3.17 9.335 3.17 9.335 3.62 11.345 3.62 11.345 3.17 11.575 3.17 11.575 3.62 12.805 3.62 13.585 3.62 13.585 3.17 13.815 3.17 13.815 3.62 15.825 3.62 15.825 3.17 16.055 3.17 16.055 3.62 18.065 3.62 18.065 3.17 18.295 3.17 18.295 3.62 20.26 3.62 20.305 3.62 20.305 2.53 20.535 2.53 20.535 3.62 21.28 3.62 21.28 4.22 20.26 4.22 12.805 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 20.69 0.3 20.69 0.765 20.35 0.765 20.35 0.3 18.45 0.3 18.45 0.71 18.11 0.71 18.11 0.3 16.21 0.3 16.21 0.71 15.87 0.71 15.87 0.3 13.97 0.3 13.97 0.71 13.63 0.71 13.63 0.3 11.73 0.3 11.73 0.71 11.39 0.71 11.39 0.3 9.49 0.3 9.49 0.71 9.15 0.71 9.15 0.3 7.25 0.3 7.25 0.765 6.91 0.765 6.91 0.3 5.01 0.3 5.01 0.765 4.67 0.765 4.67 0.3 2.77 0.3 2.77 0.765 2.43 0.765 2.43 0.3 0.53 0.3 0.53 0.765 0.19 0.765 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 2.53 6.26 2.53 6.26 1.25 1.365 1.25 1.365 0.675 1.595 0.675 1.595 1.015 3.605 1.015 3.605 0.675 3.835 0.675 3.835 1.015 5.845 1.015 5.845 0.675 6.075 0.675 6.075 1.015 6.495 1.015 6.495 1.685 12.805 1.685 12.805 2.025 6.495 2.025 6.495 2.76 5.975 2.76 5.975 3.38 5.745 3.38 5.745 2.76 3.735 2.76 3.735 3.38 3.505 3.38 3.505 2.76 1.495 2.76 1.495 3.38 1.265 3.38  ;
        POLYGON 14.625 1.685 20.26 1.685 20.26 2.03 14.625 2.03  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_12

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 28 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.816 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.71 8.185 1.71 8.185 2.15 0.62 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.4624 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.325 2.23 16.51 2.23 17.75 2.23 17.75 1.51 10.325 1.51 10.325 0.675 10.585 0.675 10.585 0.93 12.565 0.93 12.565 0.675 12.795 0.675 12.795 0.93 14.805 0.93 14.805 0.675 15.035 0.675 15.035 0.93 17.045 0.93 17.045 0.675 17.275 0.675 17.275 0.93 19.285 0.93 19.285 0.675 19.515 0.675 19.515 0.93 21.525 0.93 21.525 0.675 21.755 0.675 21.755 0.93 23.765 0.93 23.765 0.675 23.995 0.675 23.995 0.93 26.005 0.93 26.005 0.675 26.235 0.675 26.235 1.51 18.65 1.51 18.65 2.23 26.135 2.23 26.135 3.38 25.905 3.38 25.905 2.81 23.895 2.81 23.895 3.38 23.665 3.38 23.665 2.81 21.655 2.81 21.655 3.38 21.425 3.38 21.425 2.81 19.415 2.81 19.415 3.38 19.185 3.38 19.185 2.81 17.175 2.81 17.175 3.38 16.945 3.38 16.945 2.81 16.51 2.81 14.935 2.81 14.935 3.38 14.705 3.38 14.705 2.81 12.695 2.81 12.695 3.38 12.465 3.38 12.465 2.81 10.555 2.81 10.555 3.38 10.325 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.385 3.62 2.385 3 2.615 3 2.615 3.62 4.625 3.62 4.625 3 4.855 3 4.855 3.62 6.865 3.62 6.865 3 7.095 3 7.095 3.62 9.105 3.62 9.105 2.53 9.335 2.53 9.335 3.62 11.345 3.62 11.345 3.04 11.575 3.04 11.575 3.62 13.585 3.62 13.585 3.04 13.815 3.04 13.815 3.62 15.825 3.62 15.825 3.04 16.055 3.04 16.055 3.62 16.51 3.62 18.065 3.62 18.065 3.04 18.295 3.04 18.295 3.62 20.305 3.62 20.305 3.04 20.535 3.04 20.535 3.62 22.545 3.62 22.545 3.04 22.775 3.04 22.775 3.62 24.785 3.62 24.785 3.04 25.015 3.04 25.015 3.62 26.98 3.62 27.025 3.62 27.025 2.53 27.255 2.53 27.255 3.62 28 3.62 28 4.22 26.98 4.22 16.51 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 28 -0.3 28 0.3 27.41 0.3 27.41 0.765 27.07 0.765 27.07 0.3 25.17 0.3 25.17 0.7 24.83 0.7 24.83 0.3 22.93 0.3 22.93 0.7 22.59 0.7 22.59 0.3 20.69 0.3 20.69 0.7 20.35 0.7 20.35 0.3 18.45 0.3 18.45 0.7 18.11 0.7 18.11 0.3 16.21 0.3 16.21 0.7 15.87 0.7 15.87 0.3 13.97 0.3 13.97 0.7 13.63 0.7 13.63 0.3 11.73 0.3 11.73 0.7 11.39 0.7 11.39 0.3 9.49 0.3 9.49 0.765 9.15 0.765 9.15 0.3 7.25 0.3 7.25 0.765 6.91 0.765 6.91 0.3 5.01 0.3 5.01 0.765 4.67 0.765 4.67 0.3 2.77 0.3 2.77 0.765 2.43 0.765 2.43 0.3 0.53 0.3 0.53 0.765 0.19 0.765 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 2.53 8.535 2.53 8.535 1.25 1.365 1.25 1.365 0.675 1.595 0.675 1.595 1.015 3.605 1.015 3.605 0.675 3.835 0.675 3.835 1.015 5.845 1.015 5.845 0.675 6.075 0.675 6.075 1.015 8.085 1.015 8.085 0.675 8.315 0.675 8.315 1.015 8.77 1.015 8.77 1.74 16.51 1.74 16.51 1.97 8.77 1.97 8.77 2.76 8.215 2.76 8.215 3.38 7.985 3.38 7.985 2.76 5.975 2.76 5.975 3.38 5.745 3.38 5.745 2.76 3.735 2.76 3.735 3.38 3.505 3.38 3.505 2.76 1.495 2.76 1.495 3.38 1.265 3.38  ;
        POLYGON 19.56 1.74 26.98 1.74 26.98 1.97 19.56 1.97  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_16

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.61 1.015 0.61 1.015 1.625 1.65 1.625 1.65 2.15 0.705 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.675 2.21 3.24 2.21 3.48 2.21 3.48 1.3 2.675 1.3 2.675 0.57 2.905 0.57 2.905 1.065 3.8 1.065 3.8 2.7 3.24 2.7 2.905 2.7 2.905 3.39 2.675 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.405 3.62 1.405 3.01 1.745 3.01 1.745 3.62 3.24 3.62 3.64 3.62 3.64 3.01 3.98 3.01 3.98 3.62 4.48 3.62 4.48 4.22 3.24 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 4.08 0.3 4.08 0.765 3.74 0.765 3.74 0.3 1.745 0.3 1.745 0.765 1.405 0.765 1.405 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.57 0.475 0.57 0.475 2.39 1.9 2.39 1.9 1.55 3.24 1.55 3.24 1.89 2.13 1.89 2.13 2.625 0.475 2.625 0.475 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 34.72 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 11.02 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.74 9.9 1.74 9.9 2.15 0.63 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 11.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.565 2.27 21.57 2.27 22.23 2.27 22.23 1.51 12.565 1.51 12.565 0.675 12.825 0.675 12.825 0.865 14.805 0.865 14.805 0.675 15.035 0.675 15.035 0.865 17.045 0.865 17.045 0.675 17.275 0.675 17.275 0.865 19.285 0.865 19.285 0.675 19.515 0.675 19.515 0.865 21.525 0.865 21.525 0.675 21.755 0.675 21.755 0.865 23.765 0.865 23.765 0.675 23.995 0.675 23.995 0.865 26.005 0.865 26.005 0.675 26.235 0.675 26.235 0.865 28.245 0.865 28.245 0.675 28.475 0.675 28.475 0.865 30.485 0.865 30.485 0.675 30.715 0.675 30.715 0.865 32.725 0.865 32.725 0.675 32.955 0.675 32.955 1.51 23.13 1.51 23.13 2.27 32.855 2.27 32.855 3.38 32.625 3.38 32.625 3 30.615 3 30.615 3.38 30.385 3.38 30.385 3 28.375 3 28.375 3.38 28.145 3.38 28.145 3 26.135 3 26.135 3.38 25.905 3.38 25.905 3 23.895 3 23.895 3.38 23.665 3.38 23.665 3 21.655 3 21.655 3.38 21.57 3.38 21.425 3.38 21.425 3 19.415 3 19.415 3.38 19.185 3.38 19.185 3 17.175 3 17.175 3.38 16.945 3.38 16.945 3 14.935 3 14.935 3.38 14.705 3.38 14.705 3 12.795 3 12.795 3.38 12.565 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.385 3.62 2.385 3 2.615 3 2.615 3.62 4.625 3.62 4.625 3 4.855 3 4.855 3.62 6.865 3.62 6.865 3 7.095 3 7.095 3.62 9.105 3.62 9.105 3 9.335 3 9.335 3.62 11.345 3.62 11.345 2.53 11.575 2.53 11.575 3.62 13.585 3.62 13.585 3.23 13.815 3.23 13.815 3.62 15.825 3.62 15.825 3.23 16.055 3.23 16.055 3.62 18.065 3.62 18.065 3.23 18.295 3.23 18.295 3.62 20.305 3.62 20.305 3.23 20.535 3.23 20.535 3.62 21.57 3.62 22.545 3.62 22.545 3.23 22.775 3.23 22.775 3.62 24.785 3.62 24.785 3.23 25.015 3.23 25.015 3.62 27.025 3.62 27.025 3.23 27.255 3.23 27.255 3.62 29.265 3.62 29.265 3.23 29.495 3.23 29.495 3.62 31.505 3.62 31.505 3.23 31.735 3.23 31.735 3.62 33.6 3.62 33.745 3.62 33.745 2.53 33.975 2.53 33.975 3.62 34.72 3.62 34.72 4.22 33.6 4.22 21.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 34.72 -0.3 34.72 0.3 34.075 0.3 34.075 1.16 33.845 1.16 33.845 0.3 31.89 0.3 31.89 0.635 31.55 0.635 31.55 0.3 29.65 0.3 29.65 0.635 29.31 0.635 29.31 0.3 27.41 0.3 27.41 0.635 27.07 0.635 27.07 0.3 25.17 0.3 25.17 0.635 24.83 0.635 24.83 0.3 22.93 0.3 22.93 0.635 22.59 0.635 22.59 0.3 20.69 0.3 20.69 0.635 20.35 0.635 20.35 0.3 18.45 0.3 18.45 0.635 18.11 0.635 18.11 0.3 16.21 0.3 16.21 0.635 15.87 0.635 15.87 0.3 13.97 0.3 13.97 0.635 13.63 0.635 13.63 0.3 11.675 0.3 11.675 0.96 11.445 0.96 11.445 0.3 9.435 0.3 9.435 0.96 9.205 0.96 9.205 0.3 7.195 0.3 7.195 0.96 6.965 0.96 6.965 0.3 4.955 0.3 4.955 0.96 4.725 0.96 4.725 0.3 2.715 0.3 2.715 0.96 2.485 0.96 2.485 0.3 0.475 0.3 0.475 1.16 0.245 1.16 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.53 10.225 2.53 10.225 1.42 1.365 1.42 1.365 0.675 1.595 0.675 1.595 1.19 3.605 1.19 3.605 0.675 3.835 0.675 3.835 1.19 5.845 1.19 5.845 0.675 6.075 0.675 6.075 1.19 8.085 1.19 8.085 0.675 8.315 0.675 8.315 1.19 10.325 1.19 10.325 0.675 10.68 0.675 10.68 1.74 21.57 1.74 21.57 1.97 10.68 1.97 10.68 3.38 10.225 3.38 10.225 2.76 8.215 2.76 8.215 3.38 7.985 3.38 7.985 2.76 5.975 2.76 5.975 3.38 5.745 3.38 5.745 2.76 3.735 2.76 3.735 3.38 3.505 3.38 3.505 2.76 1.595 2.76 1.595 3.38 1.365 3.38  ;
        POLYGON 23.68 1.74 33.6 1.74 33.6 1.97 23.68 1.97  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_20

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.61 1.015 0.61 1.015 1.625 1.65 1.625 1.65 2.15 0.705 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.0804 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.675 2.21 4.175 2.21 4.58 2.21 4.58 1.3 2.675 1.3 2.675 0.57 2.905 0.57 2.905 1.065 4.58 1.065 4.58 0.57 5.16 0.57 5.16 3.39 4.58 3.39 4.58 2.66 4.175 2.66 2.905 2.66 2.905 3.39 2.675 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.21 3.62 1.21 2.91 1.55 2.91 1.55 3.62 3.64 3.62 3.64 2.91 3.98 2.91 3.98 3.62 4.175 3.62 5.6 3.62 5.6 4.22 4.175 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 4.08 0.3 4.08 0.765 3.74 0.765 3.74 0.3 1.84 0.3 1.84 0.765 1.5 0.765 1.5 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.57 0.475 0.57 0.475 2.39 1.9 2.39 1.9 1.55 4.175 1.55 4.175 1.89 2.13 1.89 2.13 2.625 0.475 2.625 0.475 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_3

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.84 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.1 1.06 1.1 1.06 1.715 2.15 1.715 2.15 2.15 0.62 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3656 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.605 2.36 4.095 2.36 4.36 2.36 4.36 1.42 3.605 1.42 3.605 0.675 3.865 0.675 3.865 1.14 5.845 1.14 5.845 0.675 6.075 0.675 6.075 1.42 5.16 1.42 5.16 2.36 5.975 2.36 5.975 3.38 5.745 3.38 5.745 2.68 4.095 2.68 3.835 2.68 3.835 3.38 3.605 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.57 0.475 2.57 0.475 3.62 2.385 3.62 2.385 3 2.615 3 2.615 3.62 4.095 3.62 4.625 3.62 4.625 3.05 4.855 3.05 4.855 3.62 6.81 3.62 6.865 3.62 6.865 2.57 7.095 2.57 7.095 3.62 7.84 3.62 7.84 4.22 6.81 4.22 4.095 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.84 -0.3 7.84 0.3 7.25 0.3 7.25 0.765 6.91 0.765 6.91 0.3 5.01 0.3 5.01 0.765 4.67 0.765 4.67 0.3 2.77 0.3 2.77 0.765 2.43 0.765 2.43 0.3 0.53 0.3 0.53 0.765 0.19 0.765 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 2.53 2.67 2.53 2.67 1.25 1.365 1.25 1.365 0.675 1.595 0.675 1.595 1.015 2.905 1.015 2.905 1.685 4.095 1.685 4.095 2.025 2.905 2.025 2.905 2.76 1.495 2.76 1.495 3.38 1.265 3.38  ;
        POLYGON 5.585 1.685 6.81 1.685 6.81 2.025 5.585 2.025  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__buf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__buf_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.715 3.51 1.715 3.51 2.15 0.65 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.7312 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.845 2.33 8.27 2.33 8.84 2.33 8.84 1.42 5.845 1.42 5.845 0.675 6.105 0.675 6.105 1.04 8.085 1.04 8.085 0.675 8.315 0.675 8.315 1.04 10.325 1.04 10.325 0.675 10.555 0.675 10.555 1.04 12.565 1.04 12.565 0.675 12.795 0.675 12.795 1.42 9.64 1.42 9.64 2.33 12.695 2.33 12.695 3.38 12.465 3.38 12.465 2.71 10.455 2.71 10.455 3.38 10.225 3.38 10.225 2.71 8.27 2.71 8.215 2.71 8.215 3.38 7.985 3.38 7.985 2.71 6.075 2.71 6.075 3.38 5.845 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.57 0.475 2.57 0.475 3.62 2.385 3.62 2.385 3.04 2.615 3.04 2.615 3.62 4.625 3.62 4.625 2.57 4.855 2.57 4.855 3.62 6.865 3.62 6.865 3.04 7.095 3.04 7.095 3.62 8.27 3.62 9.105 3.62 9.105 3.04 9.335 3.04 9.335 3.62 11.345 3.62 11.345 3.04 11.575 3.04 11.575 3.62 13.54 3.62 13.585 3.62 13.585 2.57 13.815 2.57 13.815 3.62 14.56 3.62 14.56 4.22 13.54 4.22 8.27 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 13.97 0.3 13.97 0.765 13.63 0.765 13.63 0.3 11.73 0.3 11.73 0.765 11.39 0.765 11.39 0.3 9.49 0.3 9.49 0.765 9.15 0.765 9.15 0.3 7.25 0.3 7.25 0.765 6.91 0.765 6.91 0.3 5.01 0.3 5.01 0.765 4.67 0.765 4.67 0.3 2.77 0.3 2.77 0.765 2.43 0.765 2.43 0.3 0.53 0.3 0.53 0.765 0.19 0.765 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 2.53 3.98 2.53 3.98 1.25 1.365 1.25 1.365 0.675 1.595 0.675 1.595 1.015 3.605 1.015 3.605 0.675 3.835 0.675 3.835 1.015 4.315 1.015 4.315 1.685 8.27 1.685 8.27 2.025 4.315 2.025 4.315 2.76 3.735 2.76 3.735 3.38 3.505 3.38 3.505 2.76 1.495 2.76 1.495 3.38 1.265 3.38  ;
        POLYGON 10.34 1.685 13.54 1.685 13.54 2.03 10.34 2.03  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__buf_8

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.84 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.052 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.36 1.78 2.36 1.78 1.65 2.19 1.65 2.19 2.68 0.87 2.68  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.526 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.795 6.33 1.795 6.33 2.12 4.6 2.12  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.77 2.92 6.855 2.92 6.95 2.92 7.18 2.92 7.18 1 6.77 1 6.77 0.6 7.71 0.6 7.71 3.38 6.95 3.38 6.855 3.38 6.77 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3.065 1.595 3.065 1.595 3.62 6.005 3.62 6.005 3.015 6.235 3.015 6.235 3.62 6.855 3.62 6.95 3.62 7.84 3.62 7.84 4.22 6.95 4.22 6.855 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.84 -0.3 7.84 0.3 6.455 0.3 6.455 0.79 6.225 0.79 6.225 0.3 1.65 0.3 1.65 0.76 1.31 0.76 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.005 2.86 1.005 2.86 2.48 3.175 2.48 3.175 2.74 2.63 2.74 2.63 1.24 0.575 1.24 0.575 3.37 0.19 3.37  ;
        POLYGON 2.29 3.16 4.14 3.16 4.14 1.22 3.76 1.22 3.76 0.99 4.37 0.99 4.37 3.16 4.92 3.16 4.92 2.36 6.625 2.36 6.625 1.88 6.855 1.88 6.855 2.59 5.235 2.59 5.235 3.39 2.29 3.39  ;
        POLYGON 2.34 0.53 5.115 0.53 5.115 1.335 6.95 1.335 6.95 1.565 4.885 1.565 4.885 0.76 3.32 0.76 3.32 1.88 3.91 1.88 3.91 2.93 3.65 2.93 3.65 2.17 3.09 2.17 3.09 0.76 2.34 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 25.76 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.77 1.59 1.77 1.59 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 6.477 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.125 1.77 11.48 1.77 11.48 2.15 5.125 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.2244 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.63 2.53 17.49 2.53 17.9 2.53 17.9 1.135 12.73 1.135 12.73 0.865 24.27 0.865 24.27 1.135 18.5 1.135 18.5 2.53 23.17 2.53 23.17 3.38 22.83 3.38 22.83 2.97 21.13 2.97 21.13 3.38 20.79 3.38 20.79 2.97 19.09 2.97 19.09 3.38 18.75 3.38 18.75 2.97 17.49 2.97 17.05 2.97 17.05 3.38 16.71 3.38 16.71 2.97 15.01 2.97 15.01 3.38 14.67 3.38 14.67 2.97 12.97 2.97 12.97 3.38 12.63 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.49 3.62 5.49 3.04 5.83 3.04 5.83 3.62 7.53 3.62 7.53 3.04 7.87 3.04 7.87 3.62 9.57 3.62 9.57 3.04 9.91 3.04 9.91 3.62 11.61 3.62 11.61 3.04 11.95 3.04 11.95 3.62 13.65 3.62 13.65 3.285 13.99 3.285 13.99 3.62 15.69 3.62 15.69 3.285 16.03 3.285 16.03 3.62 17.49 3.62 17.73 3.62 17.73 3.285 18.07 3.285 18.07 3.62 19.77 3.62 19.77 3.285 20.11 3.285 20.11 3.62 21.81 3.62 21.81 3.285 22.15 3.285 22.15 3.62 23.705 3.62 23.85 3.62 23.85 3.04 24.19 3.04 24.19 3.62 25.76 3.62 25.76 4.22 23.705 4.22 17.49 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 25.76 -0.3 25.76 0.3 25.39 0.3 25.39 0.635 25.05 0.635 25.05 0.3 23.15 0.3 23.15 0.635 22.81 0.635 22.81 0.3 20.91 0.3 20.91 0.635 20.57 0.635 20.57 0.3 18.67 0.3 18.67 0.635 18.33 0.635 18.33 0.3 16.43 0.3 16.43 0.635 16.09 0.635 16.09 0.3 14.19 0.3 14.19 0.635 13.85 0.635 13.85 0.3 11.95 0.3 11.95 0.635 11.61 0.635 11.61 0.3 9.71 0.3 9.71 0.635 9.37 0.635 9.37 0.3 7.47 0.3 7.47 0.635 7.13 0.635 7.13 0.3 5.01 0.3 5.01 0.475 4.67 0.475 4.67 0.3 1.65 0.3 1.65 0.655 1.31 0.655 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.78 1.905 2.78 1.905 1.325 0.19 1.325 0.19 0.85 0.53 0.85 0.53 1.095 2.135 1.095 2.135 2.235 3.65 2.235 3.65 2.52 2.135 2.52 2.135 3.01 0.42 3.01  ;
        POLYGON 2.485 0.53 4.44 0.53 4.44 0.705 5.945 0.705 5.945 0.865 12.01 0.865 12.01 1.365 16.875 1.365 16.875 1.595 11.78 1.595 11.78 1.095 5.695 1.095 5.695 0.935 4.215 0.935 4.215 0.76 2.715 0.76 2.715 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 2.485 2.005  ;
        POLYGON 2.685 3.16 4.595 3.16 4.595 1.545 3.77 1.545 3.77 1.14 4.11 1.14 4.11 1.315 4.825 1.315 4.825 2.53 11.78 2.53 11.78 1.965 17.49 1.965 17.49 2.195 12.01 2.195 12.01 2.76 10.93 2.76 10.93 3.38 10.59 3.38 10.59 2.76 8.89 2.76 8.89 3.38 8.55 3.38 8.55 2.76 6.85 2.76 6.85 3.38 6.51 3.38 6.51 2.76 4.825 2.76 4.825 3.39 2.685 3.39  ;
        POLYGON 19.01 1.365 23.705 1.365 23.705 1.595 19.01 1.595  ;
        POLYGON 19.33 1.965 23.705 1.965 23.705 2.195 19.33 2.195  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_12

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 32.48 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.77 1.59 1.77 1.59 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.5485 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.69 1.77 12.79 1.77 12.79 2.15 5.69 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.2992 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.95 2.505 21.92 2.505 22.23 2.505 22.23 1.095 14.97 1.095 14.97 0.865 30.99 0.865 30.99 1.095 23.13 1.095 23.13 2.505 29.57 2.505 29.57 3.38 29.23 3.38 29.23 3.055 27.53 3.055 27.53 3.38 27.19 3.38 27.19 3.055 25.49 3.055 25.49 3.38 25.15 3.38 25.15 3.055 23.45 3.055 23.45 3.38 23.13 3.38 23.13 3.055 21.92 3.055 21.41 3.055 21.41 3.38 21.07 3.38 21.07 3.055 19.37 3.055 19.37 3.38 19.03 3.38 19.03 3.055 17.33 3.055 17.33 3.38 16.99 3.38 16.99 3.055 15.29 3.055 15.29 3.38 14.95 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.29 3.62 5.29 3.04 5.63 3.04 5.63 3.62 7.33 3.62 7.33 3.04 7.67 3.04 7.67 3.62 9.37 3.62 9.37 3.04 9.71 3.04 9.71 3.62 11.71 3.62 11.71 3.04 12.05 3.04 12.05 3.62 13.93 3.62 13.93 2.53 14.27 2.53 14.27 3.62 15.97 3.62 15.97 3.285 16.31 3.285 16.31 3.62 18.01 3.62 18.01 3.285 18.35 3.285 18.35 3.62 20.05 3.62 20.05 3.285 20.39 3.285 20.39 3.62 21.92 3.62 22.09 3.62 22.09 3.285 22.43 3.285 22.43 3.62 24.13 3.62 24.13 3.285 24.47 3.285 24.47 3.62 26.17 3.62 26.17 3.285 26.51 3.285 26.51 3.62 28.21 3.62 28.21 3.285 28.55 3.285 28.55 3.62 30.08 3.62 30.305 3.62 30.305 2.53 30.535 2.53 30.535 3.62 31.52 3.62 32.48 3.62 32.48 4.22 31.52 4.22 30.08 4.22 21.92 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 32.48 -0.3 32.48 0.3 32.055 0.3 32.055 0.9 31.825 0.9 31.825 0.3 29.87 0.3 29.87 0.635 29.53 0.635 29.53 0.3 27.63 0.3 27.63 0.635 27.29 0.635 27.29 0.3 25.39 0.3 25.39 0.635 25.05 0.635 25.05 0.3 23.15 0.3 23.15 0.635 22.81 0.635 22.81 0.3 20.91 0.3 20.91 0.635 20.57 0.635 20.57 0.3 18.67 0.3 18.67 0.635 18.33 0.635 18.33 0.3 16.43 0.3 16.43 0.635 16.09 0.635 16.09 0.3 14.21 0.3 14.21 0.635 13.835 0.635 13.835 0.3 11.95 0.3 11.95 0.635 11.61 0.635 11.61 0.3 9.71 0.3 9.71 0.635 9.37 0.635 9.37 0.3 7.47 0.3 7.47 0.635 7.13 0.635 7.13 0.3 5.01 0.3 5.01 0.475 4.67 0.475 4.67 0.3 1.65 0.3 1.65 0.64 1.31 0.64 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.78 1.895 2.78 1.895 1.325 0.19 1.325 0.19 0.865 0.53 0.865 0.53 1.095 2.125 1.095 2.125 2.235 3.65 2.235 3.65 2.52 2.125 2.52 2.125 3.01 0.42 3.01  ;
        POLYGON 2.485 0.53 4.44 0.53 4.44 0.705 6.35 0.705 6.35 0.865 13.64 0.865 13.64 1.36 21.45 1.36 21.45 1.59 13.35 1.59 13.35 1.095 6.01 1.095 6.01 0.935 4.215 0.935 4.215 0.76 2.715 0.76 2.715 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 2.485 2.005  ;
        POLYGON 2.73 3.16 4.83 3.16 4.83 1.545 3.77 1.545 3.77 1.14 4.11 1.14 4.11 1.315 5.06 1.315 5.06 2.53 13.27 2.53 13.27 2 21.92 2 21.92 2.23 13.615 2.23 13.615 2.76 13.13 2.76 13.13 3.38 12.79 3.38 12.79 2.76 10.885 2.76 10.885 3.38 10.545 3.38 10.545 2.76 8.69 2.76 8.69 3.38 8.35 3.38 8.35 2.76 6.65 2.76 6.65 3.38 6.31 3.38 6.31 2.76 5.06 2.76 5.06 3.39 2.73 3.39  ;
        POLYGON 23.63 2 30.08 2 30.08 2.23 23.63 2.23  ;
        POLYGON 23.49 1.36 31.52 1.36 31.52 1.59 23.49 1.59  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_16

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.4 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 1.78 1.63 1.78 1.63 2.265 0.545 2.265  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0795 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.92 1.815 6.085 1.815 6.085 2.235 4.92 2.235  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0374 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.805 0.6 7.16 0.6 7.16 3.38 6.805 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.83 3.62 5.83 3.22 6.17 3.22 6.17 3.62 6.565 3.62 7.87 3.62 7.87 2.53 8.21 2.53 8.21 3.62 8.4 3.62 8.4 4.22 6.565 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.4 -0.3 8.4 0.3 8.155 0.3 8.155 0.9 7.925 0.9 7.925 0.3 5.915 0.3 5.915 0.9 5.685 0.9 5.685 0.3 1.65 0.3 1.65 0.64 1.31 0.64 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.78 1.9 2.78 1.9 1.325 0.19 1.325 0.19 0.865 0.53 0.865 0.53 1.095 2.13 1.095 2.13 2.235 3.65 2.235 3.65 2.52 2.13 2.52 2.13 3.01 0.42 3.01  ;
        POLYGON 2.485 0.53 5.355 0.53 5.355 1.355 6.51 1.355 6.51 1.585 5.125 1.585 5.125 0.76 2.715 0.76 2.715 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 2.485 2.005  ;
        POLYGON 2.7 3.16 4.46 3.16 4.46 1.545 3.77 1.545 3.77 0.99 4.11 0.99 4.11 1.315 4.69 1.315 4.69 2.7 6.335 2.7 6.335 1.9 6.565 1.9 6.565 2.93 5.175 2.93 5.175 3.39 2.7 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 11.2 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 1.775 1.63 1.775 1.63 2.185 0.545 2.185  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.658 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.09 1.8 7.275 1.8 7.275 2.12 5.09 2.12  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9152 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.46 2.54 10.37 2.54 10.49 2.54 10.74 2.54 10.74 1.135 8.34 1.135 8.34 0.865 11.07 0.865 11.07 2.77 10.84 2.77 10.84 3.39 10.5 3.39 10.5 2.77 10.49 2.77 10.37 2.77 8.8 2.77 8.8 3.39 8.46 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.22 3.62 5.22 3.285 5.56 3.285 5.56 3.62 7.26 3.62 7.26 3.285 7.6 3.285 7.6 3.62 9.48 3.62 9.48 3.285 9.82 3.285 9.82 3.62 10.37 3.62 10.49 3.62 11.2 3.62 11.2 4.22 10.49 4.22 10.37 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 11.2 -0.3 11.2 0.3 9.89 0.3 9.89 0.635 9.55 0.635 9.55 0.3 7.56 0.3 7.56 0.635 7.22 0.635 7.22 0.3 5.01 0.3 5.01 0.475 4.67 0.475 4.67 0.3 1.65 0.3 1.65 0.655 1.31 0.655 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.78 1.925 2.78 1.925 1.325 0.19 1.325 0.19 0.85 0.53 0.85 0.53 1.095 2.155 1.095 2.155 2.235 3.65 2.235 3.65 2.52 2.155 2.52 2.155 3.01 0.42 3.01  ;
        POLYGON 2.87 3.16 4.595 3.16 4.595 1.545 3.77 1.545 3.77 1.14 4.11 1.14 4.11 1.315 4.825 1.315 4.825 2.575 7.625 2.575 7.625 1.965 10.37 1.965 10.37 2.195 7.855 2.195 7.855 2.805 6.58 2.805 6.58 3.39 6.24 3.39 6.24 2.805 4.825 2.805 4.825 3.39 2.87 3.39  ;
        POLYGON 2.485 0.53 4.44 0.53 4.44 0.705 5.92 0.705 5.92 0.585 6.37 0.585 6.37 0.865 8.015 0.865 8.015 1.365 10.49 1.365 10.49 1.595 7.785 1.595 7.785 1.095 5.92 1.095 5.92 0.935 4.215 0.935 4.215 0.76 2.715 0.76 2.715 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 2.485 2.005  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_3

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.77 1.59 1.77 1.59 2.15 0.65 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.159 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.77 7.19 1.77 7.19 2.15 5.13 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.0748 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.35 2.52 10.15 2.52 10.73 2.52 10.73 1.135 8.16 1.135 8.16 0.865 11.11 0.865 11.11 2.76 10.73 2.76 10.73 3.38 10.39 3.38 10.39 2.8 10.15 2.8 8.69 2.8 8.69 3.38 8.35 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.29 3.62 5.29 3.285 5.63 3.285 5.63 3.62 7.33 3.62 7.33 3.285 7.67 3.285 7.67 3.62 9.37 3.62 9.37 3.285 9.71 3.285 9.71 3.62 10.15 3.62 11.41 3.62 11.41 3.285 11.75 3.285 11.75 3.62 12.32 3.62 12.32 4.22 10.15 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 11.95 0.3 11.95 0.635 11.61 0.635 11.61 0.3 9.71 0.3 9.71 0.635 9.37 0.635 9.37 0.3 7.47 0.3 7.47 0.635 7.13 0.635 7.13 0.3 5.01 0.3 5.01 0.475 4.67 0.475 4.67 0.3 1.65 0.3 1.65 0.655 1.31 0.655 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.78 1.925 2.78 1.925 1.325 0.19 1.325 0.19 0.85 0.53 0.85 0.53 1.095 2.155 1.095 2.155 2.235 3.65 2.235 3.65 2.52 2.155 2.52 2.155 3.01 0.42 3.01  ;
        POLYGON 2.485 0.53 4.44 0.53 4.44 0.705 5.945 0.705 5.945 0.865 7.745 0.865 7.745 1.365 10.15 1.365 10.15 1.595 7.515 1.595 7.515 1.095 5.695 1.095 5.695 0.935 4.215 0.935 4.215 0.76 2.715 0.76 2.715 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 2.485 2.005  ;
        POLYGON 2.87 3.16 4.595 3.16 4.595 1.545 3.77 1.545 3.77 1.14 4.11 1.14 4.11 1.315 4.825 1.315 4.825 2.53 7.515 2.53 7.515 1.965 10.15 1.965 10.15 2.195 7.745 2.195 7.745 2.76 6.65 2.76 6.65 3.38 6.31 3.38 6.31 2.76 4.825 2.76 4.825 3.39 2.87 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__bufz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__bufz_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.929 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 1.775 1.675 1.775 1.675 2.185 0.545 2.185  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.318 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.075 1.8 9.43 1.8 9.43 2.12 5.075 2.12  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.1496 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.39 2.425 12.26 2.425 12.52 2.425 13.42 2.425 13.42 1.135 10.4 1.135 10.4 0.865 17.55 0.865 17.55 1.135 14.07 1.135 14.07 2.425 16.85 2.425 16.85 3.38 16.51 3.38 16.51 2.765 14.81 2.765 14.81 3.38 14.47 3.38 14.47 2.765 12.77 2.765 12.77 3.38 12.52 3.38 12.43 3.38 12.43 2.765 12.26 2.765 10.73 2.765 10.73 3.38 10.39 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.45 3.62 1.45 3.26 1.79 3.26 1.79 3.62 5.29 3.62 5.29 3.285 5.63 3.285 5.63 3.62 7.33 3.62 7.33 3.285 7.67 3.285 7.67 3.62 9.37 3.62 9.37 3.285 9.71 3.285 9.71 3.62 11.41 3.62 11.41 3.285 11.75 3.285 11.75 3.62 12.26 3.62 12.52 3.62 13.45 3.62 13.45 3.285 13.79 3.285 13.79 3.62 15.49 3.62 15.49 3.285 15.83 3.285 15.83 3.62 17.43 3.62 17.53 3.62 17.53 3.285 17.87 3.285 17.87 3.62 17.99 3.62 19.04 3.62 19.04 4.22 17.99 4.22 17.43 4.22 12.52 4.22 12.26 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 18.67 0.3 18.67 0.635 18.33 0.635 18.33 0.3 16.43 0.3 16.43 0.635 16.09 0.635 16.09 0.3 14.19 0.3 14.19 0.635 13.85 0.635 13.85 0.3 11.95 0.3 11.95 0.635 11.61 0.635 11.61 0.3 9.71 0.3 9.71 0.635 9.37 0.635 9.37 0.3 7.47 0.3 7.47 0.635 7.13 0.635 7.13 0.3 5.01 0.3 5.01 0.475 4.67 0.475 4.67 0.3 1.65 0.3 1.65 0.655 1.31 0.655 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.42 2.78 1.925 2.78 1.925 1.325 0.19 1.325 0.19 0.85 0.53 0.85 0.53 1.095 2.155 1.095 2.155 2.235 3.65 2.235 3.65 2.52 2.155 2.52 2.155 3.01 0.42 3.01  ;
        POLYGON 2.68 3.16 4.595 3.16 4.595 1.545 3.77 1.545 3.77 1.14 4.11 1.14 4.11 1.315 4.825 1.315 4.825 2.53 9.755 2.53 9.755 1.965 12.26 1.965 12.26 2.195 9.985 2.195 9.985 2.76 8.635 2.76 8.635 3.38 8.405 3.38 8.405 2.76 6.595 2.76 6.595 3.38 6.365 3.38 6.365 2.76 4.825 2.76 4.825 3.39 2.68 3.39  ;
        POLYGON 2.39 0.53 4.44 0.53 4.44 0.705 5.945 0.705 5.945 0.865 9.985 0.865 9.985 1.365 12.52 1.365 12.52 1.595 9.755 1.595 9.755 1.095 5.695 1.095 5.695 0.935 4.215 0.935 4.215 0.76 3.435 0.76 3.435 1.775 4.23 1.775 4.23 2.93 3.89 2.93 3.89 2.005 3.205 2.005 3.205 0.76 2.39 0.76  ;
        POLYGON 15.05 1.965 17.43 1.965 17.43 2.195 15.05 2.195  ;
        POLYGON 15.415 1.365 17.99 1.365 17.99 1.595 15.415 1.595  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__bufz_8

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 3.36 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.741 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.035 1.08 1.035 1.08 1.74 1.59 1.74 1.59 2.15 0.705 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.7546 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.34 0.565 2.93 0.565 2.93 3.32 2.565 3.32 2.565 1.605 2.34 1.605  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 3.015 1.65 3.015 1.65 3.62 2.27 3.62 3.36 3.62 3.36 4.22 2.27 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 3.36 -0.3 3.36 0.3 1.65 0.3 1.65 0.925 1.31 0.925 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.565 0.475 0.565 0.475 2.52 1.93 2.52 1.93 1.88 2.27 1.88 2.27 2.755 0.575 2.755 0.575 3.38 0.245 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.555 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.765 6.07 1.765 6.07 2.15 0.62 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.036 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.265 2.495 13.09 2.495 13.83 2.495 13.83 1.535 8.265 1.535 8.265 0.69 8.495 0.69 8.495 1.215 10.505 1.215 10.505 0.69 10.735 0.69 10.735 1.215 12.745 1.215 12.745 0.69 12.975 0.69 12.975 1.215 14.985 1.215 14.985 0.69 15.215 0.69 15.215 1.215 17.225 1.215 17.225 0.69 17.455 0.69 17.455 1.215 19.465 1.215 19.465 0.69 19.695 0.69 19.695 1.535 14.73 1.535 14.73 2.495 19.595 2.495 19.595 3.39 19.365 3.39 19.365 3 17.355 3 17.355 3.39 17.125 3.39 17.125 3 15.115 3 15.115 3.39 14.885 3.39 14.885 3 13.09 3 12.875 3 12.875 3.39 12.645 3.39 12.645 3 10.635 3 10.635 3.39 10.405 3.39 10.405 3 8.495 3 8.495 3.39 8.265 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.23 0.475 3.23 0.475 3.62 2.385 3.62 2.385 3.05 2.615 3.05 2.615 3.62 4.625 3.62 4.625 3.05 4.855 3.05 4.855 3.62 7.145 3.62 7.145 3.23 7.375 3.23 7.375 3.62 9.285 3.62 9.285 3.23 9.515 3.23 9.515 3.62 11.525 3.62 11.525 3.23 11.755 3.23 11.755 3.62 13.09 3.62 13.765 3.62 13.765 3.23 13.995 3.23 13.995 3.62 16.005 3.62 16.005 3.23 16.235 3.23 16.235 3.62 18.245 3.62 18.245 3.23 18.475 3.23 18.475 3.62 20.43 3.62 20.485 3.62 20.485 2.76 20.715 2.76 20.715 3.62 21.28 3.62 21.28 4.22 20.43 4.22 13.09 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 20.87 0.3 20.87 0.985 20.53 0.985 20.53 0.3 18.63 0.3 18.63 0.985 18.29 0.985 18.29 0.3 16.39 0.3 16.39 0.985 16.05 0.985 16.05 0.3 14.15 0.3 14.15 0.985 13.81 0.985 13.81 0.3 11.91 0.3 11.91 0.985 11.57 0.985 11.57 0.3 9.67 0.3 9.67 0.985 9.33 0.985 9.33 0.3 7.43 0.3 7.43 1.075 7.09 1.075 7.09 0.3 5.01 0.3 5.01 1.075 4.67 1.075 4.67 0.3 2.77 0.3 2.77 1.075 2.43 1.075 2.43 0.3 0.53 0.3 0.53 1.075 0.19 1.075 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 2.53 6.365 2.53 6.365 1.535 1.31 1.535 1.31 0.845 1.65 0.845 1.65 1.305 3.55 1.305 3.55 0.845 3.89 0.845 3.89 1.305 5.79 1.305 5.79 0.845 6.13 0.845 6.13 1.305 6.595 1.305 6.595 1.765 13.09 1.765 13.09 2.065 6.595 2.065 6.595 2.76 5.975 2.76 5.975 3.39 5.745 3.39 5.745 2.76 3.735 2.76 3.735 3.39 3.505 3.39 3.505 2.76 1.495 2.76 1.495 3.39 1.265 3.39  ;
        POLYGON 15.39 1.765 20.43 1.765 20.43 2.065 15.39 2.065  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_12

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 28 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.738 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.74 8.31 1.74 8.31 2.15 0.37 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.0688 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.505 2.42 17.16 2.42 17.985 2.42 17.985 1.535 10.505 1.535 10.505 0.69 10.735 0.69 10.735 1.215 12.745 1.215 12.745 0.69 12.975 0.69 12.975 1.215 14.985 1.215 14.985 0.69 15.215 0.69 15.215 1.215 17.225 1.215 17.225 0.69 17.455 0.69 17.455 1.215 19.465 1.215 19.465 0.69 19.695 0.69 19.695 1.215 21.705 1.215 21.705 0.69 21.935 0.69 21.935 1.215 23.945 1.215 23.945 0.69 24.175 0.69 24.175 1.215 26.185 1.215 26.185 0.69 26.415 0.69 26.415 1.535 18.885 1.535 18.885 2.42 26.315 2.42 26.315 3.39 26.085 3.39 26.085 3 24.075 3 24.075 3.39 23.845 3.39 23.845 3 21.835 3 21.835 3.39 21.605 3.39 21.605 3 19.595 3 19.595 3.39 19.365 3.39 19.365 3 17.355 3 17.355 3.39 17.16 3.39 17.125 3.39 17.125 3 15.115 3 15.115 3.39 14.885 3.39 14.885 3 12.875 3 12.875 3.39 12.645 3.39 12.645 3 10.735 3 10.735 3.39 10.505 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.23 0.475 3.23 0.475 3.62 2.385 3.62 2.385 3.05 2.615 3.05 2.615 3.62 4.625 3.62 4.625 3.05 4.855 3.05 4.855 3.62 6.865 3.62 6.865 3.05 7.095 3.05 7.095 3.62 9.385 3.62 9.385 3.19 9.615 3.19 9.615 3.62 11.525 3.62 11.525 3.23 11.755 3.23 11.755 3.62 13.765 3.62 13.765 3.23 13.995 3.23 13.995 3.62 16.005 3.62 16.005 3.23 16.235 3.23 16.235 3.62 17.16 3.62 18.245 3.62 18.245 3.23 18.475 3.23 18.475 3.62 20.485 3.62 20.485 3.23 20.715 3.23 20.715 3.62 22.725 3.62 22.725 3.23 22.955 3.23 22.955 3.62 24.965 3.62 24.965 3.23 25.195 3.23 25.195 3.62 27.16 3.62 27.205 3.62 27.205 2.76 27.435 2.76 27.435 3.62 28 3.62 28 4.22 27.16 4.22 17.16 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 28 -0.3 28 0.3 27.59 0.3 27.59 0.985 27.25 0.985 27.25 0.3 25.35 0.3 25.35 0.985 25.01 0.985 25.01 0.3 23.11 0.3 23.11 0.985 22.77 0.985 22.77 0.3 20.87 0.3 20.87 0.985 20.53 0.985 20.53 0.3 18.63 0.3 18.63 0.985 18.29 0.985 18.29 0.3 16.39 0.3 16.39 0.985 16.05 0.985 16.05 0.3 14.15 0.3 14.15 0.985 13.81 0.985 13.81 0.3 11.91 0.3 11.91 0.985 11.57 0.985 11.57 0.3 9.67 0.3 9.67 0.96 9.33 0.96 9.33 0.3 7.25 0.3 7.25 1.04 6.91 1.04 6.91 0.3 5.01 0.3 5.01 1.04 4.67 1.04 4.67 0.3 2.77 0.3 2.77 1.04 2.43 1.04 2.43 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 2.53 8.62 2.53 8.62 1.5 1.365 1.5 1.365 0.74 1.595 0.74 1.595 1.27 3.605 1.27 3.605 0.74 3.835 0.74 3.835 1.27 5.845 1.27 5.845 0.74 6.075 0.74 6.075 1.27 8.085 1.27 8.085 0.74 8.315 0.74 8.315 1.27 8.85 1.27 8.85 1.765 17.16 1.765 17.16 2.065 8.85 2.065 8.85 2.76 8.215 2.76 8.215 3.39 7.985 3.39 7.985 2.76 5.975 2.76 5.975 3.39 5.745 3.39 5.745 2.76 3.735 2.76 3.735 3.39 3.505 3.39 3.505 2.76 1.495 2.76 1.495 3.39 1.265 3.39  ;
        POLYGON 19.74 1.765 27.16 1.765 27.16 2.065 19.74 2.065  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_16

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.726 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.55 1.08 0.55 1.08 1.74 1.65 1.74 1.65 2.15 0.705 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0086 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.665 2.36 3.21 2.36 3.47 2.36 3.47 1.51 2.665 1.51 2.665 0.8 2.895 0.8 2.895 1.28 3.81 1.28 3.81 2.71 3.21 2.71 2.895 2.71 2.895 3.39 2.665 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.36 3.62 1.36 3.05 1.7 3.05 1.7 3.62 3.21 3.62 3.685 3.62 3.685 3.05 3.915 3.05 3.915 3.62 4.48 3.62 4.48 4.22 3.21 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 4.07 0.3 4.07 1.05 3.73 1.05 3.73 0.3 1.83 0.3 1.83 1.095 1.49 1.095 1.49 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.805 0.475 0.805 0.475 2.59 1.89 2.59 1.89 1.74 3.21 1.74 3.21 2.04 2.215 2.04 2.215 2.82 0.475 2.82 0.475 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 34.72 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 5.924 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.74 9.9 1.74 9.9 2.12 0.63 2.12  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.13 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.13 2.27 32.66 2.27 33.135 2.27 33.135 3.39 32.905 3.39 32.905 3 32.66 3 30.795 3 30.795 3.39 30.565 3.39 30.565 3 28.555 3 28.555 3.39 28.325 3.39 28.325 3 26.315 3 26.315 3.39 26.085 3.39 26.085 3 24.075 3 24.075 3.39 23.845 3.39 23.845 3 21.835 3 21.835 3.39 21.605 3.39 21.605 3 21.28 3 19.595 3 19.595 3.39 19.365 3.39 19.365 3 17.355 3 17.355 3.39 17.125 3.39 17.125 3 15.115 3 15.115 3.39 14.885 3.39 14.885 3 12.975 3 12.975 3.39 12.745 3.39 12.745 2.27 21.28 2.27 22.23 2.27 22.23 1.535 12.745 1.535 12.745 0.685 13.005 0.685 13.005 1.215 14.985 1.215 14.985 0.685 15.215 0.685 15.215 1.215 17.225 1.215 17.225 0.685 17.455 0.685 17.455 1.215 19.465 1.215 19.465 0.685 19.695 0.685 19.695 1.215 21.705 1.215 21.705 0.685 21.935 0.685 21.935 1.215 23.945 1.215 23.945 0.685 24.175 0.685 24.175 1.215 26.185 1.215 26.185 0.685 26.415 0.685 26.415 1.215 28.425 1.215 28.425 0.685 28.655 0.685 28.655 1.215 30.665 1.215 30.665 0.685 30.895 0.685 30.895 1.215 32.905 1.215 32.905 0.685 33.135 0.685 33.135 1.535 23.13 1.535  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.23 0.475 3.23 0.475 3.62 2.385 3.62 2.385 3.05 2.615 3.05 2.615 3.62 4.625 3.62 4.625 3.05 4.855 3.05 4.855 3.62 6.865 3.62 6.865 3.05 7.095 3.05 7.095 3.62 9.105 3.62 9.105 3.05 9.335 3.05 9.335 3.62 11.625 3.62 11.625 3.23 11.855 3.23 11.855 3.62 13.765 3.62 13.765 3.23 13.995 3.23 13.995 3.62 16.005 3.62 16.005 3.23 16.235 3.23 16.235 3.62 18.245 3.62 18.245 3.23 18.475 3.23 18.475 3.62 20.485 3.62 20.485 3.23 20.715 3.23 20.715 3.62 21.28 3.62 22.725 3.62 22.725 3.23 22.955 3.23 22.955 3.62 24.965 3.62 24.965 3.23 25.195 3.23 25.195 3.62 27.205 3.62 27.205 3.23 27.435 3.23 27.435 3.62 29.445 3.62 29.445 3.23 29.675 3.23 29.675 3.62 31.685 3.62 31.685 3.23 31.915 3.23 31.915 3.62 32.66 3.62 34.025 3.62 34.025 2.71 34.255 2.71 34.255 3.62 34.72 3.62 34.72 4.22 32.66 4.22 21.28 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 34.72 -0.3 34.72 0.3 34.255 0.3 34.255 1.05 34.025 1.05 34.025 0.3 32.07 0.3 32.07 0.985 31.73 0.985 31.73 0.3 29.83 0.3 29.83 0.985 29.49 0.985 29.49 0.3 27.59 0.3 27.59 0.985 27.25 0.985 27.25 0.3 25.35 0.3 25.35 0.985 25.01 0.985 25.01 0.3 23.11 0.3 23.11 0.985 22.77 0.985 22.77 0.3 20.87 0.3 20.87 0.985 20.53 0.985 20.53 0.3 18.63 0.3 18.63 0.985 18.29 0.985 18.29 0.3 16.39 0.3 16.39 0.985 16.05 0.985 16.05 0.3 14.15 0.3 14.15 0.985 13.81 0.985 13.81 0.3 11.675 0.3 11.675 1.04 11.445 1.04 11.445 0.3 9.435 0.3 9.435 1.04 9.205 1.04 9.205 0.3 7.195 0.3 7.195 1.04 6.965 1.04 6.965 0.3 4.955 0.3 4.955 1.04 4.725 1.04 4.725 0.3 2.715 0.3 2.715 1.04 2.485 1.04 2.485 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.53 10.325 2.53 10.325 1.505 1.365 1.505 1.365 0.685 1.595 0.685 1.595 1.27 3.605 1.27 3.605 0.685 3.835 0.685 3.835 1.27 5.845 1.27 5.845 0.685 6.075 0.685 6.075 1.27 8.085 1.27 8.085 0.685 8.315 0.685 8.315 1.27 10.325 1.27 10.325 0.685 10.555 0.685 10.555 1.765 21.28 1.765 21.28 1.995 10.555 1.995 10.555 3.39 10.325 3.39 10.325 2.82 8.215 2.82 8.215 3.39 7.985 3.39 7.985 2.76 5.975 2.76 5.975 3.39 5.745 3.39 5.745 2.76 3.735 2.76 3.735 3.39 3.505 3.39 3.505 2.76 1.595 2.76 1.595 3.39 1.365 3.39  ;
        POLYGON 23.86 1.765 32.66 1.765 32.66 1.995 23.86 1.995  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_20

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.84 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.183 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.74 2.34 1.74 2.34 2.12 0.62 2.12  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.986 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.785 2.36 5.945 2.36 6.28 2.36 6.28 1.51 3.785 1.51 3.785 0.69 4.015 0.69 4.015 1.28 6.025 1.28 6.025 0.69 6.255 0.69 6.255 1.28 6.6 1.28 6.6 2.68 6.155 2.68 6.155 3.39 5.945 3.39 5.925 3.39 5.925 2.68 4.015 2.68 4.015 3.39 3.785 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.2 0.475 3.2 0.475 3.62 2.385 3.62 2.385 3.16 2.615 3.16 2.615 3.62 4.805 3.62 4.805 3.05 5.035 3.05 5.035 3.62 5.945 3.62 7.045 3.62 7.045 2.73 7.275 2.73 7.275 3.62 7.84 3.62 7.84 4.22 5.945 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.84 -0.3 7.84 0.3 7.43 0.3 7.43 0.985 7.09 0.985 7.09 0.3 5.19 0.3 5.19 0.985 4.85 0.985 4.85 0.3 2.95 0.3 2.95 0.985 2.61 0.985 2.61 0.3 0.53 0.3 0.53 0.985 0.19 0.985 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 2.59 2.955 2.59 2.955 1.5 1.365 1.5 1.365 0.69 1.595 0.69 1.595 1.27 3.185 1.27 3.185 1.74 5.945 1.74 5.945 2.04 3.185 2.04 3.185 2.82 1.495 2.82 1.495 3.39 1.265 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_3

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.84 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.183 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.74 2.15 1.74 2.15 2.15 0.37 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.986 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.785 2.36 4.83 2.36 5.13 2.36 5.13 1.445 3.785 1.445 3.785 0.69 4.015 0.69 4.015 1.215 6.025 1.215 6.025 0.69 6.255 0.69 6.255 1.445 5.51 1.445 5.51 2.36 6.155 2.36 6.155 3.39 5.925 3.39 5.925 2.68 4.83 2.68 4.015 2.68 4.015 3.39 3.785 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.23 0.475 3.23 0.475 3.62 2.385 3.62 2.385 3.16 2.615 3.16 2.615 3.62 4.805 3.62 4.805 3.05 4.83 3.05 5.035 3.05 5.035 3.62 6.935 3.62 7.045 3.62 7.045 2.76 7.275 2.76 7.275 3.62 7.84 3.62 7.84 4.22 6.935 4.22 4.83 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.84 -0.3 7.84 0.3 7.43 0.3 7.43 0.985 7.09 0.985 7.09 0.3 5.19 0.3 5.19 0.985 4.85 0.985 4.85 0.3 2.95 0.3 2.95 0.985 2.61 0.985 2.61 0.3 0.53 0.3 0.53 1.04 0.19 1.04 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.265 2.53 2.945 2.53 2.945 1.5 1.365 1.5 1.365 0.74 1.595 0.74 1.595 1.27 3.175 1.27 3.175 1.685 4.83 1.685 4.83 2.025 3.175 2.025 3.175 2.76 1.495 2.76 1.495 3.38 1.265 3.38  ;
        POLYGON 5.765 1.685 6.935 1.685 6.935 2.025 5.765 2.025  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.369 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.745 4.13 1.745 4.13 2.15 0.65 2.15  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.99 2.36 12.975 2.36 12.975 3.39 12.745 3.39 12.745 2.68 10.735 2.68 10.735 3.39 10.505 3.39 10.505 2.68 8.92 2.68 8.495 2.68 8.495 3.39 8.265 3.39 8.265 2.68 6.255 2.68 6.255 3.39 6.025 3.39 6.025 2.36 8.92 2.36 9.61 2.36 9.61 1.51 6.025 1.51 6.025 0.69 6.255 0.69 6.255 1.22 8.265 1.22 8.265 0.69 8.495 0.69 8.495 1.22 10.505 1.22 10.505 0.69 10.735 0.69 10.735 1.22 12.745 1.22 12.745 0.69 12.975 0.69 12.975 1.51 9.99 1.51  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 3.23 0.475 3.23 0.475 3.62 2.485 3.62 2.485 3.05 2.715 3.05 2.715 3.62 4.905 3.62 4.905 3.23 5.135 3.23 5.135 3.62 7.145 3.62 7.145 3.05 7.375 3.05 7.375 3.62 8.92 3.62 9.385 3.62 9.385 3.05 9.615 3.05 9.615 3.62 11.625 3.62 11.625 3.05 11.855 3.05 11.855 3.62 13.72 3.62 13.865 3.62 13.865 2.76 14.095 2.76 14.095 3.62 14.56 3.62 14.56 4.22 13.72 4.22 8.92 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 14.15 0.3 14.15 0.985 13.81 0.985 13.81 0.3 11.91 0.3 11.91 0.985 11.57 0.985 11.57 0.3 9.67 0.3 9.67 0.985 9.33 0.985 9.33 0.3 7.43 0.3 7.43 0.985 7.09 0.985 7.09 0.3 5.19 0.3 5.19 1.055 4.85 1.055 4.85 0.3 2.77 0.3 2.77 1.04 2.43 1.04 2.43 0.3 0.53 0.3 0.53 1.04 0.19 1.04 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 2.53 4.425 2.53 4.425 1.5 1.365 1.5 1.365 0.74 1.595 0.74 1.595 1.27 3.605 1.27 3.605 0.74 3.835 0.74 3.835 1.27 4.655 1.27 4.655 1.74 8.92 1.74 8.92 1.975 4.655 1.975 4.655 2.76 3.835 2.76 3.835 3.39 3.605 3.39 3.605 2.76 1.595 2.76 1.595 3.39 1.365 3.39  ;
        POLYGON 10.53 1.74 13.72 1.74 13.72 2.04 10.53 2.04  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__clkbuf_8

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 2.24 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.898 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.97 1.03 0.97 1.03 2.95 0.705 2.95  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.748 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.26 0.6 1.595 0.6 1.595 3.37 1.26 3.37  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.48 0.475 2.48 0.475 3.62 2.24 3.62 2.24 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 2.24 -0.3 2.24 0.3 0.475 0.3 0.475 1.04 0.245 1.04 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 10.776 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.765 5.82 1.765 5.82 2.15 0.62 2.15  ;
        POLYGON 7.99 1.765 13.54 1.765 13.54 2.15 7.99 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.036 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.57 6.55 2.57 6.55 1.535 1.365 1.535 1.365 0.585 1.595 0.585 1.595 1.1 3.605 1.1 3.605 0.585 3.835 0.585 3.835 1.1 5.845 1.1 5.845 0.585 6.075 0.585 6.075 1.1 8.085 1.1 8.085 0.585 8.315 0.585 8.315 1.1 10.325 1.1 10.325 0.585 10.555 0.585 10.555 1.1 12.565 1.1 12.565 0.585 12.795 0.585 12.795 1.535 7.45 1.535 7.45 2.57 12.695 2.57 12.695 3.38 12.465 3.38 12.465 3.045 10.455 3.045 10.455 3.38 10.225 3.38 10.225 3.045 8.215 3.045 8.215 3.38 7.985 3.38 7.985 3.045 6.07 3.045 6.07 3.38 5.69 3.38 5.69 3.05 3.735 3.05 3.735 3.38 3.505 3.38 3.505 3.05 1.495 3.05 1.495 3.38 1.265 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.57 0.475 2.57 0.475 3.62 2.33 3.62 2.33 3.28 2.67 3.28 2.67 3.62 4.57 3.62 4.57 3.28 4.91 3.28 4.91 3.62 6.81 3.62 6.81 3.28 7.15 3.28 7.15 3.62 9.05 3.62 9.05 3.28 9.39 3.28 9.39 3.62 11.29 3.62 11.29 3.28 11.63 3.28 11.63 3.62 13.585 3.62 13.585 2.57 13.815 2.57 13.815 3.62 14.56 3.62 14.56 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 13.915 0.3 13.915 0.925 13.685 0.925 13.685 0.3 11.73 0.3 11.73 0.87 11.39 0.87 11.39 0.3 9.49 0.3 9.49 0.87 9.15 0.87 9.15 0.3 7.25 0.3 7.25 0.87 6.91 0.87 6.91 0.3 5.01 0.3 5.01 0.87 4.67 0.87 4.67 0.3 2.77 0.3 2.77 0.87 2.43 0.87 2.43 0.3 0.475 0.3 0.475 0.925 0.245 0.925 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_12

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 14.368 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.64 1.76 8.13 1.76 8.13 2.15 0.64 2.15  ;
        POLYGON 10.28 1.765 17.67 1.765 17.67 2.15 10.28 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 8.048 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.475 8.79 2.475 8.79 1.455 1.31 1.455 1.31 0.53 1.65 0.53 1.65 0.875 3.55 0.875 3.55 0.53 3.89 0.53 3.89 0.875 5.79 0.875 5.79 0.53 6.13 0.53 6.13 0.875 8.03 0.875 8.03 0.53 8.37 0.53 8.37 0.875 10.27 0.875 10.27 0.53 10.61 0.53 10.61 0.875 12.51 0.875 12.51 0.53 12.85 0.53 12.85 0.875 14.75 0.875 14.75 0.53 15.09 0.53 15.09 0.875 16.99 0.875 16.99 0.53 17.33 0.53 17.33 1.455 9.69 1.455 9.69 2.475 17.175 2.475 17.175 3.38 16.945 3.38 16.945 3.055 14.935 3.055 14.935 3.38 14.705 3.38 14.705 3.055 12.695 3.055 12.695 3.38 12.465 3.38 12.465 3.055 10.455 3.055 10.455 3.38 10.225 3.38 10.225 3.055 8.31 3.055 8.31 3.38 7.93 3.38 7.93 3.055 5.975 3.055 5.975 3.38 5.745 3.38 5.745 3.055 3.735 3.055 3.735 3.38 3.505 3.38 3.505 3.055 1.495 3.055 1.495 3.38 1.265 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.57 0.475 2.57 0.475 3.62 2.33 3.62 2.33 3.285 2.67 3.285 2.67 3.62 4.57 3.62 4.57 3.285 4.91 3.285 4.91 3.62 6.81 3.62 6.81 3.285 7.15 3.285 7.15 3.62 9.05 3.62 9.05 3.285 9.39 3.285 9.39 3.62 11.29 3.62 11.29 3.285 11.63 3.285 11.63 3.62 13.53 3.62 13.53 3.285 13.87 3.285 13.87 3.62 15.77 3.62 15.77 3.285 16.11 3.285 16.11 3.62 18.065 3.62 18.065 2.53 18.295 2.53 18.295 3.62 19.04 3.62 19.04 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 18.395 0.3 18.395 0.7 18.165 0.7 18.165 0.3 16.21 0.3 16.21 0.645 15.87 0.645 15.87 0.3 13.97 0.3 13.97 0.645 13.63 0.645 13.63 0.3 11.73 0.3 11.73 0.645 11.39 0.645 11.39 0.3 9.49 0.3 9.49 0.645 9.15 0.645 9.15 0.3 7.25 0.3 7.25 0.645 6.91 0.645 6.91 0.3 5.01 0.3 5.01 0.645 4.67 0.645 4.67 0.3 2.77 0.3 2.77 0.645 2.43 0.645 2.43 0.3 0.475 0.3 0.475 0.7 0.245 0.7 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_16

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 3.36 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.796 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.19 1.035 1.19 1.035 1.735 1.97 1.735 1.97 2.12 1.035 2.12 1.035 2.875 0.705 2.875  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.006 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.36 2.33 2.36 2.33 1.505 1.365 1.505 1.365 0.68 1.595 0.68 1.595 1.27 2.71 1.27 2.71 2.735 1.495 2.735 1.495 3.38 1.265 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.33 3.62 2.33 2.965 2.67 2.965 2.67 3.62 3.36 3.62 3.36 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 3.36 -0.3 3.36 0.3 2.715 0.3 2.715 1.04 2.485 1.04 2.485 0.3 0.475 0.3 0.475 1.04 0.245 1.04 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 23.52 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 17.96 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.74 9.9 1.74 9.9 2.12 0.63 2.12  ;
        POLYGON 12.52 1.74 22.4 1.74 22.4 2.12 12.52 2.12  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 10.06 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.35 11.03 2.35 11.03 1.505 1.31 1.505 1.31 0.535 1.65 0.535 1.65 0.875 3.55 0.875 3.55 0.535 3.89 0.535 3.89 0.875 5.79 0.875 5.79 0.535 6.13 0.535 6.13 0.875 8.03 0.875 8.03 0.535 8.37 0.535 8.37 0.875 10.27 0.875 10.27 0.535 10.61 0.535 10.61 0.875 12.51 0.875 12.51 0.535 12.85 0.535 12.85 0.875 14.75 0.875 14.75 0.535 15.09 0.535 15.09 0.875 16.99 0.875 16.99 0.535 17.33 0.535 17.33 0.875 19.23 0.875 19.23 0.535 19.57 0.535 19.57 0.875 21.47 0.875 21.47 0.535 21.81 0.535 21.81 1.505 11.93 1.505 11.93 2.35 21.655 2.35 21.655 3.38 21.425 3.38 21.425 3.055 19.415 3.055 19.415 3.38 19.185 3.38 19.185 3.055 17.175 3.055 17.175 3.38 16.945 3.38 16.945 3.055 14.935 3.055 14.935 3.38 14.705 3.38 14.705 3.055 12.695 3.055 12.695 3.38 12.465 3.38 12.465 3.055 10.55 3.055 10.55 3.38 10.17 3.38 10.17 3.055 8.215 3.055 8.215 3.38 7.985 3.38 7.985 3.055 5.975 3.055 5.975 3.38 5.745 3.38 5.745 3.055 3.735 3.055 3.735 3.38 3.505 3.38 3.505 3.055 1.595 3.055 1.595 3.38 1.365 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.33 3.62 2.33 3.285 2.67 3.285 2.67 3.62 4.57 3.62 4.57 3.285 4.91 3.285 4.91 3.62 6.81 3.62 6.81 3.285 7.15 3.285 7.15 3.62 9.05 3.62 9.05 3.285 9.39 3.285 9.39 3.62 11.29 3.62 11.29 3.285 11.63 3.285 11.63 3.62 13.53 3.62 13.53 3.285 13.87 3.285 13.87 3.62 15.77 3.62 15.77 3.285 16.11 3.285 16.11 3.62 18.01 3.62 18.01 3.285 18.35 3.285 18.35 3.62 20.25 3.62 20.25 3.285 20.59 3.285 20.59 3.62 22.545 3.62 22.545 2.53 22.775 2.53 22.775 3.62 23.52 3.62 23.52 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 23.52 -0.3 23.52 0.3 22.93 0.3 22.93 0.645 22.59 0.645 22.59 0.3 20.69 0.3 20.69 0.645 20.35 0.645 20.35 0.3 18.45 0.3 18.45 0.645 18.11 0.645 18.11 0.3 16.21 0.3 16.21 0.645 15.87 0.645 15.87 0.3 13.97 0.3 13.97 0.645 13.63 0.645 13.63 0.3 11.73 0.3 11.73 0.645 11.39 0.645 11.39 0.3 9.49 0.3 9.49 0.645 9.15 0.645 9.15 0.3 7.25 0.3 7.25 0.645 6.91 0.645 6.91 0.3 5.01 0.3 5.01 0.645 4.67 0.645 4.67 0.3 2.77 0.3 2.77 0.645 2.43 0.645 2.43 0.3 0.475 0.3 0.475 0.7 0.245 0.7 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_20

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.694 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.74 2.855 1.74 2.855 2.12 0.65 2.12  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.754 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.36 3.46 2.36 3.46 1.505 1.365 1.505 1.365 0.7 1.595 0.7 1.595 1.27 3.45 1.27 3.45 0.65 3.835 0.65 3.835 3.38 3.45 3.38 3.45 2.735 1.495 2.735 1.495 3.38 1.265 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.55 0.475 2.55 0.475 3.62 2.33 3.62 2.33 2.965 2.67 2.965 2.67 3.62 4.48 3.62 4.48 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 2.715 0.3 2.715 1.04 2.485 1.04 2.485 0.3 0.475 0.3 0.475 1.04 0.245 1.04 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_3

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.592 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.765 2.71 1.765 2.71 2.15 0.65 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.256 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.385 3.45 2.385 3.45 1.535 1.365 1.535 1.365 0.7 1.595 0.7 1.595 1.215 3.45 1.215 3.45 0.7 3.835 0.7 3.835 3.27 3.45 3.27 3.45 2.705 1.595 2.705 1.595 3.27 1.365 3.27  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.59 0.475 2.59 0.475 3.62 2.43 3.62 2.43 2.965 2.77 2.965 2.77 3.62 4.725 3.62 4.725 2.59 4.955 2.59 4.955 3.62 5.6 3.62 5.6 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 4.955 0.3 4.955 1.04 4.725 1.04 4.725 0.3 2.77 0.3 2.77 0.985 2.43 0.985 2.43 0.3 0.475 0.3 0.475 1.04 0.245 1.04 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__clkinv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__clkinv_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 7.184 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.765 3.79 1.765 3.79 2.15 0.63 2.15  ;
        POLYGON 5.33 1.765 8.96 1.765 8.96 2.15 5.33 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.024 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.41 4.57 2.41 4.57 1.535 1.365 1.535 1.365 0.7 1.595 0.7 1.595 1.215 3.605 1.215 3.605 0.7 3.835 0.7 3.835 1.215 5.845 1.215 5.845 0.7 6.075 0.7 6.075 1.215 8.085 1.215 8.085 0.7 8.315 0.7 8.315 1.535 4.95 1.535 4.95 2.41 8.215 2.41 8.215 3.38 7.985 3.38 7.985 2.725 5.975 2.725 5.975 3.38 5.745 3.38 5.745 2.725 3.735 2.725 3.735 3.38 3.505 3.38 3.505 2.73 1.495 2.73 1.495 3.38 1.265 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.55 0.475 2.55 0.475 3.62 2.33 3.62 2.33 2.965 2.67 2.965 2.67 3.62 4.57 3.62 4.57 2.965 4.91 2.965 4.91 3.62 6.81 3.62 6.81 2.965 7.15 2.965 7.15 3.62 9.105 3.62 9.105 2.55 9.335 2.55 9.335 3.62 10.08 3.62 10.08 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.435 0.3 9.435 1.04 9.205 1.04 9.205 0.3 7.25 0.3 7.25 0.985 6.91 0.985 6.91 0.3 5.01 0.3 5.01 0.985 4.67 0.985 4.67 0.3 2.77 0.3 2.77 0.985 2.43 0.985 2.43 0.3 0.475 0.3 0.475 1.04 0.245 1.04 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__clkinv_8

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 16.8 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4635 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 1.77 4.39 1.77 4.39 2.15 3.45 2.15  ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7115 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.13 0.28 2.13  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.858 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.77 0.81 16.35 0.81 16.35 2.985 15.77 2.985  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.44 3.62 1.44 2.93 1.78 2.93 1.78 3.62 2.165 3.62 3.18 3.62 3.18 3.005 3.52 3.005 3.52 3.62 6.355 3.62 7.705 3.62 7.705 2.7 8.045 2.7 8.045 3.62 9.38 3.62 12.85 3.62 12.85 3.28 13.19 3.28 13.19 3.62 14.845 3.62 14.845 2.755 15.185 2.755 15.185 3.62 15.46 3.62 16.8 3.62 16.8 4.22 15.46 4.22 9.38 4.22 6.355 4.22 2.165 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 16.8 -0.3 16.8 0.3 15.23 0.3 15.23 0.69 15 0.69 15 0.3 13.06 0.3 13.06 0.95 12.72 0.95 12.72 0.3 8.04 0.3 8.04 0.81 7.7 0.81 7.7 0.3 3.62 0.3 3.62 1.075 3.28 1.075 3.28 0.3 1.78 0.3 1.78 0.915 1.44 0.915 1.44 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.36 1.935 2.36 1.935 1.375 0.375 1.375 0.375 0.735 0.605 0.735 0.605 1.145 2.165 1.145 2.165 2.59 0.705 2.59 0.705 3.225 0.475 3.225  ;
        POLYGON 4.42 2.645 5.055 2.645 5.055 1.075 4.4 1.075 4.4 0.845 5.29 0.845 5.29 2.875 4.42 2.875  ;
        POLYGON 2.515 0.735 2.845 0.735 2.845 2.48 4.06 2.48 4.06 3.16 6.355 3.16 6.355 3.39 3.83 3.39 3.83 2.71 2.845 2.71 2.845 3.225 2.515 3.225  ;
        POLYGON 5.575 0.79 5.805 0.79 5.805 1.82 6.55 1.82 6.55 1.5 8.7 1.5 8.7 1.73 6.78 1.73 6.78 2.05 5.915 2.05 5.915 2.795 5.575 2.795  ;
        POLYGON 7.095 2.05 9.04 2.05 9.04 0.99 9.38 0.99 9.38 2.93 9.04 2.93 9.04 2.39 7.095 2.39  ;
        POLYGON 6.09 1.04 8.33 1.04 8.33 0.53 11.425 0.53 11.425 2.095 11.195 2.095 11.195 0.76 8.56 0.76 8.56 1.27 6.32 1.27 6.32 1.59 6.09 1.59  ;
        POLYGON 10.16 0.99 10.5 0.99 10.5 2.355 13.29 2.355 13.29 2.105 13.63 2.105 13.63 2.585 10.5 2.585 10.5 2.93 10.16 2.93  ;
        POLYGON 12.175 1.64 13.9 1.64 13.9 0.99 14.24 0.99 14.24 1.5 15 1.5 15 1.885 14.155 1.885 14.155 2.85 13.925 2.85 13.925 1.875 12.175 1.875  ;
        POLYGON 11.79 2.815 13.66 2.815 13.66 3.1 14.385 3.1 14.385 2.115 15.23 2.115 15.23 1.15 14.54 1.15 14.54 0.76 13.52 0.76 13.52 1.41 11.655 1.41 11.655 0.89 11.885 0.89 11.885 1.18 13.29 1.18 13.29 0.53 14.77 0.53 14.77 0.92 15.46 0.92 15.46 2.345 14.615 2.345 14.615 3.33 13.43 3.33 13.43 3.05 11.79 3.05  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 18.48 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4635 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 1.77 4.39 1.77 4.39 2.15 3.45 2.15  ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7115 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.13 0.28 2.13  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.4016 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.965 1.77 16.285 1.77 16.285 0.99 16.625 0.99 16.625 1.77 17.27 1.77 17.27 2.15 16.315 2.15 16.315 2.93 15.965 2.93  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.44 3.62 1.44 2.93 1.78 2.93 1.78 3.62 2.165 3.62 3.18 3.62 3.18 3.005 3.52 3.005 3.52 3.62 6.355 3.62 7.705 3.62 7.705 2.7 8.045 2.7 8.045 3.62 9.38 3.62 12.85 3.62 12.85 3.28 13.19 3.28 13.19 3.62 14.845 3.62 14.845 2.815 15.185 2.815 15.185 3.62 15.645 3.62 17.04 3.62 17.04 2.76 17.27 2.76 17.27 3.62 18.48 3.62 18.48 4.22 15.645 4.22 9.38 4.22 6.355 4.22 2.165 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 18.48 -0.3 18.48 0.3 17.965 0.3 17.965 0.635 17.625 0.635 17.625 0.3 15.23 0.3 15.23 0.69 15 0.69 15 0.3 13.19 0.3 13.19 0.635 12.85 0.635 12.85 0.3 8.04 0.3 8.04 0.81 7.7 0.81 7.7 0.3 3.62 0.3 3.62 1.075 3.28 1.075 3.28 0.3 1.78 0.3 1.78 0.915 1.44 0.915 1.44 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.36 1.935 2.36 1.935 1.375 0.375 1.375 0.375 0.735 0.605 0.735 0.605 1.145 2.165 1.145 2.165 2.59 0.705 2.59 0.705 3.225 0.475 3.225  ;
        POLYGON 4.42 2.645 5.055 2.645 5.055 1.075 4.4 1.075 4.4 0.845 5.29 0.845 5.29 2.875 4.42 2.875  ;
        POLYGON 2.515 0.735 2.845 0.735 2.845 2.48 4.06 2.48 4.06 3.16 6.355 3.16 6.355 3.39 3.83 3.39 3.83 2.71 2.845 2.71 2.845 3.225 2.515 3.225  ;
        POLYGON 5.575 0.79 5.805 0.79 5.805 1.82 6.55 1.82 6.55 1.5 8.7 1.5 8.7 1.73 6.78 1.73 6.78 2.05 5.915 2.05 5.915 2.795 5.575 2.795  ;
        POLYGON 7.095 2.05 9.04 2.05 9.04 0.99 9.38 0.99 9.38 2.93 9.04 2.93 9.04 2.39 7.095 2.39  ;
        POLYGON 6.09 1.04 8.33 1.04 8.33 0.53 11.51 0.53 11.51 2.04 11.17 2.04 11.17 0.76 8.56 0.76 8.56 1.27 6.32 1.27 6.32 1.59 6.09 1.59  ;
        POLYGON 10.16 0.99 10.5 0.99 10.5 2.355 13.345 2.355 13.345 2.05 13.575 2.05 13.575 2.585 10.5 2.585 10.5 2.93 10.16 2.93  ;
        POLYGON 12.41 1.495 13.97 1.495 13.97 0.99 14.31 0.99 14.31 1.715 15.075 1.715 15.075 2.055 14.155 2.055 14.155 2.85 13.925 2.85 13.925 1.73 12.41 1.73  ;
        POLYGON 11.79 2.815 13.66 2.815 13.66 3.1 14.385 3.1 14.385 2.285 15.415 2.285 15.415 1.15 14.54 1.15 14.54 0.76 13.65 0.76 13.65 1.095 11.745 1.095 11.745 0.675 11.975 0.675 11.975 0.865 13.42 0.865 13.42 0.53 14.77 0.53 14.77 0.92 15.645 0.92 15.645 2.515 14.615 2.515 14.615 3.33 13.43 3.33 13.43 3.05 11.79 3.05  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4635 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 1.77 4.39 1.77 4.39 2.15 3.45 2.15  ;
    END
  END D
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7115 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.13 0.28 2.13  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.5259 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.49 2.245 17.91 2.245 18.57 2.245 18.57 1.555 16.49 1.555 16.49 0.99 16.83 0.99 16.83 1.325 19.17 1.325 19.17 0.99 19.51 0.99 19.51 2.93 18.87 2.93 18.87 2.595 17.91 2.595 16.84 2.595 16.84 2.93 16.49 2.93  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.44 3.62 1.44 2.93 1.78 2.93 1.78 3.62 2.165 3.62 3.18 3.62 3.18 3.005 3.52 3.005 3.52 3.62 6.355 3.62 7.705 3.62 7.705 2.7 8.045 2.7 8.045 3.62 9.38 3.62 12.85 3.62 12.85 3.28 13.19 3.28 13.19 3.62 15.25 3.62 15.25 2.815 15.59 2.815 15.59 3.62 17.73 3.62 17.73 3.285 18.07 3.285 18.07 3.62 20.13 3.62 20.51 3.62 20.51 2.815 20.85 2.815 20.85 3.62 21.28 3.62 21.28 4.22 20.13 4.22 9.38 4.22 6.355 4.22 2.165 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 20.795 0.3 20.795 0.765 20.565 0.765 20.565 0.3 18.17 0.3 18.17 0.635 17.83 0.635 17.83 0.3 15.435 0.3 15.435 0.69 15.205 0.69 15.205 0.3 13.19 0.3 13.19 0.635 12.85 0.635 12.85 0.3 8.04 0.3 8.04 0.81 7.7 0.81 7.7 0.3 3.62 0.3 3.62 1.075 3.28 1.075 3.28 0.3 1.78 0.3 1.78 0.915 1.44 0.915 1.44 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.36 1.935 2.36 1.935 1.375 0.375 1.375 0.375 0.735 0.605 0.735 0.605 1.145 2.165 1.145 2.165 2.59 0.705 2.59 0.705 3.225 0.475 3.225  ;
        POLYGON 4.42 2.645 5.055 2.645 5.055 1.075 4.4 1.075 4.4 0.845 5.29 0.845 5.29 2.875 4.42 2.875  ;
        POLYGON 2.515 0.735 2.845 0.735 2.845 2.48 4.06 2.48 4.06 3.16 6.355 3.16 6.355 3.39 3.83 3.39 3.83 2.71 2.845 2.71 2.845 3.225 2.515 3.225  ;
        POLYGON 5.575 0.79 5.805 0.79 5.805 1.82 6.55 1.82 6.55 1.5 8.7 1.5 8.7 1.73 6.78 1.73 6.78 2.05 5.915 2.05 5.915 2.795 5.575 2.795  ;
        POLYGON 7.095 2.05 9.04 2.05 9.04 0.99 9.38 0.99 9.38 2.93 9.04 2.93 9.04 2.39 7.095 2.39  ;
        POLYGON 6.09 1.04 8.33 1.04 8.33 0.53 11.51 0.53 11.51 2.04 11.17 2.04 11.17 0.76 8.56 0.76 8.56 1.27 6.32 1.27 6.32 1.59 6.09 1.59  ;
        POLYGON 10.16 0.99 10.5 0.99 10.5 2.355 13.43 2.355 13.43 2.105 13.77 2.105 13.77 2.585 10.5 2.585 10.5 2.93 10.16 2.93  ;
        POLYGON 12.41 1.495 14.15 1.495 14.15 0.99 14.49 0.99 14.49 1.785 17.91 1.785 17.91 2.015 14.43 2.015 14.43 2.795 14.09 2.795 14.09 1.73 12.41 1.73  ;
        POLYGON 11.79 2.815 13.73 2.815 13.73 3.025 14.79 3.025 14.79 2.295 16.055 2.295 16.055 3.16 17.27 3.16 17.27 2.825 18.53 2.825 18.53 3.16 19.9 3.16 19.9 0.76 18.63 0.76 18.63 1.095 17.37 1.095 17.37 0.76 15.895 0.76 15.895 1.15 14.745 1.15 14.745 0.76 13.65 0.76 13.65 1.095 11.745 1.095 11.745 0.675 11.975 0.675 11.975 0.865 13.42 0.865 13.42 0.53 14.975 0.53 14.975 0.92 15.665 0.92 15.665 0.53 17.6 0.53 17.6 0.865 18.4 0.865 18.4 0.53 20.13 0.53 20.13 3.39 18.3 3.39 18.3 3.055 17.5 3.055 17.5 3.39 15.825 3.39 15.825 2.525 15.02 2.525 15.02 3.255 13.5 3.255 13.5 3.05 11.79 3.05  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.614 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 3.895 1.77 3.895 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.318 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.65 0.6 16.3 0.6 16.3 1.02 15.14 1.02 15.14 1.83 14.65 1.83  ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.29 1.77 1.575 1.77 1.575 2.15 0.29 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8668 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.45 2.33 18.04 2.33 18.57 2.33 18.57 0.83 18.38 0.83 18.38 0.6 18.92 0.6 18.92 3.32 18.365 3.32 18.365 2.765 18.04 2.765 17.45 2.765  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 2.035 3.62 3.17 3.62 3.17 2.845 3.51 2.845 3.51 3.62 5.015 3.62 7.59 3.62 7.59 3.005 7.93 3.005 7.93 3.62 9.17 3.62 9.605 3.62 9.605 2.79 9.835 2.79 9.835 3.62 10.33 3.62 10.855 3.62 14.22 3.62 14.22 3.28 14.56 3.28 14.56 3.62 16.385 3.62 16.595 3.62 16.595 2.69 16.825 2.69 16.825 3.62 17.415 3.62 17.415 3.16 17.645 3.16 17.645 3.62 18.04 3.62 19.04 3.62 19.04 4.22 18.04 4.22 16.385 4.22 10.855 4.22 10.33 4.22 9.17 4.22 5.015 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 17.545 0.3 17.545 0.93 17.315 0.93 17.315 0.3 14.405 0.3 14.405 1.13 14.175 1.13 14.175 0.3 8.87 0.3 8.87 0.915 8.53 0.915 8.53 0.3 3.49 0.3 3.49 1.075 3.15 1.075 3.15 0.3 1.65 0.3 1.65 0.915 1.31 0.915 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.465 1.805 2.465 1.805 1.375 0.245 1.375 0.245 0.63 0.475 0.63 0.475 1.145 2.035 1.145 2.035 2.7 0.575 2.7 0.575 2.805 0.345 2.805  ;
        POLYGON 4.245 0.79 4.555 0.79 4.555 2.8 4.245 2.8  ;
        POLYGON 2.615 2.38 4.015 2.38 4.015 3.16 4.785 3.16 4.785 1.555 5.015 1.555 5.015 3.39 3.785 3.39 3.785 2.61 2.615 2.61 2.615 2.805 2.385 2.805 2.385 0.63 2.715 0.63 2.715 0.97 2.615 0.97  ;
        POLYGON 6.285 2.545 8.39 2.545 8.39 2.83 9.17 2.83 9.17 3.06 8.16 3.06 8.16 2.775 6.515 2.775 6.515 3.115 6.285 3.115  ;
        POLYGON 5.265 0.79 5.675 0.79 5.675 2.085 8.85 2.085 8.85 2.24 10.33 2.24 10.33 2.47 8.62 2.47 8.62 2.315 5.495 2.315 5.495 2.8 5.265 2.8  ;
        POLYGON 6.93 1.625 10.09 1.625 10.09 0.99 10.43 0.99 10.43 1.78 10.855 1.78 10.855 3.13 10.625 3.13 10.625 2.01 10.06 2.01 10.06 1.855 6.93 1.855  ;
        POLYGON 6.17 1.165 9.1 1.165 9.1 0.53 12.625 0.53 12.625 2.525 12.395 2.525 12.395 0.76 11.255 0.76 11.255 1.62 11.025 1.62 11.025 0.76 9.33 0.76 9.33 1.395 6.515 1.395 6.515 1.565 6.17 1.565  ;
        POLYGON 12.98 0.82 13.32 0.82 13.32 2.93 12.98 2.93  ;
        POLYGON 11.645 0.99 11.995 0.99 11.995 2.065 12.105 2.065 12.105 3.16 13.67 3.16 13.67 2.815 15.02 2.815 15.02 3.16 16.135 3.16 16.135 2.035 16.385 2.035 16.385 2.375 16.365 2.375 16.365 3.39 14.79 3.39 14.79 3.05 13.9 3.05 13.9 3.39 11.875 3.39 11.875 2.405 11.645 2.405  ;
        POLYGON 13.56 2.235 15.56 2.235 15.56 1.505 16.595 1.505 16.595 0.79 16.825 0.79 16.825 1.505 18.04 1.505 18.04 1.735 15.79 1.735 15.79 2.93 15.45 2.93 15.45 2.47 13.56 2.47  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.614 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 3.895 1.77 3.895 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.393 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.65 0.65 15.14 0.65 15.14 1.59 14.65 1.59  ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.575 1.77 1.575 2.15 0.71 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0296 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.38 2.33 18.61 2.33 19.13 2.33 19.13 1.175 18.435 1.175 18.435 0.79 18.665 0.79 18.665 0.945 19.51 0.945 19.51 2.765 18.72 2.765 18.72 3.235 18.61 3.235 18.38 3.235  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 2.035 3.62 3.17 3.62 3.17 2.845 3.51 2.845 3.51 3.62 5.015 3.62 7.59 3.62 7.59 3.005 7.93 3.005 7.93 3.62 9.17 3.62 9.605 3.62 9.605 2.79 9.835 2.79 9.835 3.62 10.33 3.62 10.855 3.62 14.22 3.62 14.22 3.28 14.56 3.28 14.56 3.62 16.385 3.62 16.595 3.62 16.595 2.69 16.825 2.69 16.825 3.62 17.415 3.62 17.415 2.69 17.645 2.69 17.645 3.62 18.61 3.62 19.455 3.62 19.455 3.16 19.685 3.16 19.685 3.62 20.16 3.62 20.16 4.22 18.61 4.22 16.385 4.22 10.855 4.22 10.33 4.22 9.17 4.22 5.015 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 19.84 0.3 19.84 0.715 19.5 0.715 19.5 0.3 17.545 0.3 17.545 0.765 17.315 0.765 17.315 0.3 14.405 0.3 14.405 1.13 14.175 1.13 14.175 0.3 8.87 0.3 8.87 0.915 8.53 0.915 8.53 0.3 3.49 0.3 3.49 1.075 3.15 1.075 3.15 0.3 1.65 0.3 1.65 0.915 1.31 0.915 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.465 1.805 2.465 1.805 1.375 0.245 1.375 0.245 0.63 0.475 0.63 0.475 1.145 2.035 1.145 2.035 2.7 0.575 2.7 0.575 2.805 0.345 2.805  ;
        POLYGON 4.245 0.79 4.555 0.79 4.555 2.8 4.245 2.8  ;
        POLYGON 2.615 2.38 4.015 2.38 4.015 3.16 4.785 3.16 4.785 1.555 5.015 1.555 5.015 3.39 3.785 3.39 3.785 2.61 2.615 2.61 2.615 2.805 2.385 2.805 2.385 0.63 2.715 0.63 2.715 0.97 2.615 0.97  ;
        POLYGON 6.285 2.545 8.39 2.545 8.39 2.83 9.17 2.83 9.17 3.06 8.16 3.06 8.16 2.775 6.515 2.775 6.515 3.115 6.285 3.115  ;
        POLYGON 5.265 0.79 5.675 0.79 5.675 2.085 8.85 2.085 8.85 2.24 10.33 2.24 10.33 2.47 8.62 2.47 8.62 2.315 5.495 2.315 5.495 2.8 5.265 2.8  ;
        POLYGON 6.93 1.625 10.09 1.625 10.09 0.99 10.43 0.99 10.43 1.78 10.855 1.78 10.855 3.13 10.625 3.13 10.625 2.01 10.06 2.01 10.06 1.855 6.93 1.855  ;
        POLYGON 6.17 1.165 9.1 1.165 9.1 0.53 12.625 0.53 12.625 2.525 12.395 2.525 12.395 0.76 11.255 0.76 11.255 1.62 11.025 1.62 11.025 0.76 9.33 0.76 9.33 1.395 6.515 1.395 6.515 1.565 6.17 1.565  ;
        POLYGON 12.98 0.82 13.32 0.82 13.32 2.93 12.98 2.93  ;
        POLYGON 11.645 0.99 11.995 0.99 11.995 2.065 12.105 2.065 12.105 3.16 13.67 3.16 13.67 2.815 15.02 2.815 15.02 3.155 16.135 3.155 16.135 2.035 16.385 2.035 16.385 2.375 16.365 2.375 16.365 3.39 14.79 3.39 14.79 3.05 13.9 3.05 13.9 3.39 11.875 3.39 11.875 2.405 11.645 2.405  ;
        POLYGON 13.56 1.77 13.9 1.77 13.9 2.235 15.56 2.235 15.56 1.505 16.595 1.505 16.595 0.74 16.825 0.74 16.825 1.505 18.61 1.505 18.61 1.735 15.79 1.735 15.79 2.87 15.45 2.87 15.45 2.47 13.56 2.47  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.614 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 3.895 1.77 3.895 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.3955 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.65 0.65 15.14 0.65 15.14 1.59 14.65 1.59  ;
    END
  END RN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.77 1.575 1.77 1.575 2.15 0.71 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.08 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.38 2.33 20.28 2.33 20.81 2.33 20.81 1.175 18.435 1.175 18.435 0.79 18.665 0.79 18.665 0.945 20.635 0.945 20.635 0.79 21.19 0.79 21.19 2.765 20.76 2.765 20.76 3.235 20.42 3.235 20.42 2.765 20.28 2.765 18.72 2.765 18.72 3.235 18.38 3.235  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 2.035 3.62 3.17 3.62 3.17 2.845 3.51 2.845 3.51 3.62 5.015 3.62 7.59 3.62 7.59 3.005 7.93 3.005 7.93 3.62 9.17 3.62 9.605 3.62 9.605 2.79 9.835 2.79 9.835 3.62 10.33 3.62 10.855 3.62 14.22 3.62 14.22 3.28 14.56 3.28 14.56 3.62 16.385 3.62 16.595 3.62 16.595 2.69 16.825 2.69 16.825 3.62 17.415 3.62 17.415 2.69 17.645 2.69 17.645 3.62 19.455 3.62 19.455 3.16 19.685 3.16 19.685 3.62 20.28 3.62 21.495 3.62 21.495 2.69 21.725 2.69 21.725 3.62 22.4 3.62 22.4 4.22 20.28 4.22 16.385 4.22 10.855 4.22 10.33 4.22 9.17 4.22 5.015 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 22.025 0.3 22.025 0.765 21.795 0.765 21.795 0.3 19.84 0.3 19.84 0.715 19.5 0.715 19.5 0.3 17.545 0.3 17.545 0.765 17.315 0.765 17.315 0.3 14.405 0.3 14.405 1.13 14.175 1.13 14.175 0.3 8.87 0.3 8.87 0.915 8.53 0.915 8.53 0.3 3.49 0.3 3.49 1.075 3.15 1.075 3.15 0.3 1.65 0.3 1.65 0.915 1.31 0.915 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.465 1.805 2.465 1.805 1.375 0.245 1.375 0.245 0.63 0.475 0.63 0.475 1.145 2.035 1.145 2.035 2.7 0.575 2.7 0.575 2.805 0.345 2.805  ;
        POLYGON 4.245 0.79 4.555 0.79 4.555 2.8 4.245 2.8  ;
        POLYGON 2.615 2.38 4.015 2.38 4.015 3.16 4.785 3.16 4.785 1.555 5.015 1.555 5.015 3.39 3.785 3.39 3.785 2.61 2.615 2.61 2.615 2.805 2.385 2.805 2.385 0.63 2.715 0.63 2.715 0.97 2.615 0.97  ;
        POLYGON 6.285 2.545 8.39 2.545 8.39 2.83 9.17 2.83 9.17 3.06 8.16 3.06 8.16 2.775 6.515 2.775 6.515 3.115 6.285 3.115  ;
        POLYGON 5.265 0.79 5.675 0.79 5.675 2.085 8.85 2.085 8.85 2.24 10.33 2.24 10.33 2.47 8.62 2.47 8.62 2.315 5.495 2.315 5.495 2.8 5.265 2.8  ;
        POLYGON 6.93 1.625 10.09 1.625 10.09 0.99 10.43 0.99 10.43 1.78 10.855 1.78 10.855 3.13 10.625 3.13 10.625 2.01 10.06 2.01 10.06 1.855 6.93 1.855  ;
        POLYGON 6.17 1.165 9.1 1.165 9.1 0.53 12.625 0.53 12.625 2.525 12.395 2.525 12.395 0.76 11.255 0.76 11.255 1.62 11.025 1.62 11.025 0.76 9.33 0.76 9.33 1.395 6.515 1.395 6.515 1.565 6.17 1.565  ;
        POLYGON 12.98 0.82 13.32 0.82 13.32 2.93 12.98 2.93  ;
        POLYGON 11.645 0.99 11.995 0.99 11.995 2.065 12.105 2.065 12.105 3.16 13.67 3.16 13.67 2.815 15.02 2.815 15.02 3.155 16.135 3.155 16.135 2.035 16.385 2.035 16.385 2.375 16.365 2.375 16.365 3.39 14.79 3.39 14.79 3.05 13.9 3.05 13.9 3.39 11.875 3.39 11.875 2.405 11.645 2.405  ;
        POLYGON 13.56 1.77 13.9 1.77 13.9 2.235 15.56 2.235 15.56 1.435 16.595 1.435 16.595 0.74 16.825 0.74 16.825 1.435 20.28 1.435 20.28 1.665 15.79 1.665 15.79 2.87 15.45 2.87 15.45 2.47 13.56 2.47  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 24.08 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.433 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 4.05 1.77 4.05 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.284 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.38 1.77 20.63 1.77 20.63 2.15 19.38 2.15  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1495 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.45 1.77 18.28 1.77 18.28 1.32 18.55 1.32 18.55 2.15 17.45 2.15  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.15 0.28 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8954 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.585 0.55 23.96 0.55 23.96 3.38 23.585 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 3.005 1.65 3.005 1.65 3.62 2.055 3.62 3.05 3.62 3.05 3 3.39 3 3.39 3.62 7.585 3.62 7.585 3.165 7.93 3.165 7.93 3.62 13.45 3.62 13.45 3.035 13.68 3.035 13.68 3.62 15.48 3.62 17.705 3.62 17.705 2.94 18.045 2.94 18.045 3.62 19.745 3.62 19.745 2.94 20.085 2.94 20.085 3.62 21.61 3.62 21.84 3.62 21.84 2.415 22.07 2.415 22.07 3.62 22.58 3.62 22.58 2.565 22.81 2.565 22.81 3.62 23.25 3.62 24.08 3.62 24.08 4.22 23.25 4.22 21.61 4.22 15.48 4.22 2.055 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 24.08 -0.3 24.08 0.3 22.71 0.3 22.71 0.93 22.48 0.93 22.48 0.3 20.085 0.3 20.085 1.075 19.745 1.075 19.745 0.3 10.92 0.3 10.92 0.915 10.58 0.915 10.58 0.3 3.61 0.3 3.61 1.075 3.27 1.075 3.27 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.435 1.825 2.435 1.825 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.055 1.28 2.055 2.67 0.575 2.67 0.575 3.3 0.345 3.3  ;
        POLYGON 4.29 0.845 4.73 0.845 4.73 2.83 4.29 2.83  ;
        POLYGON 6.405 2.245 8.97 2.245 8.97 2.585 10.85 2.585 10.85 2.875 10.51 2.875 10.51 2.815 8.74 2.815 8.74 2.475 6.635 2.475 6.635 2.87 6.405 2.87  ;
        POLYGON 5.31 1.785 5.565 1.785 5.565 0.79 5.795 0.79 5.795 1.785 9.43 1.785 9.43 2.07 12.07 2.07 12.07 1.545 12.47 1.545 12.47 1.775 12.3 1.775 12.3 2.3 9.2 2.3 9.2 2.015 5.65 2.015 5.65 2.83 5.31 2.83  ;
        POLYGON 11.79 2.645 12.53 2.645 12.53 2.115 14.465 2.115 14.465 1.315 11.84 1.315 11.84 1.835 9.66 1.835 9.66 1.555 7.03 1.555 7.03 1.325 9.89 1.325 9.89 1.605 11.61 1.605 11.61 1.085 14.75 1.085 14.75 2.125 14.975 2.125 14.975 2.875 14.635 2.875 14.635 2.345 12.76 2.345 12.76 2.875 11.79 2.875  ;
        POLYGON 2.615 2.54 4.015 2.54 4.015 3.105 6.865 3.105 6.865 2.705 8.51 2.705 8.51 3.16 12.99 3.16 12.99 2.575 14.405 2.575 14.405 3.16 15.25 3.16 15.25 2.07 15.48 2.07 15.48 3.39 14.175 3.39 14.175 2.805 13.22 2.805 13.22 3.39 8.28 3.39 8.28 2.935 7.095 2.935 7.095 3.335 3.785 3.335 3.785 2.77 2.615 2.77 2.615 3.3 2.385 3.3 2.385 0.81 2.715 0.81 2.715 1.15 2.615 1.15  ;
        POLYGON 6.135 0.79 10.35 0.79 10.35 1.145 11.15 1.145 11.15 0.53 17.115 0.53 17.115 0.855 16.775 0.855 16.775 0.76 14.77 0.76 14.77 0.855 14.43 0.855 14.43 0.76 11.38 0.76 11.38 1.375 10.12 1.375 10.12 1.02 6.475 1.02 6.475 1.555 6.135 1.555  ;
        POLYGON 16.17 1.03 16.455 1.03 16.455 1.085 17.64 1.085 17.64 0.79 19.01 0.79 19.01 2.855 18.78 2.855 18.78 1.075 17.925 1.075 17.925 1.315 17.015 1.315 17.015 2.895 16.675 2.895 16.675 1.37 16.17 1.37  ;
        POLYGON 14.98 1.085 15.94 1.085 15.94 3.16 17.245 3.16 17.245 2.475 18.505 2.475 18.505 3.085 19.24 3.085 19.24 2.48 20.545 2.48 20.545 3.085 21.38 3.085 21.38 1.91 21.61 1.91 21.61 3.32 20.315 3.32 20.315 2.71 19.47 2.71 19.47 3.32 18.275 3.32 18.275 2.71 17.475 2.71 17.475 3.39 15.71 3.39 15.71 1.315 14.98 1.315  ;
        POLYGON 20.82 2.515 20.92 2.515 20.92 1.54 19.305 1.54 19.305 1.31 21.76 1.31 21.76 0.79 21.99 0.79 21.99 1.33 23.25 1.33 23.25 1.56 21.15 1.56 21.15 2.855 20.82 2.855  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 25.2 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.433 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 4.05 1.77 4.05 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.284 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.38 1.77 20.63 1.77 20.63 2.15 19.38 2.15  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1495 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.45 1.77 18.225 1.77 18.225 1.34 18.54 1.34 18.54 2.15 17.45 2.15  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.15 0.28 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0582 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.545 2.07 23.72 2.07 24.17 2.07 24.17 1.17 23.6 1.17 23.6 0.55 23.98 0.55 23.98 0.94 24.55 0.94 24.55 2.32 23.98 2.32 23.98 3.38 23.72 3.38 23.545 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 3.005 1.65 3.005 1.65 3.62 2.055 3.62 3.05 3.62 3.05 3 3.39 3 3.39 3.62 7.585 3.62 7.585 3.165 7.93 3.165 7.93 3.62 13.45 3.62 13.45 3.035 13.68 3.035 13.68 3.62 15.48 3.62 17.705 3.62 17.705 2.94 18.045 2.94 18.045 3.62 19.745 3.62 19.745 2.94 20.085 2.94 20.085 3.62 21.61 3.62 21.84 3.62 21.84 2.415 22.07 2.415 22.07 3.62 22.58 3.62 22.58 2.57 22.81 2.57 22.81 3.62 23.72 3.62 24.62 3.62 24.62 2.57 24.85 2.57 24.85 3.62 25.2 3.62 25.2 4.22 23.72 4.22 21.61 4.22 15.48 4.22 2.055 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 25.2 -0.3 25.2 0.3 25.005 0.3 25.005 0.71 24.665 0.71 24.665 0.3 22.71 0.3 22.71 0.765 22.48 0.765 22.48 0.3 20.085 0.3 20.085 1.075 19.745 1.075 19.745 0.3 10.92 0.3 10.92 0.915 10.58 0.915 10.58 0.3 3.61 0.3 3.61 1.075 3.27 1.075 3.27 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.435 1.825 2.435 1.825 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.055 1.28 2.055 2.67 0.575 2.67 0.575 3.3 0.345 3.3  ;
        POLYGON 4.29 0.845 4.73 0.845 4.73 2.83 4.29 2.83  ;
        POLYGON 6.405 2.245 8.97 2.245 8.97 2.585 10.85 2.585 10.85 2.875 10.51 2.875 10.51 2.815 8.74 2.815 8.74 2.475 6.635 2.475 6.635 2.87 6.405 2.87  ;
        POLYGON 5.31 1.785 5.565 1.785 5.565 0.79 5.795 0.79 5.795 1.785 9.43 1.785 9.43 2.07 12.07 2.07 12.07 1.545 12.47 1.545 12.47 1.775 12.3 1.775 12.3 2.3 9.2 2.3 9.2 2.015 5.65 2.015 5.65 2.83 5.31 2.83  ;
        POLYGON 11.79 2.645 12.53 2.645 12.53 2.115 14.465 2.115 14.465 1.315 11.84 1.315 11.84 1.835 9.66 1.835 9.66 1.555 7.03 1.555 7.03 1.325 9.89 1.325 9.89 1.605 11.61 1.605 11.61 1.085 14.75 1.085 14.75 2.125 14.975 2.125 14.975 2.875 14.635 2.875 14.635 2.345 12.76 2.345 12.76 2.875 11.79 2.875  ;
        POLYGON 2.615 2.54 4.015 2.54 4.015 3.105 6.865 3.105 6.865 2.705 8.51 2.705 8.51 3.16 12.99 3.16 12.99 2.575 14.405 2.575 14.405 3.16 15.25 3.16 15.25 2.07 15.48 2.07 15.48 3.39 14.175 3.39 14.175 2.805 13.22 2.805 13.22 3.39 8.28 3.39 8.28 2.935 7.095 2.935 7.095 3.335 3.785 3.335 3.785 2.77 2.615 2.77 2.615 3.3 2.385 3.3 2.385 0.81 2.715 0.81 2.715 1.15 2.615 1.15  ;
        POLYGON 6.135 0.79 10.35 0.79 10.35 1.145 11.15 1.145 11.15 0.53 17.115 0.53 17.115 0.855 16.775 0.855 16.775 0.76 14.77 0.76 14.77 0.855 14.43 0.855 14.43 0.76 11.38 0.76 11.38 1.375 10.12 1.375 10.12 1.02 6.475 1.02 6.475 1.555 6.135 1.555  ;
        POLYGON 16.17 1.03 16.455 1.03 16.455 1.085 17.71 1.085 17.71 0.79 19.01 0.79 19.01 2.855 18.78 2.855 18.78 1.075 17.995 1.075 17.995 1.315 17.015 1.315 17.015 2.895 16.675 2.895 16.675 1.37 16.17 1.37  ;
        POLYGON 14.98 1.085 15.94 1.085 15.94 3.16 17.245 3.16 17.245 2.475 18.505 2.475 18.505 3.085 19.24 3.085 19.24 2.48 20.545 2.48 20.545 3.085 21.38 3.085 21.38 1.91 21.61 1.91 21.61 3.32 20.315 3.32 20.315 2.71 19.47 2.71 19.47 3.32 18.275 3.32 18.275 2.71 17.475 2.71 17.475 3.39 15.71 3.39 15.71 1.315 14.98 1.315  ;
        POLYGON 20.82 2.515 20.92 2.515 20.92 1.54 19.305 1.54 19.305 1.31 21.76 1.31 21.76 0.79 21.99 0.79 21.99 1.33 23.305 1.33 23.305 1.475 23.72 1.475 23.72 1.82 22.965 1.82 22.965 1.56 21.15 1.56 21.15 2.855 20.82 2.855  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 27.44 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.433 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 4.05 1.77 4.05 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.284 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.38 1.77 20.63 1.77 20.63 2.15 19.38 2.15  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1495 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.45 1.77 18.225 1.77 18.225 1.32 18.54 1.32 18.54 2.15 17.45 2.15  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.15 0.28 2.15  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1112 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.545 2.1 25.39 2.1 25.85 2.1 25.85 1.17 23.6 1.17 23.6 0.55 23.83 0.55 23.83 0.94 25.84 0.94 25.84 0.55 26.23 0.55 26.23 3.38 25.585 3.38 25.585 2.33 25.39 2.33 23.885 2.33 23.885 3.38 23.545 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 3.005 1.65 3.005 1.65 3.62 2.055 3.62 3.05 3.62 3.05 3 3.39 3 3.39 3.62 7.585 3.62 7.585 3.165 7.93 3.165 7.93 3.62 13.45 3.62 13.45 3.035 13.68 3.035 13.68 3.62 15.48 3.62 17.705 3.62 17.705 2.94 18.045 2.94 18.045 3.62 19.745 3.62 19.745 2.94 20.085 2.94 20.085 3.62 21.61 3.62 21.84 3.62 21.84 2.415 22.07 2.415 22.07 3.62 22.58 3.62 22.58 2.57 22.81 2.57 22.81 3.62 24.62 3.62 24.62 2.57 24.85 2.57 24.85 3.62 25.39 3.62 26.66 3.62 26.66 2.57 26.89 2.57 26.89 3.62 27.44 3.62 27.44 4.22 25.39 4.22 21.61 4.22 15.48 4.22 2.055 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 27.44 -0.3 27.44 0.3 27.19 0.3 27.19 0.765 26.96 0.765 26.96 0.3 25.005 0.3 25.005 0.71 24.665 0.71 24.665 0.3 22.71 0.3 22.71 0.765 22.48 0.765 22.48 0.3 20.085 0.3 20.085 1.075 19.745 1.075 19.745 0.3 10.92 0.3 10.92 0.915 10.58 0.915 10.58 0.3 3.61 0.3 3.61 1.075 3.27 1.075 3.27 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.435 1.825 2.435 1.825 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.055 1.28 2.055 2.67 0.575 2.67 0.575 3.3 0.345 3.3  ;
        POLYGON 4.29 0.845 4.73 0.845 4.73 2.83 4.29 2.83  ;
        POLYGON 6.405 2.245 8.97 2.245 8.97 2.585 10.85 2.585 10.85 2.875 10.51 2.875 10.51 2.815 8.74 2.815 8.74 2.475 6.635 2.475 6.635 2.87 6.405 2.87  ;
        POLYGON 5.31 1.785 5.565 1.785 5.565 0.79 5.795 0.79 5.795 1.785 9.43 1.785 9.43 2.07 12.07 2.07 12.07 1.545 12.47 1.545 12.47 1.775 12.3 1.775 12.3 2.3 9.2 2.3 9.2 2.015 5.65 2.015 5.65 2.83 5.31 2.83  ;
        POLYGON 11.79 2.645 12.53 2.645 12.53 2.115 14.465 2.115 14.465 1.315 11.84 1.315 11.84 1.835 9.66 1.835 9.66 1.555 7.03 1.555 7.03 1.325 9.89 1.325 9.89 1.605 11.61 1.605 11.61 1.085 14.75 1.085 14.75 2.125 14.975 2.125 14.975 2.875 14.635 2.875 14.635 2.345 12.76 2.345 12.76 2.875 11.79 2.875  ;
        POLYGON 2.615 2.54 4.015 2.54 4.015 3.105 6.865 3.105 6.865 2.705 8.51 2.705 8.51 3.16 12.99 3.16 12.99 2.575 14.405 2.575 14.405 3.16 15.25 3.16 15.25 2.07 15.48 2.07 15.48 3.39 14.175 3.39 14.175 2.805 13.22 2.805 13.22 3.39 8.28 3.39 8.28 2.935 7.095 2.935 7.095 3.335 3.785 3.335 3.785 2.77 2.615 2.77 2.615 3.3 2.385 3.3 2.385 0.81 2.715 0.81 2.715 1.15 2.615 1.15  ;
        POLYGON 6.135 0.79 10.35 0.79 10.35 1.145 11.15 1.145 11.15 0.53 17.115 0.53 17.115 0.855 16.775 0.855 16.775 0.76 14.77 0.76 14.77 0.855 14.43 0.855 14.43 0.76 11.38 0.76 11.38 1.375 10.12 1.375 10.12 1.02 6.475 1.02 6.475 1.555 6.135 1.555  ;
        POLYGON 16.17 1.03 16.455 1.03 16.455 1.085 17.675 1.085 17.675 0.79 19.01 0.79 19.01 2.855 18.78 2.855 18.78 1.075 17.96 1.075 17.96 1.315 17.015 1.315 17.015 2.895 16.675 2.895 16.675 1.37 16.17 1.37  ;
        POLYGON 14.98 1.085 15.94 1.085 15.94 3.16 17.245 3.16 17.245 2.475 18.505 2.475 18.505 3.085 19.24 3.085 19.24 2.48 20.545 2.48 20.545 3.085 21.38 3.085 21.38 1.91 21.61 1.91 21.61 3.32 20.315 3.32 20.315 2.71 19.47 2.71 19.47 3.32 18.275 3.32 18.275 2.71 17.475 2.71 17.475 3.39 15.71 3.39 15.71 1.315 14.98 1.315  ;
        POLYGON 20.82 2.515 20.92 2.515 20.92 1.54 19.305 1.54 19.305 1.31 21.76 1.31 21.76 0.79 21.99 0.79 21.99 1.33 23.305 1.33 23.305 1.475 25.39 1.475 25.39 1.82 22.965 1.82 22.965 1.56 21.15 1.56 21.15 2.855 20.82 2.855  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnrsnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5305 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 1.77 4.39 1.77 4.39 2.15 3.45 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1565 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.56 1.22 15.59 1.22 15.59 1.67 14.56 1.67  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.794 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.13 0.28 2.13  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8932 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.61 0.55 20.04 0.55 20.04 3.38 19.61 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 3.005 1.65 3.005 1.65 3.62 2.155 3.62 3.05 3.62 3.05 3.005 3.39 3.005 3.39 3.62 7.29 3.62 7.29 3.24 7.63 3.24 7.63 3.62 9.825 3.62 9.825 2.885 10.055 2.885 10.055 3.62 11.67 3.62 14.11 3.62 14.11 2.945 14.45 2.945 14.45 3.62 16.745 3.62 16.745 2.6 16.975 2.6 16.975 3.62 17.47 3.62 18.645 3.62 18.645 2.53 18.875 2.53 18.875 3.62 19.215 3.62 20.16 3.62 20.16 4.22 19.215 4.22 17.47 4.22 11.67 4.22 2.155 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 18.775 0.3 18.775 0.835 18.545 0.835 18.545 0.3 16.99 0.3 16.99 1.08 16.65 1.08 16.65 0.3 7.81 0.3 7.81 1.09 7.47 1.09 7.47 0.3 3.455 0.3 3.455 1.145 3.225 1.145 3.225 0.3 1.65 0.3 1.65 0.935 1.31 0.935 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.36 1.925 2.36 1.925 1.395 0.245 1.395 0.245 0.66 0.475 0.66 0.475 1.165 2.155 1.165 2.155 2.595 0.575 2.595 0.575 3.3 0.345 3.3  ;
        POLYGON 4.29 2.52 4.86 2.52 4.86 1.095 4.29 1.095 4.29 0.865 5.09 0.865 5.09 2.75 4.29 2.75  ;
        POLYGON 5.365 0.865 5.85 0.865 5.85 1.395 8.29 1.395 8.29 1.63 5.595 1.63 5.595 2.71 5.365 2.71  ;
        POLYGON 6.63 1.965 9.825 1.965 9.825 0.81 10.055 0.81 10.055 1.93 11.23 1.93 11.23 2.655 10.89 2.655 10.89 2.195 8.87 2.195 8.87 2.655 8.53 2.655 8.53 2.195 6.63 2.195  ;
        POLYGON 2.385 0.66 2.715 0.66 2.715 2.545 3.85 2.545 3.85 3.12 5.94 3.12 5.94 2.65 8.205 2.65 8.205 2.885 9.1 2.885 9.1 2.425 10.515 2.425 10.515 3.065 11.67 3.065 11.67 3.295 10.285 3.295 10.285 2.655 9.33 2.655 9.33 3.115 7.975 3.115 7.975 2.88 6.23 2.88 6.23 3.36 3.62 3.36 3.62 2.775 2.715 2.775 2.715 3.3 2.385 3.3  ;
        POLYGON 13.395 1.965 15.73 1.965 15.73 2.655 15.38 2.655 15.38 2.195 13.395 2.195 13.395 2.71 13.165 2.71 13.165 1.075 12.01 1.075 12.01 0.795 14.295 0.795 14.295 1.135 13.395 1.135  ;
        POLYGON 10.945 0.81 11.175 0.81 11.175 1.355 12.375 1.355 12.375 2.94 13.625 2.94 13.625 2.48 14.985 2.48 14.985 2.885 16.15 2.885 16.15 1.96 17.47 1.96 17.47 2.195 16.38 2.195 16.38 3.12 14.755 3.12 14.755 2.715 13.855 2.715 13.855 3.175 12.145 3.175 12.145 1.585 10.945 1.585  ;
        POLYGON 15.99 1.385 17.825 1.385 17.825 0.795 18.055 0.795 18.055 1.545 19.215 1.545 19.215 1.895 17.995 1.895 17.995 2.875 17.765 2.875 17.765 1.615 15.99 1.615  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnsnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5305 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 1.77 4.39 1.77 4.39 2.15 3.45 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1565 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.56 1.22 15.59 1.22 15.59 1.67 14.56 1.67  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.794 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.13 0.28 2.13  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.61 2.09 19.93 2.09 20.26 2.09 20.26 1.29 19.665 1.29 19.665 0.55 20.06 0.55 20.06 1.06 20.62 1.06 20.62 2.32 20.06 2.32 20.06 3.38 19.93 3.38 19.61 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 3.005 1.65 3.005 1.65 3.62 2.155 3.62 3.05 3.62 3.05 3.005 3.39 3.005 3.39 3.62 7.29 3.62 7.29 3.24 7.63 3.24 7.63 3.62 9.825 3.62 9.825 2.885 10.055 2.885 10.055 3.62 11.67 3.62 14.11 3.62 14.11 2.945 14.45 2.945 14.45 3.62 16.745 3.62 16.745 2.6 16.975 2.6 16.975 3.62 17.47 3.62 18.645 3.62 18.645 2.57 18.875 2.57 18.875 3.62 19.93 3.62 20.685 3.62 20.685 2.57 20.915 2.57 20.915 3.62 21.28 3.62 21.28 4.22 19.93 4.22 17.47 4.22 11.67 4.22 2.155 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 21.015 0.3 21.015 0.765 20.785 0.765 20.785 0.3 18.775 0.3 18.775 0.765 18.545 0.765 18.545 0.3 16.99 0.3 16.99 1.08 16.65 1.08 16.65 0.3 7.81 0.3 7.81 1.09 7.47 1.09 7.47 0.3 3.455 0.3 3.455 1.145 3.225 1.145 3.225 0.3 1.65 0.3 1.65 0.935 1.31 0.935 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.36 1.925 2.36 1.925 1.395 0.245 1.395 0.245 0.66 0.475 0.66 0.475 1.165 2.155 1.165 2.155 2.595 0.575 2.595 0.575 3.3 0.345 3.3  ;
        POLYGON 4.29 2.52 4.86 2.52 4.86 1.095 4.29 1.095 4.29 0.865 5.09 0.865 5.09 2.75 4.29 2.75  ;
        POLYGON 5.365 0.865 5.85 0.865 5.85 1.395 8.29 1.395 8.29 1.63 5.595 1.63 5.595 2.71 5.365 2.71  ;
        POLYGON 6.63 1.965 9.825 1.965 9.825 0.81 10.055 0.81 10.055 1.93 11.23 1.93 11.23 2.655 10.89 2.655 10.89 2.195 8.87 2.195 8.87 2.655 8.53 2.655 8.53 2.195 6.63 2.195  ;
        POLYGON 2.385 0.66 2.715 0.66 2.715 2.545 3.85 2.545 3.85 3.12 5.94 3.12 5.94 2.65 8.205 2.65 8.205 2.885 9.1 2.885 9.1 2.425 10.515 2.425 10.515 3.065 11.67 3.065 11.67 3.295 10.285 3.295 10.285 2.655 9.33 2.655 9.33 3.115 7.975 3.115 7.975 2.88 6.23 2.88 6.23 3.36 3.62 3.36 3.62 2.775 2.715 2.775 2.715 3.3 2.385 3.3  ;
        POLYGON 13.395 1.965 15.73 1.965 15.73 2.655 15.38 2.655 15.38 2.195 13.395 2.195 13.395 2.71 13.165 2.71 13.165 1.075 12.01 1.075 12.01 0.795 14.295 0.795 14.295 1.135 13.395 1.135  ;
        POLYGON 10.945 0.81 11.175 0.81 11.175 1.355 12.375 1.355 12.375 2.94 13.625 2.94 13.625 2.48 14.985 2.48 14.985 2.885 16.15 2.885 16.15 1.96 17.47 1.96 17.47 2.195 16.38 2.195 16.38 3.12 14.755 3.12 14.755 2.715 13.855 2.715 13.855 3.175 12.145 3.175 12.145 1.585 10.945 1.585  ;
        POLYGON 15.99 1.385 17.825 1.385 17.825 0.795 18.055 0.795 18.055 1.605 19.93 1.605 19.93 1.835 17.995 1.835 17.995 2.875 17.765 2.875 17.765 1.615 15.99 1.615  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnsnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 23.52 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5305 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.45 1.77 4.39 1.77 4.39 2.15 3.45 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1565 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.56 1.22 15.59 1.22 15.59 1.67 14.56 1.67  ;
    END
  END SETN
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.794 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.13 0.28 2.13  ;
    END
  END CLKN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1112 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.665 2.09 21.56 2.09 21.93 2.09 21.93 1.29 19.665 1.29 19.665 0.805 19.895 0.805 19.895 1.06 21.905 1.06 21.905 0.55 22.31 0.55 22.31 3.38 21.69 3.38 21.69 2.32 21.56 2.32 19.895 2.32 19.895 3.38 19.665 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 3.005 1.65 3.005 1.65 3.62 2.155 3.62 3.05 3.62 3.05 3.005 3.39 3.005 3.39 3.62 7.29 3.62 7.29 3.24 7.63 3.24 7.63 3.62 9.825 3.62 9.825 2.885 10.055 2.885 10.055 3.62 11.67 3.62 14.11 3.62 14.11 2.945 14.45 2.945 14.45 3.62 16.745 3.62 16.745 2.6 16.975 2.6 16.975 3.62 17.47 3.62 18.645 3.62 18.645 2.57 18.875 2.57 18.875 3.62 20.685 3.62 20.685 2.57 20.915 2.57 20.915 3.62 21.56 3.62 22.725 3.62 22.725 2.57 22.955 2.57 22.955 3.62 23.52 3.62 23.52 4.22 21.56 4.22 17.47 4.22 11.67 4.22 2.155 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 23.52 -0.3 23.52 0.3 23.255 0.3 23.255 0.765 23.025 0.765 23.025 0.3 21.015 0.3 21.015 0.765 20.785 0.765 20.785 0.3 18.775 0.3 18.775 0.765 18.545 0.765 18.545 0.3 16.99 0.3 16.99 1.08 16.65 1.08 16.65 0.3 7.81 0.3 7.81 1.09 7.47 1.09 7.47 0.3 3.455 0.3 3.455 1.145 3.225 1.145 3.225 0.3 1.65 0.3 1.65 0.935 1.31 0.935 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.36 1.925 2.36 1.925 1.395 0.245 1.395 0.245 0.66 0.475 0.66 0.475 1.165 2.155 1.165 2.155 2.595 0.575 2.595 0.575 3.3 0.345 3.3  ;
        POLYGON 4.29 2.52 4.86 2.52 4.86 1.095 4.29 1.095 4.29 0.865 5.09 0.865 5.09 2.75 4.29 2.75  ;
        POLYGON 5.365 0.865 5.85 0.865 5.85 1.395 8.29 1.395 8.29 1.63 5.595 1.63 5.595 2.71 5.365 2.71  ;
        POLYGON 6.63 1.965 9.825 1.965 9.825 0.81 10.055 0.81 10.055 1.93 11.23 1.93 11.23 2.655 10.89 2.655 10.89 2.195 8.87 2.195 8.87 2.655 8.53 2.655 8.53 2.195 6.63 2.195  ;
        POLYGON 2.385 0.66 2.715 0.66 2.715 2.545 3.85 2.545 3.85 3.12 5.94 3.12 5.94 2.65 8.205 2.65 8.205 2.885 9.1 2.885 9.1 2.425 10.515 2.425 10.515 3.065 11.67 3.065 11.67 3.295 10.285 3.295 10.285 2.655 9.33 2.655 9.33 3.115 7.975 3.115 7.975 2.88 6.23 2.88 6.23 3.36 3.62 3.36 3.62 2.775 2.715 2.775 2.715 3.3 2.385 3.3  ;
        POLYGON 13.395 1.965 15.73 1.965 15.73 2.655 15.38 2.655 15.38 2.195 13.395 2.195 13.395 2.71 13.165 2.71 13.165 1.075 12.01 1.075 12.01 0.795 14.295 0.795 14.295 1.135 13.395 1.135  ;
        POLYGON 10.945 0.81 11.175 0.81 11.175 1.355 12.375 1.355 12.375 2.94 13.625 2.94 13.625 2.48 14.985 2.48 14.985 2.885 16.15 2.885 16.15 1.96 17.47 1.96 17.47 2.195 16.38 2.195 16.38 3.12 14.755 3.12 14.755 2.715 13.855 2.715 13.855 3.175 12.145 3.175 12.145 1.585 10.945 1.585  ;
        POLYGON 15.99 1.385 17.825 1.385 17.825 0.795 18.055 0.795 18.055 1.605 21.56 1.605 21.56 1.84 17.995 1.84 17.995 2.875 17.765 2.875 17.765 1.615 15.99 1.615  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffnsnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 16.24 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.57 1.21 4.975 1.21 4.975 2.71 4.57 2.71  ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.77 1.59 1.77 1.59 2.15 0.65 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.835 2.33 15.095 2.33 15.47 2.33 15.47 0.55 15.85 0.55 15.85 2.975 15.095 2.975 14.835 2.975  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 3.305 3.62 3.305 3.185 3.535 3.185 3.535 3.62 6.59 3.62 7.63 3.62 7.63 2.7 7.97 2.7 7.97 3.62 8.41 3.62 11.33 3.62 12.625 3.62 12.625 2.635 12.855 2.635 12.855 3.62 13.35 3.62 14.365 3.62 14.365 2.635 14.595 2.635 14.595 3.62 15.095 3.62 16.24 3.62 16.24 4.22 15.095 4.22 13.35 4.22 11.33 4.22 8.41 4.22 6.59 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 16.24 -0.3 16.24 0.3 14.655 0.3 14.655 0.89 14.425 0.89 14.425 0.3 12.715 0.3 12.715 1.105 12.485 1.105 12.485 0.3 8.13 0.3 8.13 0.585 7.79 0.585 7.79 0.3 3.49 0.3 3.49 1.09 3.15 1.09 3.15 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.47 1.915 2.47 1.915 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.145 1.28 2.145 2.98 2.845 2.98 2.845 2.65 4.12 2.65 4.12 3.16 6.59 3.16 6.59 3.39 3.89 3.39 3.89 2.885 3.075 2.885 3.075 3.215 1.915 3.215 1.915 2.7 0.575 2.7 0.575 3.155 0.345 3.155  ;
        POLYGON 5.325 0.99 5.67 0.99 5.67 2.24 8.41 2.24 8.41 2.47 5.95 2.47 5.95 2.93 5.61 2.93 5.61 2.47 5.325 2.47  ;
        POLYGON 7.13 1.32 9.13 1.32 9.13 0.86 9.47 0.86 9.47 2.93 9.125 2.93 9.125 1.55 7.13 1.55  ;
        POLYGON 2.385 2.09 3.845 2.09 3.845 1.555 2.485 1.555 2.485 0.81 2.715 0.81 2.715 1.325 3.845 1.325 3.845 0.53 6.395 0.53 6.395 1.78 8.87 1.78 8.87 3.16 9.72 3.16 9.72 1.225 9.95 1.225 9.95 3.16 11.33 3.16 11.33 3.39 8.64 3.39 8.64 2.01 6.165 2.01 6.165 0.76 4.075 0.76 4.075 2.325 2.615 2.325 2.615 2.71 2.385 2.71  ;
        POLYGON 10.25 0.86 10.59 0.86 10.59 1.895 13.35 1.895 13.35 2.13 10.59 2.13 10.59 2.93 10.25 2.93  ;
        POLYGON 11.77 1.4 13.605 1.4 13.605 0.755 13.87 0.755 13.87 1.5 15.095 1.5 15.095 1.84 13.875 1.84 13.875 3.03 13.645 3.03 13.645 1.63 11.77 1.63  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.36 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.57 1.21 4.975 1.21 4.975 2.71 4.57 2.71  ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.77 1.59 1.77 1.59 2.15 0.65 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.33 2.33 15.565 2.33 16.03 2.33 16.03 1.02 15.45 1.02 15.45 0.55 16.41 0.55 16.41 2.975 15.565 2.975 15.33 2.975  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 3.305 3.62 3.305 3.185 3.535 3.185 3.535 3.62 6.59 3.62 7.63 3.62 7.63 2.7 7.97 2.7 7.97 3.62 8.41 3.62 11.33 3.62 12.625 3.62 12.625 2.635 12.855 2.635 12.855 3.62 13.35 3.62 14.365 3.62 14.365 2.635 14.595 2.635 14.595 3.62 15.565 3.62 16.665 3.62 16.665 2.635 16.895 2.635 16.895 3.62 17.36 3.62 17.36 4.22 15.565 4.22 13.35 4.22 11.33 4.22 8.41 4.22 6.59 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.36 -0.3 17.36 0.3 16.895 0.3 16.895 0.97 16.665 0.97 16.665 0.3 14.655 0.3 14.655 0.89 14.425 0.89 14.425 0.3 12.715 0.3 12.715 1.105 12.485 1.105 12.485 0.3 8.13 0.3 8.13 0.585 7.79 0.585 7.79 0.3 3.49 0.3 3.49 1.09 3.15 1.09 3.15 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.47 1.915 2.47 1.915 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.145 1.28 2.145 2.98 2.845 2.98 2.845 2.65 4.12 2.65 4.12 3.16 6.59 3.16 6.59 3.39 3.89 3.39 3.89 2.885 3.075 2.885 3.075 3.215 1.915 3.215 1.915 2.7 0.575 2.7 0.575 3.155 0.345 3.155  ;
        POLYGON 5.325 0.99 5.67 0.99 5.67 2.24 8.41 2.24 8.41 2.47 5.95 2.47 5.95 2.93 5.61 2.93 5.61 2.47 5.325 2.47  ;
        POLYGON 7.13 1.32 9.13 1.32 9.13 0.86 9.47 0.86 9.47 2.93 9.125 2.93 9.125 1.55 7.13 1.55  ;
        POLYGON 2.385 2.09 3.845 2.09 3.845 1.555 2.485 1.555 2.485 0.81 2.715 0.81 2.715 1.325 3.845 1.325 3.845 0.53 6.395 0.53 6.395 1.78 8.87 1.78 8.87 3.16 9.72 3.16 9.72 1.225 9.95 1.225 9.95 3.16 11.33 3.16 11.33 3.39 8.64 3.39 8.64 2.01 6.165 2.01 6.165 0.76 4.075 0.76 4.075 2.325 2.615 2.325 2.615 2.71 2.385 2.71  ;
        POLYGON 10.25 0.86 10.59 0.86 10.59 1.895 13.35 1.895 13.35 2.13 10.59 2.13 10.59 2.93 10.25 2.93  ;
        POLYGON 11.77 1.4 13.605 1.4 13.605 0.805 13.87 0.805 13.87 1.5 15.565 1.5 15.565 1.84 13.875 1.84 13.875 3.03 13.645 3.03 13.645 1.63 11.77 1.63  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.57 1.21 4.975 1.21 4.975 2.71 4.57 2.71  ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.59 1.77 1.59 2.13 0.28 2.13  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.6044 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.735 2.33 17.795 2.33 18.13 2.33 18.13 1.17 15.965 1.17 15.965 0.805 16.195 0.805 16.195 0.94 17.795 0.94 17.795 0.835 18.51 0.835 18.51 2.93 17.795 2.93 15.735 2.93  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 3.305 3.62 3.305 3.185 3.535 3.185 3.535 3.62 6.59 3.62 7.63 3.62 7.63 2.7 7.97 2.7 7.97 3.62 8.41 3.62 11.33 3.62 12.625 3.62 12.625 2.72 12.855 2.72 12.855 3.62 13.35 3.62 14.725 3.62 14.725 2.72 14.955 2.72 14.955 3.62 17.03 3.62 17.03 3.285 17.37 3.285 17.37 3.62 17.795 3.62 19.325 3.62 19.325 2.72 19.555 2.72 19.555 3.62 20.16 3.62 20.16 4.22 17.795 4.22 13.35 4.22 11.33 4.22 8.41 4.22 6.59 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 19.555 0.3 19.555 0.765 19.325 0.765 19.325 0.3 17.37 0.3 17.37 0.71 17.03 0.71 17.03 0.3 14.955 0.3 14.955 0.765 14.725 0.765 14.725 0.3 12.715 0.3 12.715 0.765 12.485 0.765 12.485 0.3 8.13 0.3 8.13 0.585 7.79 0.585 7.79 0.3 3.49 0.3 3.49 1.09 3.15 1.09 3.15 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.36 1.915 2.36 1.915 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.145 1.28 2.145 2.98 2.845 2.98 2.845 2.65 4.12 2.65 4.12 3.16 6.59 3.16 6.59 3.39 3.89 3.39 3.89 2.885 3.075 2.885 3.075 3.215 1.915 3.215 1.915 2.59 0.575 2.59 0.575 3.225 0.345 3.225  ;
        POLYGON 5.325 0.99 5.67 0.99 5.67 2.24 8.41 2.24 8.41 2.47 5.95 2.47 5.95 2.93 5.61 2.93 5.61 2.47 5.325 2.47  ;
        POLYGON 7.13 1.32 9.13 1.32 9.13 0.86 9.47 0.86 9.47 2.93 9.125 2.93 9.125 1.55 7.13 1.55  ;
        POLYGON 2.385 2.09 3.845 2.09 3.845 1.555 2.485 1.555 2.485 0.81 2.715 0.81 2.715 1.325 3.845 1.325 3.845 0.53 6.395 0.53 6.395 1.78 8.87 1.78 8.87 3.16 9.72 3.16 9.72 1.225 9.95 1.225 9.95 3.16 11.33 3.16 11.33 3.39 8.64 3.39 8.64 2.01 6.165 2.01 6.165 0.76 4.075 0.76 4.075 2.325 2.615 2.325 2.615 2.71 2.385 2.71  ;
        POLYGON 10.25 0.86 10.59 0.86 10.59 1.895 13.35 1.895 13.35 2.13 10.59 2.13 10.59 2.93 10.25 2.93  ;
        POLYGON 11.77 1.4 13.605 1.4 13.605 0.805 13.87 0.805 13.87 1.5 17.795 1.5 17.795 1.84 13.875 1.84 13.875 3.07 13.645 3.07 13.645 1.63 11.77 1.63  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.606 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 3.92 1.77 3.92 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.322 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.66 0.66 16.295 0.66 16.295 1.02 15.205 1.02 15.205 1.83 14.66 1.83  ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.57 1.77 1.57 2.15 0.28 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8932 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.475 0.55 18.91 0.55 18.91 3.38 18.475 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.865 1.65 2.865 1.65 3.62 2.035 3.62 3.05 3.62 3.05 2.845 3.39 2.845 3.39 3.62 4.915 3.62 7.35 3.62 7.35 2.99 7.69 2.99 7.69 3.62 8.995 3.62 9.485 3.62 9.485 2.79 9.715 2.79 9.715 3.62 10.155 3.62 11.08 3.62 14.655 3.62 14.655 3.28 14.995 3.28 14.995 3.62 16.42 3.62 16.75 3.62 16.75 2.59 16.98 2.59 16.98 3.62 17.47 3.62 17.47 2.53 17.7 2.53 17.7 3.62 18.23 3.62 19.04 3.62 19.04 4.22 18.23 4.22 16.42 4.22 11.08 4.22 10.155 4.22 8.995 4.22 4.915 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 17.655 0.3 17.655 0.875 17.315 0.875 17.315 0.3 14.3 0.3 14.3 1.13 14.07 1.13 14.07 0.3 8.77 0.3 8.77 0.915 8.43 0.915 8.43 0.3 3.51 0.3 3.51 1.075 3.17 1.075 3.17 0.3 1.655 0.3 1.655 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.405 1.805 2.405 1.805 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.035 1.28 2.035 2.635 0.575 2.635 0.575 3.225 0.345 3.225  ;
        POLYGON 4.125 2.42 4.225 2.42 4.225 0.845 4.63 0.845 4.63 1.075 4.455 1.075 4.455 2.76 4.125 2.76  ;
        POLYGON 2.495 2.385 3.895 2.385 3.895 2.99 4.685 2.99 4.685 1.91 4.915 1.91 4.915 3.22 3.665 3.22 3.665 2.615 2.615 2.615 2.615 3.215 2.265 3.215 2.265 0.865 2.77 0.865 2.77 1.095 2.495 1.095  ;
        POLYGON 6.165 2.53 8.995 2.53 8.995 3.13 8.765 3.13 8.765 2.76 6.395 2.76 6.395 2.955 6.165 2.955  ;
        POLYGON 5.145 2.07 5.465 2.07 5.465 0.79 5.695 0.79 5.695 2.07 10.155 2.07 10.155 2.525 9.855 2.525 9.855 2.3 5.375 2.3 5.375 2.76 5.145 2.76  ;
        POLYGON 6.69 1.61 9.99 1.61 9.99 1 10.33 1 10.33 1.61 10.67 1.61 10.67 2.845 11.08 2.845 11.08 3.075 10.44 3.075 10.44 1.84 6.69 1.84  ;
        POLYGON 6.045 1.15 9 1.15 9 0.53 12.35 0.53 12.35 1.36 13.12 1.36 13.12 2.525 12.89 2.525 12.89 1.59 12.12 1.59 12.12 0.76 11.155 0.76 11.155 1.59 10.925 1.59 10.925 0.76 9.23 0.76 9.23 1.38 6.275 1.38 6.275 1.59 6.045 1.59  ;
        POLYGON 12.95 0.79 13.755 0.79 13.755 2.93 13.415 2.93 13.415 1.13 12.95 1.13  ;
        POLYGON 11.55 1 11.89 1 11.89 1.82 12.44 1.82 12.44 3.16 14.195 3.16 14.195 2.82 15.465 2.82 15.465 3.16 16.19 3.16 16.19 1.91 16.42 1.91 16.42 3.39 15.235 3.39 15.235 3.05 14.425 3.05 14.425 3.39 12.21 3.39 12.21 2.05 11.55 2.05  ;
        POLYGON 13.995 2.175 15.73 2.175 15.73 1.45 16.65 1.45 16.65 0.79 16.88 0.79 16.88 1.45 18.23 1.45 18.23 1.68 15.96 1.68 15.96 2.93 15.73 2.93 15.73 2.405 13.995 2.405  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.606 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 3.92 1.77 3.92 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.4295 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.66 0.66 16.255 0.66 16.255 1.02 15.205 1.02 15.205 1.83 14.66 1.83  ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.57 1.77 1.57 2.15 0.28 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.475 2.05 18.69 2.05 19.14 2.05 19.14 1.27 18.475 1.27 18.475 0.55 18.94 0.55 18.94 1.04 19.5 1.04 19.5 2.28 18.94 2.28 18.94 3.38 18.69 3.38 18.475 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.865 1.65 2.865 1.65 3.62 2.035 3.62 3.05 3.62 3.05 2.845 3.39 2.845 3.39 3.62 4.915 3.62 7.35 3.62 7.35 2.99 7.69 2.99 7.69 3.62 8.995 3.62 9.485 3.62 9.485 2.79 9.715 2.79 9.715 3.62 10.155 3.62 11.08 3.62 14.655 3.62 14.655 3.28 14.995 3.28 14.995 3.62 16.42 3.62 16.75 3.62 16.75 2.57 16.985 2.57 16.985 3.62 17.465 3.62 17.465 2.57 17.7 2.57 17.7 3.62 18.69 3.62 19.455 3.62 19.455 2.53 19.795 2.53 19.795 3.62 20.16 3.62 20.16 4.22 18.69 4.22 16.42 4.22 11.08 4.22 10.155 4.22 8.995 4.22 4.915 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 19.895 0.3 19.895 0.79 19.555 0.79 19.555 0.3 17.655 0.3 17.655 0.79 17.315 0.79 17.315 0.3 14.3 0.3 14.3 1.13 14.07 1.13 14.07 0.3 8.77 0.3 8.77 0.915 8.43 0.915 8.43 0.3 3.51 0.3 3.51 1.075 3.17 1.075 3.17 0.3 1.655 0.3 1.655 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.405 1.805 2.405 1.805 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.035 1.28 2.035 2.635 0.575 2.635 0.575 3.225 0.345 3.225  ;
        POLYGON 4.125 2.42 4.225 2.42 4.225 0.845 4.63 0.845 4.63 1.075 4.455 1.075 4.455 2.76 4.125 2.76  ;
        POLYGON 2.495 2.385 3.895 2.385 3.895 2.99 4.685 2.99 4.685 1.91 4.915 1.91 4.915 3.22 3.665 3.22 3.665 2.615 2.615 2.615 2.615 3.215 2.265 3.215 2.265 0.865 2.77 0.865 2.77 1.095 2.495 1.095  ;
        POLYGON 6.165 2.53 8.995 2.53 8.995 3.13 8.765 3.13 8.765 2.76 6.395 2.76 6.395 2.955 6.165 2.955  ;
        POLYGON 5.145 2.07 5.465 2.07 5.465 0.79 5.695 0.79 5.695 2.07 10.155 2.07 10.155 2.525 9.855 2.525 9.855 2.3 5.375 2.3 5.375 2.76 5.145 2.76  ;
        POLYGON 6.69 1.61 9.99 1.61 9.99 1 10.33 1 10.33 1.61 10.67 1.61 10.67 2.845 11.08 2.845 11.08 3.075 10.44 3.075 10.44 1.84 6.69 1.84  ;
        POLYGON 6.045 1.15 9 1.15 9 0.53 12.35 0.53 12.35 1.36 13.12 1.36 13.12 2.525 12.89 2.525 12.89 1.59 12.12 1.59 12.12 0.76 11.155 0.76 11.155 1.59 10.925 1.59 10.925 0.76 9.23 0.76 9.23 1.38 6.275 1.38 6.275 1.59 6.045 1.59  ;
        POLYGON 12.95 0.79 13.755 0.79 13.755 2.93 13.415 2.93 13.415 1.13 12.95 1.13  ;
        POLYGON 11.55 1 11.89 1 11.89 1.82 12.44 1.82 12.44 3.16 14.195 3.16 14.195 2.82 15.465 2.82 15.465 3.16 16.19 3.16 16.19 1.91 16.42 1.91 16.42 3.39 15.235 3.39 15.235 3.05 14.425 3.05 14.425 3.39 12.21 3.39 12.21 2.05 11.55 2.05  ;
        POLYGON 13.995 2.175 15.73 2.175 15.73 1.45 16.65 1.45 16.65 0.81 16.88 0.81 16.88 1.525 18.69 1.525 18.69 1.755 16.65 1.755 16.65 1.68 15.96 1.68 15.96 2.93 15.73 2.93 15.73 2.405 13.995 2.405  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.606 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 3.92 1.77 3.92 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.4295 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.66 0.66 16.255 0.66 16.255 1.025 15.21 1.025 15.21 1.685 14.66 1.685  ;
    END
  END RN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.57 1.77 1.57 2.15 0.28 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1112 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.435 2.03 20.485 2.03 20.715 2.03 20.715 1.175 18.49 1.175 18.49 0.78 18.72 0.78 18.72 0.94 20.715 0.94 20.715 0.55 21.18 0.55 21.18 3.38 20.485 3.38 20.475 3.38 20.475 2.28 18.8 2.28 18.8 3.38 18.435 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.865 1.65 2.865 1.65 3.62 2.035 3.62 3.05 3.62 3.05 2.845 3.39 2.845 3.39 3.62 4.915 3.62 7.35 3.62 7.35 2.99 7.69 2.99 7.69 3.62 8.995 3.62 9.485 3.62 9.485 2.79 9.715 2.79 9.715 3.62 10.155 3.62 11.08 3.62 14.655 3.62 14.655 3.28 14.995 3.28 14.995 3.62 16.44 3.62 16.75 3.62 16.75 2.57 16.985 2.57 16.985 3.62 17.465 3.62 17.465 2.57 17.7 2.57 17.7 3.62 19.455 3.62 19.455 2.53 19.795 2.53 19.795 3.62 20.485 3.62 21.55 3.62 21.55 2.57 21.78 2.57 21.78 3.62 22.4 3.62 22.4 4.22 20.485 4.22 16.44 4.22 11.08 4.22 10.155 4.22 8.995 4.22 4.915 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 22.08 0.3 22.08 0.765 21.85 0.765 21.85 0.3 19.895 0.3 19.895 0.71 19.555 0.71 19.555 0.3 17.655 0.3 17.655 0.64 17.315 0.64 17.315 0.3 14.3 0.3 14.3 1.13 14.07 1.13 14.07 0.3 8.77 0.3 8.77 0.915 8.43 0.915 8.43 0.3 3.51 0.3 3.51 1.075 3.17 1.075 3.17 0.3 1.655 0.3 1.655 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.405 1.805 2.405 1.805 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.035 1.28 2.035 2.635 0.575 2.635 0.575 3.225 0.345 3.225  ;
        POLYGON 4.125 2.42 4.225 2.42 4.225 0.845 4.63 0.845 4.63 1.075 4.455 1.075 4.455 2.76 4.125 2.76  ;
        POLYGON 2.495 2.385 3.895 2.385 3.895 2.99 4.685 2.99 4.685 1.91 4.915 1.91 4.915 3.22 3.665 3.22 3.665 2.615 2.615 2.615 2.615 3.215 2.265 3.215 2.265 0.865 2.77 0.865 2.77 1.095 2.495 1.095  ;
        POLYGON 6.165 2.53 8.995 2.53 8.995 3.13 8.765 3.13 8.765 2.76 6.395 2.76 6.395 2.955 6.165 2.955  ;
        POLYGON 5.145 2.07 5.465 2.07 5.465 0.79 5.695 0.79 5.695 2.07 10.155 2.07 10.155 2.525 9.855 2.525 9.855 2.3 5.375 2.3 5.375 2.76 5.145 2.76  ;
        POLYGON 6.69 1.61 9.99 1.61 9.99 1 10.33 1 10.33 1.61 10.67 1.61 10.67 2.845 11.08 2.845 11.08 3.075 10.44 3.075 10.44 1.84 6.69 1.84  ;
        POLYGON 6.045 1.15 9 1.15 9 0.53 12.35 0.53 12.35 1.36 13.12 1.36 13.12 2.525 12.89 2.525 12.89 1.59 12.12 1.59 12.12 0.76 11.155 0.76 11.155 1.59 10.925 1.59 10.925 0.76 9.23 0.76 9.23 1.38 6.275 1.38 6.275 1.59 6.045 1.59  ;
        POLYGON 12.95 0.79 13.755 0.79 13.755 2.93 13.415 2.93 13.415 1.13 12.95 1.13  ;
        POLYGON 11.55 1 11.89 1 11.89 1.82 12.44 1.82 12.44 3.16 14.195 3.16 14.195 2.82 15.465 2.82 15.465 3.16 16.21 3.16 16.21 1.91 16.44 1.91 16.44 3.39 15.235 3.39 15.235 3.05 14.425 3.05 14.425 3.39 12.21 3.39 12.21 2.05 11.55 2.05  ;
        POLYGON 13.995 2.175 15.73 2.175 15.73 1.45 16.65 1.45 16.65 0.81 16.88 0.81 16.88 1.45 20.485 1.45 20.485 1.68 15.96 1.68 15.96 2.93 15.73 2.93 15.73 2.405 13.995 2.405  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.84 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4015 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 3.96 1.77 3.96 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.2095 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.715 1.785 18.115 1.785 18.115 2.15 16.715 2.15  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.65 1.7 15.955 1.7 15.955 2.15 14.65 2.15  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.575 1.77 1.575 2.13 0.28 2.13  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8932 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.825 0.86 21.335 0.86 21.335 3.38 20.825 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.205 3.62 1.205 2.93 1.555 2.93 1.555 3.62 2.055 3.62 3.01 3.62 3.01 3.005 3.35 3.005 3.35 3.62 5.095 3.62 7.53 3.62 7.53 3.445 7.87 3.445 7.87 3.62 10.73 3.62 10.73 3.445 11.07 3.445 11.07 3.62 12.75 3.62 15.125 3.62 15.125 2.93 15.465 2.93 15.465 3.62 17.27 3.62 17.27 2.93 17.61 2.93 17.61 3.62 19.035 3.62 19.365 3.62 19.365 2.81 19.595 2.81 19.595 3.62 20.085 3.62 20.085 2.53 20.315 2.53 20.315 3.62 20.595 3.62 21.84 3.62 21.84 4.22 20.595 4.22 19.035 4.22 12.75 4.22 5.095 4.22 2.055 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 21.84 -0.3 21.84 0.3 20.155 0.3 20.155 0.765 19.925 0.765 19.925 0.3 17.51 0.3 17.51 1.075 17.17 1.075 17.17 0.3 9.19 0.3 9.19 0.915 8.85 0.915 8.85 0.3 3.85 0.3 3.85 1.15 3.51 1.15 3.51 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.36 1.825 2.36 1.825 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.055 1.28 2.055 2.59 0.475 2.59 0.475 3.225 0.245 3.225  ;
        POLYGON 4.25 0.865 4.915 0.865 4.915 1.205 4.59 1.205 4.59 2.88 4.25 2.88  ;
        POLYGON 2.515 2.49 3.88 2.49 3.88 3.11 4.865 3.11 4.865 1.895 5.095 1.895 5.095 3.34 3.65 3.34 3.65 2.725 2.515 2.725 2.515 3.225 2.285 3.225 2.285 0.765 2.715 0.765 2.715 1.105 2.515 1.105  ;
        POLYGON 6.29 2.525 9.11 2.525 9.11 2.925 8.77 2.925 8.77 2.755 6.63 2.755 6.63 2.88 6.29 2.88  ;
        POLYGON 5.325 2.04 5.805 2.04 5.805 0.865 6.035 0.865 6.035 2.065 10.27 2.065 10.27 2.295 5.555 2.295 5.555 2.94 5.325 2.94  ;
        POLYGON 9.49 2.525 11.28 2.525 11.28 1.835 7.03 1.835 7.03 1.605 11.17 1.605 11.17 0.99 11.51 0.99 11.51 2.525 12.31 2.525 12.31 2.835 11.97 2.835 11.97 2.755 9.83 2.755 9.83 2.925 9.49 2.925  ;
        POLYGON 5.85 3.11 7.07 3.11 7.07 2.985 8.41 2.985 8.41 3.155 10.245 3.155 10.245 2.985 11.53 2.985 11.53 3.065 12.75 3.065 12.75 3.295 11.3 3.295 11.3 3.215 10.48 3.215 10.48 3.39 8.18 3.39 8.18 3.215 7.3 3.215 7.3 3.345 5.85 3.345  ;
        POLYGON 6.265 1.145 10.65 1.145 10.65 0.53 13.125 0.53 13.125 1.6 13.735 1.6 13.735 2.43 13.505 2.43 13.505 1.83 12.895 1.83 12.895 0.76 12 0.76 12 1.735 11.745 1.735 11.745 0.76 10.88 0.76 10.88 1.375 6.495 1.375 6.495 1.685 6.265 1.685  ;
        POLYGON 13.41 0.99 14.065 0.99 14.065 0.845 16.415 0.845 16.415 2.465 16.535 2.465 16.535 2.805 16.185 2.805 16.185 1.075 14.295 1.075 14.295 2.89 14.065 2.89 14.065 1.22 13.41 1.22  ;
        POLYGON 12.29 0.99 12.63 0.99 12.63 2.06 13.275 2.06 13.275 3.12 14.585 3.12 14.585 2.465 15.925 2.465 15.925 3.09 16.805 3.09 16.805 2.465 18.115 2.465 18.115 3.035 18.805 3.035 18.805 2.005 19.035 2.005 19.035 3.27 17.885 3.27 17.885 2.7 17.035 2.7 17.035 3.325 15.695 3.325 15.695 2.7 14.815 2.7 14.815 3.355 13.045 3.355 13.045 2.295 12.4 2.295 12.4 1.22 12.29 1.22  ;
        POLYGON 16.645 1.325 19.205 1.325 19.205 0.79 19.435 0.79 19.435 1.27 20.595 1.27 20.595 1.61 18.575 1.61 18.575 2.805 18.345 2.805 18.345 1.555 16.645 1.555  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrsnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.96 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4015 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 3.96 1.77 3.96 2.15 2.89 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.2095 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.715 1.785 18.115 1.785 18.115 2.15 16.715 2.15  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.65 1.7 15.955 1.7 15.955 2.15 14.65 2.15  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.31 1.77 1.575 1.77 1.575 2.13 0.31 2.13  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.1 2.33 21.12 2.33 21.37 2.33 21.37 1.09 20.99 1.09 20.99 0.86 21.755 0.86 21.755 3.38 21.12 3.38 21.1 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.205 3.62 1.205 2.93 1.555 2.93 1.555 3.62 2.055 3.62 3.01 3.62 3.01 3.005 3.35 3.005 3.35 3.62 5.095 3.62 7.53 3.62 7.53 3.445 7.87 3.445 7.87 3.62 10.73 3.62 10.73 3.445 11.07 3.445 11.07 3.62 12.75 3.62 15.125 3.62 15.125 2.93 15.465 2.93 15.465 3.62 17.27 3.62 17.27 2.93 17.61 2.93 17.61 3.62 19.035 3.62 19.365 3.62 19.365 2.81 19.595 2.81 19.595 3.62 20.085 3.62 20.085 2.57 20.315 2.57 20.315 3.62 21.12 3.62 22.125 3.62 22.125 2.57 22.355 2.57 22.355 3.62 22.96 3.62 22.96 4.22 21.12 4.22 19.035 4.22 12.75 4.22 5.095 4.22 2.055 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 22.96 -0.3 22.96 0.3 22.55 0.3 22.55 0.64 22.21 0.64 22.21 0.3 20.155 0.3 20.155 0.765 19.925 0.765 19.925 0.3 17.51 0.3 17.51 1.075 17.17 1.075 17.17 0.3 9.19 0.3 9.19 0.915 8.85 0.915 8.85 0.3 3.85 0.3 3.85 1.15 3.51 1.15 3.51 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.36 1.825 2.36 1.825 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.055 1.28 2.055 2.59 0.475 2.59 0.475 3.225 0.245 3.225  ;
        POLYGON 4.25 0.865 4.915 0.865 4.915 1.205 4.59 1.205 4.59 2.88 4.25 2.88  ;
        POLYGON 2.515 2.49 3.88 2.49 3.88 3.11 4.865 3.11 4.865 1.895 5.095 1.895 5.095 3.34 3.65 3.34 3.65 2.725 2.515 2.725 2.515 3.225 2.285 3.225 2.285 0.765 2.715 0.765 2.715 1.105 2.515 1.105  ;
        POLYGON 6.29 2.525 9.11 2.525 9.11 2.925 8.77 2.925 8.77 2.755 6.63 2.755 6.63 2.88 6.29 2.88  ;
        POLYGON 5.325 2.04 5.805 2.04 5.805 0.865 6.035 0.865 6.035 2.065 10.27 2.065 10.27 2.295 5.555 2.295 5.555 2.94 5.325 2.94  ;
        POLYGON 9.49 2.525 11.28 2.525 11.28 1.835 7.03 1.835 7.03 1.605 11.17 1.605 11.17 0.99 11.51 0.99 11.51 2.525 12.31 2.525 12.31 2.835 11.97 2.835 11.97 2.755 9.83 2.755 9.83 2.925 9.49 2.925  ;
        POLYGON 5.85 3.11 7.07 3.11 7.07 2.985 8.41 2.985 8.41 3.155 10.245 3.155 10.245 2.985 11.53 2.985 11.53 3.065 12.75 3.065 12.75 3.295 11.3 3.295 11.3 3.215 10.48 3.215 10.48 3.39 8.18 3.39 8.18 3.215 7.3 3.215 7.3 3.345 5.85 3.345  ;
        POLYGON 6.265 1.145 10.65 1.145 10.65 0.53 13.125 0.53 13.125 1.6 13.735 1.6 13.735 2.43 13.505 2.43 13.505 1.83 12.895 1.83 12.895 0.76 12 0.76 12 1.735 11.745 1.735 11.745 0.76 10.88 0.76 10.88 1.375 6.495 1.375 6.495 1.685 6.265 1.685  ;
        POLYGON 13.41 0.99 14.065 0.99 14.065 0.845 16.415 0.845 16.415 2.465 16.535 2.465 16.535 2.805 16.185 2.805 16.185 1.075 14.295 1.075 14.295 2.89 14.065 2.89 14.065 1.22 13.41 1.22  ;
        POLYGON 12.29 0.99 12.63 0.99 12.63 2.06 13.275 2.06 13.275 3.12 14.585 3.12 14.585 2.465 15.925 2.465 15.925 3.09 16.805 3.09 16.805 2.465 18.115 2.465 18.115 3.035 18.805 3.035 18.805 2.005 19.035 2.005 19.035 3.27 17.885 3.27 17.885 2.7 17.035 2.7 17.035 3.325 15.695 3.325 15.695 2.7 14.815 2.7 14.815 3.355 13.045 3.355 13.045 2.295 12.4 2.295 12.4 1.22 12.29 1.22  ;
        POLYGON 16.645 1.325 19.205 1.325 19.205 0.79 19.435 0.79 19.435 1.325 20.595 1.325 20.595 1.525 21.12 1.525 21.12 1.755 20.305 1.755 20.305 1.555 18.575 1.555 18.575 2.805 18.345 2.805 18.345 1.555 16.645 1.555  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrsnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 25.2 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4565 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.85 1.65 3.96 1.65 3.96 2.15 2.85 2.15  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.177 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.715 1.785 18.115 1.785 18.115 2.13 16.715 2.13  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.096 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.565 1.67 15.955 1.67 15.955 2.225 14.565 2.225  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.6 1.07 0.6 1.07 2.15 0.705 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1112 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.045 2.125 22.89 2.125 23.14 2.125 23.14 1.315 21.045 1.315 21.045 0.655 21.275 0.655 21.275 1.085 23.14 1.085 23.14 0.6 24.005 0.6 24.005 2.28 23.42 2.28 23.42 3.38 23.06 3.38 23.06 2.36 22.89 2.36 21.335 2.36 21.335 3.38 21.045 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.205 3.62 1.205 2.93 1.555 2.93 1.555 3.62 2.035 3.62 3.01 3.62 3.01 3.005 3.35 3.005 3.35 3.62 4.995 3.62 7.53 3.62 7.53 3.445 7.87 3.445 7.87 3.62 10.73 3.62 10.73 3.445 11.07 3.445 11.07 3.62 12.75 3.62 15.125 3.62 15.125 2.93 15.465 2.93 15.465 3.62 17.27 3.62 17.27 2.93 17.61 2.93 17.61 3.62 19.035 3.62 19.365 3.62 19.365 2.73 19.595 2.73 19.595 3.62 20.085 3.62 20.085 2.53 20.315 2.53 20.315 3.62 22.07 3.62 22.07 2.62 22.41 2.62 22.41 3.62 22.89 3.62 24.165 3.62 24.165 2.53 24.395 2.53 24.395 3.62 25.2 3.62 25.2 4.22 22.89 4.22 19.035 4.22 12.75 4.22 4.995 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 25.2 -0.3 25.2 0.3 24.635 0.3 24.635 0.905 24.405 0.905 24.405 0.3 22.395 0.3 22.395 0.765 22.165 0.765 22.165 0.3 20.155 0.3 20.155 0.905 19.925 0.905 19.925 0.3 17.51 0.3 17.51 1.075 17.17 1.075 17.17 0.3 9.19 0.3 9.19 0.915 8.85 0.915 8.85 0.3 3.85 0.3 3.85 1.15 3.51 1.15 3.51 0.3 1.595 0.3 1.595 1.16 1.365 1.16 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.81 0.475 0.81 0.475 2.38 1.805 2.38 1.805 1.28 2.035 1.28 2.035 2.7 0.475 2.7 0.475 3.225 0.245 3.225  ;
        POLYGON 4.305 0.865 4.915 0.865 4.915 1.205 4.535 1.205 4.535 2.93 4.305 2.93  ;
        POLYGON 2.515 2.49 3.88 2.49 3.88 3.16 4.765 3.16 4.765 1.895 4.995 1.895 4.995 3.39 3.65 3.39 3.65 2.725 2.515 2.725 2.515 3.225 2.285 3.225 2.285 0.765 2.715 0.765 2.715 1.105 2.515 1.105  ;
        POLYGON 6.29 2.525 9.11 2.525 9.11 2.93 8.77 2.93 8.77 2.755 6.63 2.755 6.63 2.885 6.29 2.885  ;
        POLYGON 5.325 2.04 5.805 2.04 5.805 0.865 6.035 0.865 6.035 2.065 10.36 2.065 10.36 2.295 5.555 2.295 5.555 2.94 5.325 2.94  ;
        POLYGON 9.49 2.525 11.28 2.525 11.28 1.835 7.03 1.835 7.03 1.605 11.17 1.605 11.17 0.99 11.51 0.99 11.51 2.525 12.31 2.525 12.31 2.835 11.97 2.835 11.97 2.755 9.83 2.755 9.83 2.93 9.49 2.93  ;
        POLYGON 5.78 3.16 7.07 3.16 7.07 2.985 8.41 2.985 8.41 3.16 10.245 3.16 10.245 2.985 11.53 2.985 11.53 3.065 12.75 3.065 12.75 3.295 11.3 3.295 11.3 3.215 10.48 3.215 10.48 3.39 8.18 3.39 8.18 3.215 7.3 3.215 7.3 3.39 5.78 3.39  ;
        POLYGON 6.265 1.145 10.65 1.145 10.65 0.53 13.125 0.53 13.125 1.6 13.735 1.6 13.735 2.43 13.505 2.43 13.505 1.83 12.895 1.83 12.895 0.76 12 0.76 12 1.735 11.745 1.735 11.745 0.76 10.88 0.76 10.88 1.375 6.495 1.375 6.495 1.685 6.265 1.685  ;
        POLYGON 13.41 0.99 14.065 0.99 14.065 0.845 16.415 0.845 16.415 2.465 16.535 2.465 16.535 2.805 16.185 2.805 16.185 1.075 14.295 1.075 14.295 2.89 14.065 2.89 14.065 1.22 13.41 1.22  ;
        POLYGON 12.29 0.99 12.63 0.99 12.63 2.06 13.275 2.06 13.275 3.12 14.585 3.12 14.585 2.465 15.925 2.465 15.925 3.09 16.805 3.09 16.805 2.465 18.115 2.465 18.115 3.035 18.805 3.035 18.805 2.005 19.035 2.005 19.035 3.27 17.885 3.27 17.885 2.7 17.035 2.7 17.035 3.325 15.695 3.325 15.695 2.7 14.815 2.7 14.815 3.355 13.045 3.355 13.045 2.295 12.4 2.295 12.4 1.22 12.29 1.22  ;
        POLYGON 16.645 1.325 19.205 1.325 19.205 0.79 19.435 0.79 19.435 1.325 20.595 1.325 20.595 1.555 22.89 1.555 22.89 1.785 20.305 1.785 20.305 1.555 18.575 1.555 18.575 2.805 18.345 2.805 18.345 1.555 16.645 1.555  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffrsnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4685 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 4.03 1.77 4.03 2.15 2.89 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.09 1.77 15.285 1.77 15.285 2.15 14.09 2.15  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.765 1.59 1.765 1.59 2.13 0.28 2.13  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0147 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.045 2.19 19.12 2.19 19.425 2.19 19.425 1.16 19.3 1.16 19.3 0.55 19.815 0.55 19.815 3.38 19.12 3.38 19.045 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 2.09 3.62 3.24 3.62 3.24 2.845 3.58 2.845 3.58 3.62 5.115 3.62 7.675 3.62 7.675 3.445 8.015 3.445 8.015 3.62 10.275 3.62 10.275 3.005 10.615 3.005 10.615 3.62 12.315 3.62 14.295 3.62 14.295 3.005 14.635 3.005 14.635 3.62 15.6 3.62 16.71 3.62 16.71 2.53 16.94 2.53 16.94 3.62 18.45 3.62 18.45 2.53 18.68 2.53 18.68 3.62 19.12 3.62 20.16 3.62 20.16 4.22 19.12 4.22 15.6 4.22 12.315 4.22 5.115 4.22 2.09 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 18.68 0.3 18.68 0.765 18.45 0.765 18.45 0.3 16.895 0.3 16.895 1.05 16.555 1.05 16.555 0.3 7.795 0.3 7.795 1.075 7.455 1.075 7.455 0.3 3.49 0.3 3.49 1.075 3.15 1.075 3.15 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.36 1.86 2.36 1.86 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.09 1.28 2.09 2.595 0.575 2.595 0.575 3.225 0.345 3.225  ;
        POLYGON 4.27 0.79 4.61 0.79 4.61 2.93 4.27 2.93  ;
        POLYGON 2.62 2.38 4.04 2.38 4.04 3.16 4.885 3.16 4.885 1.93 5.115 1.93 5.115 3.39 3.81 3.39 3.81 2.615 2.615 2.615 2.615 3.225 2.385 3.225 2.385 0.81 2.715 0.81 2.715 1.15 2.62 1.15  ;
        POLYGON 5.345 0.79 5.675 0.79 5.675 1.765 8.235 1.765 8.235 1.995 5.575 1.995 5.575 2.985 5.345 2.985  ;
        POLYGON 6 1.305 8.11 1.305 8.11 0.53 11.04 0.53 11.04 1.615 10.81 1.615 10.81 0.76 8.34 0.76 8.34 1.535 6 1.535  ;
        POLYGON 7.015 2.225 9.035 2.225 9.035 2.08 9.875 2.08 9.875 0.99 10.215 0.99 10.215 2.08 11.645 2.08 11.645 2.78 11.305 2.78 11.305 2.31 9.375 2.31 9.375 2.93 9.035 2.93 9.035 2.455 7.015 2.455  ;
        POLYGON 6.115 2.24 6.455 2.24 6.455 2.985 8.5 2.985 8.5 3.16 9.685 3.16 9.685 2.54 11.075 2.54 11.075 3.065 12.315 3.065 12.315 3.295 10.845 3.295 10.845 2.775 9.915 2.775 9.915 3.39 8.27 3.39 8.27 3.215 6.115 3.215  ;
        POLYGON 13.86 2.54 15.6 2.54 15.6 2.885 15.37 2.885 15.37 2.775 13.86 2.775 13.86 2.845 13.63 2.845 13.63 1.22 12.555 1.22 12.555 0.99 14.495 0.99 14.495 1.22 13.86 1.22  ;
        POLYGON 11.27 0.79 11.93 0.79 11.93 0.53 16.11 0.53 16.11 1.395 17.335 1.395 17.335 1.63 15.88 1.63 15.88 0.76 12.16 0.76 12.16 2.55 12.895 2.55 12.895 2.78 11.93 2.78 11.93 1.13 11.27 1.13  ;
        POLYGON 15.755 1.86 17.73 1.86 17.73 0.805 17.96 0.805 17.96 1.5 19.12 1.5 19.12 1.84 17.96 1.84 17.96 3.38 17.73 3.38 17.73 2.105 15.755 2.105  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffsnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4685 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 4.03 1.77 4.03 2.15 2.89 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.09 1.77 15.285 1.77 15.285 2.15 14.09 2.15  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.765 1.59 1.765 1.59 2.13 0.65 2.13  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.2986 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.53 2.33 19.69 2.33 19.95 2.33 19.95 1.02 19.33 1.02 19.33 0.55 20.37 0.55 20.37 3.38 19.69 3.38 19.53 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 2.09 3.62 3.24 3.62 3.24 2.845 3.58 2.845 3.58 3.62 5.115 3.62 7.675 3.62 7.675 3.445 8.015 3.445 8.015 3.62 10.275 3.62 10.275 3.005 10.615 3.005 10.615 3.62 12.315 3.62 14.295 3.62 14.295 3.005 14.635 3.005 14.635 3.62 15.6 3.62 16.81 3.62 16.81 2.53 17.04 2.53 17.04 3.62 18.55 3.62 18.55 2.53 18.78 2.53 18.78 3.62 19.69 3.62 20.79 3.62 20.79 2.53 21.02 2.53 21.02 3.62 21.28 3.62 21.28 4.22 19.69 4.22 15.6 4.22 12.315 4.22 5.115 4.22 2.09 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 21.02 0.3 21.02 0.89 20.79 0.89 20.79 0.3 18.78 0.3 18.78 0.89 18.55 0.89 18.55 0.3 16.895 0.3 16.895 0.835 16.555 0.835 16.555 0.3 7.795 0.3 7.795 1.075 7.455 1.075 7.455 0.3 3.49 0.3 3.49 1.075 3.15 1.075 3.15 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.36 1.86 2.36 1.86 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.09 1.28 2.09 2.595 0.575 2.595 0.575 3.225 0.345 3.225  ;
        POLYGON 4.27 0.79 4.61 0.79 4.61 2.93 4.27 2.93  ;
        POLYGON 2.62 2.38 4.04 2.38 4.04 3.16 4.885 3.16 4.885 1.93 5.115 1.93 5.115 3.39 3.81 3.39 3.81 2.615 2.615 2.615 2.615 3.225 2.385 3.225 2.385 0.81 2.715 0.81 2.715 1.15 2.62 1.15  ;
        POLYGON 5.345 0.79 5.675 0.79 5.675 1.765 8.235 1.765 8.235 1.995 5.575 1.995 5.575 2.985 5.345 2.985  ;
        POLYGON 6 1.305 8.11 1.305 8.11 0.53 11.04 0.53 11.04 1.615 10.81 1.615 10.81 0.76 8.34 0.76 8.34 1.535 6 1.535  ;
        POLYGON 7.015 2.225 9.035 2.225 9.035 2.08 9.875 2.08 9.875 0.99 10.215 0.99 10.215 2.08 11.645 2.08 11.645 2.78 11.305 2.78 11.305 2.31 9.375 2.31 9.375 2.93 9.035 2.93 9.035 2.455 7.015 2.455  ;
        POLYGON 6.115 2.24 6.455 2.24 6.455 2.985 8.5 2.985 8.5 3.16 9.685 3.16 9.685 2.54 11.075 2.54 11.075 3.065 12.315 3.065 12.315 3.295 10.845 3.295 10.845 2.775 9.915 2.775 9.915 3.39 8.27 3.39 8.27 3.215 6.115 3.215  ;
        POLYGON 13.86 2.54 15.6 2.54 15.6 2.885 15.37 2.885 15.37 2.775 13.86 2.775 13.86 2.845 13.63 2.845 13.63 1.22 12.555 1.22 12.555 0.99 14.495 0.99 14.495 1.22 13.86 1.22  ;
        POLYGON 11.27 0.79 11.93 0.79 11.93 0.53 16.11 0.53 16.11 1.395 17.335 1.395 17.335 1.63 15.88 1.63 15.88 0.76 12.16 0.76 12.16 2.55 12.895 2.55 12.895 2.78 11.93 2.78 11.93 1.13 11.27 1.13  ;
        POLYGON 15.755 1.86 17.73 1.86 17.73 0.55 17.96 0.55 17.96 1.5 19.69 1.5 19.69 1.84 18.06 1.84 18.06 3.38 17.83 3.38 17.83 2.105 15.755 2.105  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffsnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dffsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 24.08 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4685 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.77 4.03 1.77 4.03 2.15 2.89 2.15  ;
    END
  END D
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.1415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.09 1.77 15.285 1.77 15.285 2.15 14.09 2.15  ;
    END
  END SETN
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6755 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.765 1.59 1.765 1.59 2.13 0.28 2.13  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.5972 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.05 2.06 21.605 2.06 22.01 2.06 22.01 1.315 20.045 1.315 20.045 0.55 20.28 0.55 20.28 1.085 22.01 1.085 22.01 0.55 22.535 0.55 22.535 3.38 21.67 3.38 21.67 2.29 21.605 2.29 20.28 2.29 20.28 3.38 20.05 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.31 3.62 1.31 2.93 1.65 2.93 1.65 3.62 2.09 3.62 3.24 3.62 3.24 2.845 3.58 2.845 3.58 3.62 5.115 3.62 7.675 3.62 7.675 3.445 8.015 3.445 8.015 3.62 10.275 3.62 10.275 3.005 10.615 3.005 10.615 3.62 12.315 3.62 14.295 3.62 14.295 3.005 14.635 3.005 14.635 3.62 15.6 3.62 16.705 3.62 16.705 2.53 16.935 2.53 16.935 3.62 18.75 3.62 18.75 2.53 18.98 2.53 18.98 3.62 21.17 3.62 21.17 2.53 21.4 2.53 21.4 3.62 21.605 3.62 23.41 3.62 23.41 2.53 23.64 2.53 23.64 3.62 24.08 3.62 24.08 4.22 21.605 4.22 15.6 4.22 12.315 4.22 5.115 4.22 2.09 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 24.08 -0.3 24.08 0.3 23.64 0.3 23.64 0.89 23.41 0.89 23.41 0.3 21.455 0.3 21.455 0.835 21.115 0.835 21.115 0.3 19.08 0.3 19.08 0.89 18.85 0.89 18.85 0.3 16.895 0.3 16.895 0.835 16.555 0.835 16.555 0.3 7.795 0.3 7.795 1.075 7.455 1.075 7.455 0.3 3.49 0.3 3.49 1.075 3.15 1.075 3.15 0.3 1.65 0.3 1.65 1.05 1.31 1.05 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.36 1.86 2.36 1.86 1.51 0.245 1.51 0.245 0.81 0.475 0.81 0.475 1.28 2.09 1.28 2.09 2.595 0.575 2.595 0.575 3.225 0.345 3.225  ;
        POLYGON 4.27 0.79 4.61 0.79 4.61 2.93 4.27 2.93  ;
        POLYGON 2.62 2.38 4.04 2.38 4.04 3.16 4.885 3.16 4.885 1.93 5.115 1.93 5.115 3.39 3.81 3.39 3.81 2.615 2.615 2.615 2.615 3.225 2.385 3.225 2.385 0.81 2.715 0.81 2.715 1.15 2.62 1.15  ;
        POLYGON 5.345 0.79 5.675 0.79 5.675 1.765 8.235 1.765 8.235 1.995 5.575 1.995 5.575 2.985 5.345 2.985  ;
        POLYGON 6 1.305 8.11 1.305 8.11 0.53 11.04 0.53 11.04 1.615 10.81 1.615 10.81 0.76 8.34 0.76 8.34 1.535 6 1.535  ;
        POLYGON 7.015 2.225 9.035 2.225 9.035 2.08 9.875 2.08 9.875 0.99 10.215 0.99 10.215 2.08 11.645 2.08 11.645 2.78 11.305 2.78 11.305 2.31 9.375 2.31 9.375 2.93 9.035 2.93 9.035 2.455 7.015 2.455  ;
        POLYGON 6.115 2.24 6.455 2.24 6.455 2.985 8.5 2.985 8.5 3.16 9.685 3.16 9.685 2.54 11.075 2.54 11.075 3.065 12.315 3.065 12.315 3.295 10.845 3.295 10.845 2.775 9.915 2.775 9.915 3.39 8.27 3.39 8.27 3.215 6.115 3.215  ;
        POLYGON 13.86 2.54 15.6 2.54 15.6 2.885 15.37 2.885 15.37 2.775 13.86 2.775 13.86 2.845 13.63 2.845 13.63 1.22 12.555 1.22 12.555 0.99 14.495 0.99 14.495 1.22 13.86 1.22  ;
        POLYGON 11.27 0.79 11.93 0.79 11.93 0.53 16.11 0.53 16.11 1.395 17.335 1.395 17.335 1.63 15.88 1.63 15.88 0.76 12.16 0.76 12.16 2.55 12.895 2.55 12.895 2.78 11.93 2.78 11.93 1.13 11.27 1.13  ;
        POLYGON 15.755 1.86 17.73 1.86 17.73 0.55 17.96 0.55 17.96 1.555 21.605 1.555 21.605 1.785 17.96 1.785 17.96 3.38 17.73 3.38 17.73 2.105 15.755 2.105  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dffsnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlya_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlya_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.16 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.21 1.845 1.21 1.845 1.61 0.705 1.61  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.65 0.55 6.02 0.55 6.02 3.38 5.65 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.21 3.62 1.21 2.54 1.55 2.54 1.55 3.62 2.135 3.62 4.645 3.62 4.645 2.53 4.875 2.53 4.875 3.62 5.215 3.62 6.16 3.62 6.16 4.22 5.215 4.22 2.135 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.16 -0.3 6.16 0.3 4.775 0.3 4.775 0.69 4.545 0.69 4.545 0.3 1.595 0.3 1.595 0.98 1.365 0.98 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.64 0.475 0.64 0.475 2.025 2.135 2.025 2.135 2.255 0.475 2.255 0.475 2.825 0.245 2.825  ;
        POLYGON 2.385 0.64 2.715 0.64 2.715 1.495 4.18 1.495 4.18 1.725 2.615 1.725 2.615 2.825 2.385 2.825  ;
        POLYGON 3.105 2.05 4.985 2.05 4.985 1.18 3.87 1.18 3.87 0.765 3.145 0.765 3.145 0.53 4.105 0.53 4.105 0.95 5.215 0.95 5.215 2.28 3.335 2.28 3.335 2.71 3.105 2.71  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlya_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlya_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlya_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.28 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.21 1.59 1.21 1.59 1.61 0.705 1.61  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1889 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.66 0.805 6.07 0.805 6.07 3.38 5.66 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.21 3.62 1.21 2.54 1.55 2.54 1.55 3.62 2.035 3.62 4.64 3.62 4.64 2.53 4.87 2.53 4.87 3.62 5.375 3.62 6.785 3.62 6.785 2.53 7.02 2.53 7.02 3.62 7.28 3.62 7.28 4.22 5.375 4.22 2.035 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.28 -0.3 7.28 0.3 7.015 0.3 7.015 1.145 6.785 1.145 6.785 0.3 4.775 0.3 4.775 0.69 4.545 0.69 4.545 0.3 1.595 0.3 1.595 0.98 1.365 0.98 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.64 0.475 0.64 0.475 2.075 1.805 2.075 1.805 1.97 2.035 1.97 2.035 2.31 0.475 2.31 0.475 2.825 0.245 2.825  ;
        POLYGON 2.385 0.64 2.715 0.64 2.715 1.55 4.055 1.55 4.055 1.79 2.615 1.79 2.615 2.825 2.385 2.825  ;
        POLYGON 3.105 2.05 5.145 2.05 5.145 1.25 4.05 1.25 4.05 0.765 3.145 0.765 3.145 0.53 4.285 0.53 4.285 1.02 5.375 1.02 5.375 2.28 3.335 2.28 3.335 2.71 3.105 2.71  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlya_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlya_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlya_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 9.52 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.21 2.15 1.21 2.15 1.59 0.71 1.59  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3656 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.68 2.35 7.06 2.35 7.82 2.35 7.82 1.405 5.63 1.405 5.63 0.6 5.86 0.6 5.86 1.17 7.87 1.17 7.87 0.6 8.39 0.6 8.39 3.16 7.82 3.16 7.82 2.58 7.06 2.58 5.91 2.58 5.91 3.16 5.68 3.16  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.27 3.62 1.27 2.635 1.5 2.635 1.5 3.62 2.095 3.62 4.455 3.62 4.455 2.66 4.795 2.66 4.795 3.62 6.645 3.62 6.645 2.81 6.985 2.81 6.985 3.62 7.06 3.62 8.89 3.62 8.89 2.605 9.12 2.605 9.12 3.62 9.52 3.62 9.52 4.22 7.06 4.22 2.095 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 9.52 -0.3 9.52 0.3 9.22 0.3 9.22 0.94 8.99 0.94 8.99 0.3 6.98 0.3 6.98 0.94 6.75 0.94 6.75 0.3 4.56 0.3 4.56 0.905 4.33 0.905 4.33 0.3 1.655 0.3 1.655 0.845 1.315 0.845 1.315 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.25 0.56 0.48 0.56 0.48 2.175 2.095 2.175 2.095 2.405 0.48 2.405 0.48 2.98 0.25 2.98  ;
        POLYGON 2.39 2.64 2.49 2.64 2.49 0.56 2.72 0.56 2.72 1.6 3.985 1.6 3.985 1.83 2.72 1.83 2.72 2.98 2.39 2.98  ;
        POLYGON 3.26 2.06 4.215 2.06 4.215 1.37 3.21 1.37 3.21 0.56 3.44 0.56 3.44 1.135 4.445 1.135 4.445 1.685 7.06 1.685 7.06 2.025 4.445 2.025 4.445 2.295 3.49 2.295 3.49 2.98 3.26 2.98  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlya_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlyb_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyb_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.96 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.93 1.2 3.355 1.2 3.355 1.6 0.93 1.6  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.81 2.33 7.975 2.33 8.37 2.33 8.37 0.675 8.6 0.675 8.6 3.195 8.215 3.195 8.215 2.71 7.975 2.71 6.81 2.71  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.485 3.62 1.485 3.285 1.825 3.285 1.825 3.62 3.265 3.62 6.565 3.62 6.565 3.175 6.905 3.175 6.905 3.62 7.975 3.62 8.96 3.62 8.96 4.22 7.975 4.22 3.265 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.96 -0.3 8.96 0.3 6.95 0.3 6.95 0.69 6.72 0.69 6.72 0.3 1.925 0.3 1.925 0.635 1.585 0.635 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.065 3.265 2.065 3.265 2.405 0.585 2.405 0.585 3.105 0.245 3.105 0.245 0.67 0.585 0.67 0.585 0.9 0.475 0.9  ;
        POLYGON 3.72 0.77 4.105 0.77 4.105 1.68 5.485 1.68 5.485 1.91 3.95 1.91 3.95 3.16 3.72 3.16  ;
        POLYGON 4.54 2.235 5.835 2.235 5.835 1.055 4.54 1.055 4.54 0.715 6.155 0.715 6.155 1.395 7.975 1.395 7.975 1.625 6.155 1.625 6.155 2.465 4.77 2.465 4.77 3.16 4.54 3.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyb_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlyb_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyb_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.93 1.2 3.355 1.2 3.355 1.6 0.93 1.6  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.42 2.105 8.54 2.105 8.93 2.105 8.93 1.215 8.37 1.215 8.37 0.53 8.6 0.53 8.6 0.96 9.38 0.96 9.38 2.34 8.86 2.34 8.86 3.39 8.54 3.39 8.42 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.485 3.62 1.485 3.285 1.825 3.285 1.825 3.62 3.265 3.62 6.565 3.62 6.565 3.175 7.345 3.175 7.345 2.53 7.685 2.53 7.685 3.62 8.54 3.62 9.435 3.62 9.435 2.57 9.775 2.57 9.775 3.62 10.08 3.62 10.08 4.22 8.54 4.22 3.265 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.775 0.3 9.775 0.635 9.435 0.635 9.435 0.3 6.95 0.3 6.95 0.69 6.72 0.69 6.72 0.3 1.925 0.3 1.925 0.635 1.585 0.635 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.065 3.265 2.065 3.265 2.405 0.585 2.405 0.585 3.105 0.245 3.105 0.245 0.67 0.585 0.67 0.585 0.9 0.475 0.9  ;
        POLYGON 3.72 0.77 4.105 0.77 4.105 1.68 5.485 1.68 5.485 1.91 3.95 1.91 3.95 3.16 3.72 3.16  ;
        POLYGON 4.54 2.235 5.835 2.235 5.835 1.055 4.54 1.055 4.54 0.715 6.155 0.715 6.155 1.625 8.54 1.625 8.54 1.855 6.155 1.855 6.155 2.465 4.77 2.465 4.77 3.16 4.54 3.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyb_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlyb_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyb_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.93 1.2 3.36 1.2 3.36 1.6 0.93 1.6  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3046 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.42 2.105 10.36 2.105 10.61 2.105 10.61 1.215 8.37 1.215 8.37 0.53 8.6 0.53 8.6 0.96 10.61 0.96 10.61 0.55 11.18 0.55 11.18 3.38 10.61 3.38 10.61 2.34 10.36 2.34 8.65 2.34 8.65 3.38 8.42 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.485 3.62 1.485 3.285 1.825 3.285 1.825 3.62 3.265 3.62 6.565 3.62 6.565 3.175 7.355 3.175 7.355 2.53 7.685 2.53 7.685 3.62 9.44 3.62 9.44 2.57 9.67 2.57 9.67 3.62 10.36 3.62 11.63 3.62 11.63 2.53 11.86 2.53 11.86 3.62 12.32 3.62 12.32 4.22 10.36 4.22 3.265 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 11.96 0.3 11.96 1.115 11.73 1.115 11.73 0.3 9.775 0.3 9.775 0.635 9.435 0.635 9.435 0.3 6.95 0.3 6.95 0.69 6.72 0.69 6.72 0.3 1.925 0.3 1.925 0.635 1.585 0.635 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.065 3.265 2.065 3.265 2.405 0.585 2.405 0.585 3.105 0.245 3.105 0.245 0.67 0.585 0.67 0.585 0.9 0.475 0.9  ;
        POLYGON 3.72 0.77 4.105 0.77 4.105 1.68 5.485 1.68 5.485 1.91 3.95 1.91 3.95 3.16 3.72 3.16  ;
        POLYGON 4.54 2.235 5.835 2.235 5.835 1.055 4.54 1.055 4.54 0.715 6.155 0.715 6.155 1.625 10.36 1.625 10.36 1.855 6.155 1.855 6.155 2.465 4.77 2.465 4.77 3.16 4.54 3.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyb_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlyc_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyc_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.905 1.2 3.33 1.2 3.33 1.6 0.905 1.6  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.965 2.33 13.13 2.33 13.525 2.33 13.525 0.675 13.755 0.675 13.755 3.195 13.37 3.195 13.37 2.71 13.13 2.71 11.965 2.71  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.46 3.62 1.46 3.285 1.8 3.285 1.8 3.62 3.24 3.62 6.44 3.62 6.44 3.285 6.78 3.285 6.78 3.62 8.09 3.62 11.72 3.62 11.72 3.175 12.06 3.175 12.06 3.62 13.13 3.62 14 3.62 14 4.22 13.13 4.22 8.09 4.22 3.24 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14 -0.3 14 0.3 12.345 0.3 12.345 0.69 12.115 0.69 12.115 0.3 6.98 0.3 6.98 0.635 6.64 0.635 6.64 0.3 1.9 0.3 1.9 0.635 1.56 0.635 1.56 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.22 0.67 0.56 0.67 0.56 2.065 3.24 2.065 3.24 2.405 0.56 2.405 0.56 3.105 0.22 3.105  ;
        POLYGON 3.695 0.77 4.08 0.77 4.08 1.465 5.305 1.465 5.305 1.805 3.925 1.805 3.925 3.16 3.695 3.16  ;
        POLYGON 4.36 2.875 5.535 2.875 5.535 1 4.46 1 4.46 0.77 5.765 0.77 5.765 1.52 8.09 1.52 8.09 1.75 5.765 1.75 5.765 3.105 4.36 3.105  ;
        POLYGON 8.875 0.715 9.105 0.715 9.105 1.535 11.055 1.535 11.055 1.965 9.26 1.965 9.26 3.16 8.875 3.16  ;
        POLYGON 9.695 2.235 11.345 2.235 11.345 1.055 9.695 1.055 9.695 0.715 11.665 0.715 11.665 1.395 13.13 1.395 13.13 1.625 11.665 1.625 11.665 2.465 9.925 2.465 9.925 3.16 9.695 3.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyc_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlyc_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyc_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.12 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.93 1.2 3.35 1.2 3.35 1.6 0.93 1.6  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.2817 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.395 0.675 13.91 0.675 13.91 3.195 13.395 3.195  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.485 3.62 1.485 3.285 1.825 3.285 1.825 3.62 3.265 3.62 6.465 3.62 6.465 3.285 6.805 3.285 6.805 3.62 8.115 3.62 11.745 3.62 11.745 3.175 12.085 3.175 12.085 3.62 12.81 3.62 14.465 3.62 14.465 2.705 14.805 2.705 14.805 3.62 15.12 3.62 15.12 4.22 12.81 4.22 8.115 4.22 3.265 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 15.12 -0.3 15.12 0.3 14.75 0.3 14.75 0.69 14.52 0.69 14.52 0.3 12.155 0.3 12.155 0.69 11.925 0.69 11.925 0.3 7.005 0.3 7.005 0.635 6.665 0.635 6.665 0.3 1.925 0.3 1.925 0.635 1.585 0.635 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.065 3.265 2.065 3.265 2.405 0.585 2.405 0.585 3.105 0.245 3.105 0.245 0.67 0.585 0.67 0.585 0.9 0.475 0.9  ;
        POLYGON 3.72 0.77 4.105 0.77 4.105 1.465 5.33 1.465 5.33 1.805 3.95 1.805 3.95 3.16 3.72 3.16  ;
        POLYGON 4.385 2.875 5.56 2.875 5.56 1 4.485 1 4.485 0.77 5.79 0.77 5.79 1.52 8.115 1.52 8.115 1.75 5.79 1.75 5.79 3.105 4.385 3.105  ;
        POLYGON 8.9 0.715 9.13 0.715 9.13 1.535 11.08 1.535 11.08 1.875 9.13 1.875 9.13 2.82 9.285 2.82 9.285 3.16 8.9 3.16  ;
        POLYGON 9.72 2.235 11.37 2.235 11.37 1.055 9.72 1.055 9.72 0.715 11.69 0.715 11.69 1.5 12.81 1.5 12.81 1.73 11.69 1.73 11.69 2.465 9.95 2.465 9.95 3.16 9.72 3.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyc_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlyc_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyc_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.36 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.93 1.2 3.405 1.2 3.405 1.6 0.93 1.6  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.4035 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.395 2.425 14.69 2.425 15.54 2.425 15.54 1.155 13.395 1.155 13.395 0.675 13.63 0.675 13.63 0.925 15.54 0.925 15.54 0.73 16.15 0.73 16.15 3.255 15.54 3.255 15.54 2.66 14.69 2.66 13.735 2.66 13.735 3.195 13.395 3.195  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.485 3.62 1.485 3.285 1.825 3.285 1.825 3.62 3.265 3.62 6.465 3.62 6.465 3.285 6.805 3.285 6.805 3.62 8.115 3.62 11.745 3.62 11.745 3.175 12.085 3.175 12.085 3.62 14.465 3.62 14.465 3.175 14.69 3.175 14.805 3.175 14.805 3.62 16.555 3.62 16.555 2.705 16.895 2.705 16.895 3.62 17.36 3.62 17.36 4.22 14.69 4.22 8.115 4.22 3.265 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.36 -0.3 17.36 0.3 16.99 0.3 16.99 0.695 16.76 0.695 16.76 0.3 14.75 0.3 14.75 0.695 14.52 0.695 14.52 0.3 12.155 0.3 12.155 0.695 11.925 0.695 11.925 0.3 7.005 0.3 7.005 0.635 6.665 0.635 6.665 0.3 1.925 0.3 1.925 0.635 1.585 0.635 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.065 3.265 2.065 3.265 2.405 0.585 2.405 0.585 3.105 0.245 3.105 0.245 0.67 0.585 0.67 0.585 0.9 0.475 0.9  ;
        POLYGON 3.72 0.77 4.105 0.77 4.105 1.465 5.8 1.465 5.8 1.805 3.95 1.805 3.95 3.16 3.72 3.16  ;
        POLYGON 4.385 2.875 6.03 2.875 6.03 1 4.485 1 4.485 0.77 6.26 0.77 6.26 1.52 8.115 1.52 8.115 1.75 6.26 1.75 6.26 3.105 4.385 3.105  ;
        POLYGON 8.9 0.715 9.13 0.715 9.13 1.535 11.08 1.535 11.08 1.875 9.13 1.875 9.13 2.82 9.285 2.82 9.285 3.16 8.9 3.16  ;
        POLYGON 9.72 2.235 11.37 2.235 11.37 1.055 9.72 1.055 9.72 0.715 11.69 0.715 11.69 1.53 14.69 1.53 14.69 1.76 11.69 1.76 11.69 2.465 9.95 2.465 9.95 3.16 9.72 3.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyc_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlyd_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyd_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.93 1.2 3.355 1.2 3.355 1.6 0.93 1.6  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.48 0.6 18.92 0.6 18.92 3.32 18.48 3.32  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.485 3.62 1.485 3.285 1.825 3.285 1.825 3.62 3.265 3.62 6.465 3.62 6.465 3.285 6.805 3.285 6.805 3.62 8.115 3.62 11.745 3.62 11.745 3.285 12.085 3.285 12.085 3.62 13.395 3.62 17.025 3.62 17.025 3.175 17.365 3.175 17.365 3.62 18.185 3.62 19.04 3.62 19.04 4.22 18.185 4.22 13.395 4.22 8.115 4.22 3.265 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 17.41 0.3 17.41 0.69 17.18 0.69 17.18 0.3 12.285 0.3 12.285 0.635 11.945 0.635 11.945 0.3 7.005 0.3 7.005 0.635 6.665 0.635 6.665 0.3 1.925 0.3 1.925 0.635 1.585 0.635 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.065 3.265 2.065 3.265 2.405 0.585 2.405 0.585 3.105 0.245 3.105 0.245 0.67 0.585 0.67 0.585 0.9 0.475 0.9  ;
        POLYGON 3.72 0.77 4.105 0.77 4.105 1.465 5.33 1.465 5.33 1.805 3.95 1.805 3.95 3.16 3.72 3.16  ;
        POLYGON 4.385 2.875 5.56 2.875 5.56 1 4.485 1 4.485 0.77 5.79 0.77 5.79 1.52 8.115 1.52 8.115 1.75 5.79 1.75 5.79 3.105 4.385 3.105  ;
        POLYGON 8.9 0.715 9.13 0.715 9.13 1.465 10.61 1.465 10.61 1.805 9.13 1.805 9.13 2.82 9.285 2.82 9.285 3.16 8.9 3.16  ;
        POLYGON 9.665 2.875 10.84 2.875 10.84 1 9.765 1 9.765 0.77 11.07 0.77 11.07 1.52 13.395 1.52 13.395 1.75 11.07 1.75 11.07 3.105 9.665 3.105  ;
        POLYGON 14.18 0.715 14.41 0.715 14.41 1.535 16.36 1.535 16.36 1.875 14.41 1.875 14.41 2.82 14.565 2.82 14.565 3.16 14.18 3.16  ;
        POLYGON 15 2.235 16.65 2.235 16.65 1 14.945 1 14.945 0.77 16.88 0.77 16.88 1.395 18.185 1.395 18.185 1.625 16.88 1.625 16.88 2.465 15.23 2.465 15.23 3.16 15 3.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyd_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlyd_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyd_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.16 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.93 1.2 3.395 1.2 3.395 1.6 0.93 1.6  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.48 0.675 18.95 0.675 18.95 3.38 18.48 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.485 3.62 1.485 3.285 1.825 3.285 1.825 3.62 3.265 3.62 6.465 3.62 6.465 3.285 6.805 3.285 6.805 3.62 8.115 3.62 11.745 3.62 11.745 3.285 12.085 3.285 12.085 3.62 13.395 3.62 17.46 3.62 17.46 2.53 17.69 2.53 17.69 3.62 18.185 3.62 19.5 3.62 19.5 2.53 19.73 2.53 19.73 3.62 20.16 3.62 20.16 4.22 18.185 4.22 13.395 4.22 8.115 4.22 3.265 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.16 -0.3 20.16 0.3 19.83 0.3 19.83 0.69 19.6 0.69 19.6 0.3 17.41 0.3 17.41 0.69 17.18 0.69 17.18 0.3 12.285 0.3 12.285 0.635 11.945 0.635 11.945 0.3 7.005 0.3 7.005 0.635 6.665 0.635 6.665 0.3 1.925 0.3 1.925 0.635 1.585 0.635 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.065 3.265 2.065 3.265 2.405 0.585 2.405 0.585 3.105 0.245 3.105 0.245 0.67 0.585 0.67 0.585 0.9 0.475 0.9  ;
        POLYGON 3.72 0.77 4.105 0.77 4.105 1.465 5.33 1.465 5.33 1.805 3.95 1.805 3.95 3.16 3.72 3.16  ;
        POLYGON 4.385 2.875 5.56 2.875 5.56 1 4.485 1 4.485 0.77 5.79 0.77 5.79 1.52 8.115 1.52 8.115 1.75 5.79 1.75 5.79 3.105 4.385 3.105  ;
        POLYGON 8.9 0.715 9.13 0.715 9.13 1.465 10.61 1.465 10.61 1.805 9.13 1.805 9.13 2.82 9.285 2.82 9.285 3.16 8.9 3.16  ;
        POLYGON 9.665 2.875 10.84 2.875 10.84 1 9.765 1 9.765 0.77 11.07 0.77 11.07 1.52 13.395 1.52 13.395 1.75 11.07 1.75 11.07 3.105 9.665 3.105  ;
        POLYGON 14.18 0.715 14.41 0.715 14.41 1.535 16.36 1.535 16.36 1.875 14.41 1.875 14.41 2.82 14.565 2.82 14.565 3.16 14.18 3.16  ;
        POLYGON 15 2.235 16.65 2.235 16.65 1 14.945 1 14.945 0.77 16.88 0.77 16.88 1.395 18.185 1.395 18.185 1.625 16.88 1.625 16.88 2.465 15.23 2.465 15.23 3.16 15 3.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyd_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__dlyd_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__dlyd_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.93 1.2 3.355 1.2 3.355 1.6 0.93 1.6  ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1216 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.48 2.165 20.065 2.165 20.72 2.165 20.72 1.15 18.425 1.15 18.425 0.73 18.765 0.73 18.765 0.92 20.72 0.92 20.72 0.675 21.19 0.675 21.19 3.38 20.72 3.38 20.72 2.395 20.065 2.395 18.71 2.395 18.71 3.38 18.48 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.485 3.62 1.485 3.285 1.825 3.285 1.825 3.62 3.265 3.62 6.465 3.62 6.465 3.285 6.805 3.285 6.805 3.62 8.115 3.62 11.745 3.62 11.745 3.285 12.085 3.285 12.085 3.62 13.395 3.62 17.46 3.62 17.46 2.53 17.69 2.53 17.69 3.62 19.525 3.62 19.525 2.625 19.865 2.625 19.865 3.62 20.065 3.62 21.74 3.62 21.74 2.53 21.97 2.53 21.97 3.62 22.4 3.62 22.4 4.22 20.065 4.22 13.395 4.22 8.115 4.22 3.265 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 22.07 0.3 22.07 0.69 21.84 0.69 21.84 0.3 19.83 0.3 19.83 0.69 19.6 0.69 19.6 0.3 17.41 0.3 17.41 0.69 17.18 0.69 17.18 0.3 12.285 0.3 12.285 0.635 11.945 0.635 11.945 0.3 7.005 0.3 7.005 0.635 6.665 0.635 6.665 0.3 1.925 0.3 1.925 0.635 1.585 0.635 1.585 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.475 2.065 3.265 2.065 3.265 2.405 0.585 2.405 0.585 3.105 0.245 3.105 0.245 0.67 0.585 0.67 0.585 0.9 0.475 0.9  ;
        POLYGON 3.72 0.77 4.105 0.77 4.105 1.465 5.33 1.465 5.33 1.805 3.95 1.805 3.95 3.16 3.72 3.16  ;
        POLYGON 4.385 2.875 5.56 2.875 5.56 1 4.485 1 4.485 0.77 5.79 0.77 5.79 1.52 8.115 1.52 8.115 1.75 5.79 1.75 5.79 3.105 4.385 3.105  ;
        POLYGON 8.9 0.715 9.13 0.715 9.13 1.465 10.61 1.465 10.61 1.805 9.13 1.805 9.13 2.82 9.285 2.82 9.285 3.16 8.9 3.16  ;
        POLYGON 9.665 2.875 10.84 2.875 10.84 1 9.765 1 9.765 0.77 11.07 0.77 11.07 1.52 13.395 1.52 13.395 1.75 11.07 1.75 11.07 3.105 9.665 3.105  ;
        POLYGON 14.18 0.715 14.41 0.715 14.41 1.535 16.36 1.535 16.36 1.875 14.41 1.875 14.41 2.82 14.565 2.82 14.565 3.16 14.18 3.16  ;
        POLYGON 15 2.235 16.65 2.235 16.65 1 14.945 1 14.945 0.77 16.88 0.77 16.88 1.59 20.065 1.59 20.065 1.82 16.88 1.82 16.88 2.465 15.23 2.465 15.23 3.16 15 3.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__dlyd_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__endcap
  CLASS ENDCAP PRE ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__endcap 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 1.12 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.37 3.62 0.37 1.92 0.71 1.92 0.71 3.62 1.12 3.62 1.12 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 1.12 -0.3 1.12 0.3 0.71 0.3 0.71 1.19 0.37 1.19 0.37 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__endcap

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fill_1
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 0.56 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.56 3.62 0.56 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 0.56 -0.3 0.56 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fill_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.96 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 8.96 3.62 8.96 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.96 -0.3 8.96 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_16

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fill_2
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 1.12 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.12 3.62 1.12 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 1.12 -0.3 1.12 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fill_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.92 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 17.92 3.62 17.92 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.92 -0.3 17.92 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_32

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fill_4
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 2.24 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.24 3.62 2.24 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 2.24 -0.3 2.24 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fill_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_64 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 35.84 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 35.84 3.62 35.84 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 35.84 -0.3 35.84 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_64

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fill_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fill_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 4.48 3.62 4.48 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__fill_8

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_16
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.96 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.765 3.62 1.765 2.49 1.995 2.49 1.995 3.62 4.005 3.62 4.005 2.49 4.235 2.49 4.235 3.62 6.245 3.62 6.245 2.49 6.475 2.49 6.475 3.62 8.485 3.62 8.485 2.49 8.715 2.49 8.715 3.62 8.96 3.62 8.96 4.22 8.715 4.22 6.475 4.22 4.235 4.22 1.995 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.96 -0.3 8.96 0.3 7.195 0.3 7.195 1.07 6.965 1.07 6.965 0.3 4.955 0.3 4.955 1.07 4.725 1.07 4.725 0.3 2.715 0.3 2.715 1.07 2.485 1.07 2.485 0.3 0.475 0.3 0.475 1.07 0.245 1.07 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.325 1.52 1.325 1.52 1.555 0.475 1.555 0.475 3.39 0.245 3.39  ;
        POLYGON 0.73 1.96 1.765 1.96 1.765 0.53 1.995 0.53 1.995 2.19 0.73 2.19  ;
        POLYGON 2.485 1.325 3.76 1.325 3.76 1.555 2.715 1.555 2.715 3.39 2.485 3.39  ;
        POLYGON 2.97 1.96 4.005 1.96 4.005 0.53 4.235 0.53 4.235 2.19 2.97 2.19  ;
        POLYGON 4.725 1.325 6 1.325 6 1.555 4.955 1.555 4.955 3.39 4.725 3.39  ;
        POLYGON 5.21 1.96 6.245 1.96 6.245 0.53 6.475 0.53 6.475 2.19 5.21 2.19  ;
        POLYGON 6.965 1.325 8.24 1.325 8.24 1.555 7.195 1.555 7.195 3.39 6.965 3.39  ;
        POLYGON 7.45 1.96 8.485 1.96 8.485 0.53 8.715 0.53 8.715 2.19 7.45 2.19  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_16

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_32
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_32 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.92 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.765 3.62 1.765 2.49 1.995 2.49 1.995 3.62 4.005 3.62 4.005 2.49 4.235 2.49 4.235 3.62 6.245 3.62 6.245 2.49 6.475 2.49 6.475 3.62 8.485 3.62 8.485 2.49 8.715 2.49 8.715 3.62 10.725 3.62 10.725 2.49 10.955 2.49 10.955 3.62 12.965 3.62 12.965 2.49 13.195 2.49 13.195 3.62 15.205 3.62 15.205 2.49 15.435 2.49 15.435 3.62 17.445 3.62 17.445 2.49 17.675 2.49 17.675 3.62 17.92 3.62 17.92 4.22 17.675 4.22 15.435 4.22 13.195 4.22 10.955 4.22 8.715 4.22 6.475 4.22 4.235 4.22 1.995 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.92 -0.3 17.92 0.3 16.155 0.3 16.155 1.045 15.925 1.045 15.925 0.3 13.915 0.3 13.915 1.045 13.685 1.045 13.685 0.3 11.675 0.3 11.675 1.045 11.445 1.045 11.445 0.3 9.435 0.3 9.435 1.045 9.205 1.045 9.205 0.3 7.195 0.3 7.195 1.045 6.965 1.045 6.965 0.3 4.955 0.3 4.955 1.045 4.725 1.045 4.725 0.3 2.715 0.3 2.715 1.045 2.485 1.045 2.485 0.3 0.475 0.3 0.475 1.045 0.245 1.045 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.325 1.52 1.325 1.52 1.555 0.475 1.555 0.475 3.39 0.245 3.39  ;
        POLYGON 0.73 1.96 1.765 1.96 1.765 0.53 1.995 0.53 1.995 2.19 0.73 2.19  ;
        POLYGON 2.485 1.325 3.76 1.325 3.76 1.555 2.715 1.555 2.715 3.39 2.485 3.39  ;
        POLYGON 2.97 1.96 4.005 1.96 4.005 0.53 4.235 0.53 4.235 2.19 2.97 2.19  ;
        POLYGON 4.725 1.325 6 1.325 6 1.555 4.955 1.555 4.955 3.39 4.725 3.39  ;
        POLYGON 5.21 1.96 6.245 1.96 6.245 0.53 6.475 0.53 6.475 2.19 5.21 2.19  ;
        POLYGON 6.965 1.325 8.24 1.325 8.24 1.555 7.195 1.555 7.195 3.39 6.965 3.39  ;
        POLYGON 7.45 1.96 8.485 1.96 8.485 0.53 8.715 0.53 8.715 2.19 7.45 2.19  ;
        POLYGON 9.205 1.325 10.48 1.325 10.48 1.555 9.435 1.555 9.435 3.39 9.205 3.39  ;
        POLYGON 9.69 1.96 10.725 1.96 10.725 0.53 10.955 0.53 10.955 2.19 9.69 2.19  ;
        POLYGON 11.445 1.325 12.72 1.325 12.72 1.555 11.675 1.555 11.675 3.39 11.445 3.39  ;
        POLYGON 11.93 1.96 12.965 1.96 12.965 0.53 13.195 0.53 13.195 2.19 11.93 2.19  ;
        POLYGON 13.685 1.325 14.96 1.325 14.96 1.555 13.915 1.555 13.915 3.39 13.685 3.39  ;
        POLYGON 14.17 1.96 15.205 1.96 15.205 0.53 15.435 0.53 15.435 2.19 14.17 2.19  ;
        POLYGON 15.925 1.325 17.2 1.325 17.2 1.555 16.155 1.555 16.155 3.39 15.925 3.39  ;
        POLYGON 16.41 1.96 17.445 1.96 17.445 0.53 17.675 0.53 17.675 2.19 16.41 2.19  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_32

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_4
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 2.24 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.765 3.62 1.765 2.49 1.995 2.49 1.995 3.62 2.24 3.62 2.24 4.22 1.995 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 2.24 -0.3 2.24 0.3 0.475 0.3 0.475 1.095 0.245 1.095 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.325 1.52 1.325 1.52 1.555 0.475 1.555 0.475 3.39 0.245 3.39  ;
        POLYGON 0.73 1.96 1.765 1.96 1.765 0.53 1.995 0.53 1.995 2.19 0.73 2.19  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_64
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_64 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 35.84 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.765 3.62 1.765 2.49 1.995 2.49 1.995 3.62 4.005 3.62 4.005 2.49 4.235 2.49 4.235 3.62 6.245 3.62 6.245 2.49 6.475 2.49 6.475 3.62 8.485 3.62 8.485 2.49 8.715 2.49 8.715 3.62 10.725 3.62 10.725 2.49 10.955 2.49 10.955 3.62 12.965 3.62 12.965 2.49 13.195 2.49 13.195 3.62 15.205 3.62 15.205 2.49 15.435 2.49 15.435 3.62 17.445 3.62 17.445 2.49 17.675 2.49 17.675 3.62 19.685 3.62 19.685 2.49 19.915 2.49 19.915 3.62 21.925 3.62 21.925 2.49 22.155 2.49 22.155 3.62 24.165 3.62 24.165 2.49 24.395 2.49 24.395 3.62 26.405 3.62 26.405 2.49 26.635 2.49 26.635 3.62 28.645 3.62 28.645 2.49 28.875 2.49 28.875 3.62 30.885 3.62 30.885 2.49 31.115 2.49 31.115 3.62 33.125 3.62 33.125 2.49 33.355 2.49 33.355 3.62 35.365 3.62 35.365 2.49 35.595 2.49 35.595 3.62 35.84 3.62 35.84 4.22 35.595 4.22 33.355 4.22 31.115 4.22 28.875 4.22 26.635 4.22 24.395 4.22 22.155 4.22 19.915 4.22 17.675 4.22 15.435 4.22 13.195 4.22 10.955 4.22 8.715 4.22 6.475 4.22 4.235 4.22 1.995 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 35.84 -0.3 35.84 0.3 34.075 0.3 34.075 1.055 33.845 1.055 33.845 0.3 31.835 0.3 31.835 1.055 31.605 1.055 31.605 0.3 29.595 0.3 29.595 1.055 29.365 1.055 29.365 0.3 27.355 0.3 27.355 1.055 27.125 1.055 27.125 0.3 25.115 0.3 25.115 1.055 24.885 1.055 24.885 0.3 22.875 0.3 22.875 1.055 22.645 1.055 22.645 0.3 20.635 0.3 20.635 1.055 20.405 1.055 20.405 0.3 18.395 0.3 18.395 1.055 18.165 1.055 18.165 0.3 16.155 0.3 16.155 1.055 15.925 1.055 15.925 0.3 13.915 0.3 13.915 1.055 13.685 1.055 13.685 0.3 11.675 0.3 11.675 1.055 11.445 1.055 11.445 0.3 9.435 0.3 9.435 1.055 9.205 1.055 9.205 0.3 7.195 0.3 7.195 1.055 6.965 1.055 6.965 0.3 4.955 0.3 4.955 1.055 4.725 1.055 4.725 0.3 2.715 0.3 2.715 1.055 2.485 1.055 2.485 0.3 0.475 0.3 0.475 1.055 0.245 1.055 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.325 1.52 1.325 1.52 1.555 0.475 1.555 0.475 3.39 0.245 3.39  ;
        POLYGON 0.73 1.96 1.765 1.96 1.765 0.53 1.995 0.53 1.995 2.19 0.73 2.19  ;
        POLYGON 2.485 1.325 3.76 1.325 3.76 1.555 2.715 1.555 2.715 3.39 2.485 3.39  ;
        POLYGON 2.97 1.96 4.005 1.96 4.005 0.53 4.235 0.53 4.235 2.19 2.97 2.19  ;
        POLYGON 4.725 1.325 6 1.325 6 1.555 4.955 1.555 4.955 3.39 4.725 3.39  ;
        POLYGON 5.21 1.96 6.245 1.96 6.245 0.53 6.475 0.53 6.475 2.19 5.21 2.19  ;
        POLYGON 6.965 1.325 8.24 1.325 8.24 1.555 7.195 1.555 7.195 3.39 6.965 3.39  ;
        POLYGON 7.45 1.96 8.485 1.96 8.485 0.53 8.715 0.53 8.715 2.19 7.45 2.19  ;
        POLYGON 9.205 1.325 10.48 1.325 10.48 1.555 9.435 1.555 9.435 3.39 9.205 3.39  ;
        POLYGON 9.69 1.96 10.725 1.96 10.725 0.53 10.955 0.53 10.955 2.19 9.69 2.19  ;
        POLYGON 11.445 1.325 12.72 1.325 12.72 1.555 11.675 1.555 11.675 3.39 11.445 3.39  ;
        POLYGON 11.93 1.96 12.965 1.96 12.965 0.53 13.195 0.53 13.195 2.19 11.93 2.19  ;
        POLYGON 13.685 1.325 14.96 1.325 14.96 1.555 13.915 1.555 13.915 3.39 13.685 3.39  ;
        POLYGON 14.17 1.96 15.205 1.96 15.205 0.53 15.435 0.53 15.435 2.19 14.17 2.19  ;
        POLYGON 15.925 1.325 17.2 1.325 17.2 1.555 16.155 1.555 16.155 3.39 15.925 3.39  ;
        POLYGON 16.41 1.96 17.445 1.96 17.445 0.53 17.675 0.53 17.675 2.19 16.41 2.19  ;
        POLYGON 18.165 1.325 19.44 1.325 19.44 1.555 18.395 1.555 18.395 3.39 18.165 3.39  ;
        POLYGON 18.65 1.96 19.685 1.96 19.685 0.53 19.915 0.53 19.915 2.19 18.65 2.19  ;
        POLYGON 20.405 1.325 21.68 1.325 21.68 1.555 20.635 1.555 20.635 3.39 20.405 3.39  ;
        POLYGON 20.89 1.96 21.925 1.96 21.925 0.53 22.155 0.53 22.155 2.19 20.89 2.19  ;
        POLYGON 22.645 1.325 23.92 1.325 23.92 1.555 22.875 1.555 22.875 3.39 22.645 3.39  ;
        POLYGON 23.13 1.96 24.165 1.96 24.165 0.53 24.395 0.53 24.395 2.19 23.13 2.19  ;
        POLYGON 24.885 1.325 26.16 1.325 26.16 1.555 25.115 1.555 25.115 3.39 24.885 3.39  ;
        POLYGON 25.37 1.96 26.405 1.96 26.405 0.53 26.635 0.53 26.635 2.19 25.37 2.19  ;
        POLYGON 27.125 1.325 28.4 1.325 28.4 1.555 27.355 1.555 27.355 3.39 27.125 3.39  ;
        POLYGON 27.61 1.96 28.645 1.96 28.645 0.53 28.875 0.53 28.875 2.19 27.61 2.19  ;
        POLYGON 29.365 1.325 30.64 1.325 30.64 1.555 29.595 1.555 29.595 3.39 29.365 3.39  ;
        POLYGON 29.85 1.96 30.885 1.96 30.885 0.53 31.115 0.53 31.115 2.19 29.85 2.19  ;
        POLYGON 31.605 1.325 32.88 1.325 32.88 1.555 31.835 1.555 31.835 3.39 31.605 3.39  ;
        POLYGON 32.09 1.96 33.125 1.96 33.125 0.53 33.355 0.53 33.355 2.19 32.09 2.19  ;
        POLYGON 33.845 1.325 35.12 1.325 35.12 1.555 34.075 1.555 34.075 3.39 33.845 3.39  ;
        POLYGON 34.33 1.96 35.365 1.96 35.365 0.53 35.595 0.53 35.595 2.19 34.33 2.19  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_64

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__fillcap_8
  CLASS core SPACER ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__fillcap_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.765 3.62 1.765 2.49 1.995 2.49 1.995 3.62 4.005 3.62 4.005 2.49 4.235 2.49 4.235 3.62 4.48 3.62 4.48 4.22 4.235 4.22 1.995 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 2.715 0.3 2.715 1.085 2.485 1.085 2.485 0.3 0.475 0.3 0.475 1.085 0.245 1.085 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 1.325 1.52 1.325 1.52 1.555 0.475 1.555 0.475 3.39 0.245 3.39  ;
        POLYGON 0.73 1.96 1.765 1.96 1.765 0.53 1.995 0.53 1.995 2.19 0.73 2.19  ;
        POLYGON 2.485 1.325 3.76 1.325 3.76 1.555 2.715 1.555 2.715 3.39 2.485 3.39  ;
        POLYGON 2.97 1.96 4.005 1.96 4.005 0.53 4.235 0.53 4.235 2.19 2.97 2.19  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__fillcap_8

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__filltie
  CLASS core WELLTAP ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__filltie 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 1.12 BY 3.92 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.39 3.62 0.39 1.93 0.73 1.93 0.73 3.62 1.12 3.62 1.12 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 1.12 -0.3 1.12 0.3 0.73 0.3 0.73 1.185 0.39 1.185 0.39 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__filltie

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__hold
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__hold 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.04 BY 3.92 ;
  PIN Z
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.4512 ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.245 0.565 0.475 0.565 0.475 1.155 3.95 1.155 3.95 1.56 0.575 1.56 0.575 2.895 0.245 2.895  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 3.225 3.62 3.225 2.535 3.455 2.535 3.455 3.62 4.575 3.62 5.04 3.62 5.04 4.22 4.575 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.04 -0.3 5.04 0.3 3.455 0.3 3.455 0.925 3.225 0.925 3.225 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.45 1.885 4.345 1.885 4.345 0.575 4.575 0.575 4.575 3.18 4.245 3.18 4.245 2.185 2.45 2.185  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__hold

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__icgtn_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtn_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.36 BY 3.92 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.394 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.81 1.21 13.865 1.21 13.865 1.45 14.255 1.45 14.255 2.195 14.025 2.195 14.025 1.68 13.57 1.68 13.57 1.59 11.81 1.59  ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.845 1.77 2.73 1.77 2.73 3.37 2.32 3.37 2.32 2.15 1.845 2.15  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.27 1.77 1.57 1.77 1.57 2.15 0.27 2.15  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8118 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.3 0.63 17.035 0.63 17.035 3.27 16.3 3.27  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.48 0.575 2.48 0.575 3.62 2.77 3.62 6.3 3.62 6.3 2.79 6.53 2.79 6.53 3.62 8.79 3.62 9.11 3.62 9.11 2.47 9.34 2.47 9.34 3.62 9.91 3.62 12.8 3.62 12.8 2.46 13.03 2.46 13.03 3.62 13.63 3.62 15.345 3.62 15.345 2.425 15.685 2.425 15.685 3.62 16.07 3.62 17.36 3.62 17.36 4.22 16.07 4.22 13.63 4.22 9.91 4.22 8.79 4.22 2.77 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.36 -0.3 17.36 0.3 15.91 0.3 15.91 1.095 15.68 1.095 15.68 0.3 15.245 0.3 15.245 0.76 14.905 0.76 14.905 0.3 13.005 0.3 13.005 0.76 12.665 0.76 12.665 0.3 9.445 0.3 9.445 1.075 9.105 1.075 9.105 0.3 6.405 0.3 6.405 1.075 6.065 1.075 6.065 0.3 1.65 0.3 1.65 1.06 1.31 1.06 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.845 0.53 0.845 0.53 1.29 1.885 1.29 1.885 0.845 2.77 0.845 2.77 1.075 2.115 1.075 2.115 1.52 0.19 1.52  ;
        POLYGON 3.46 1.42 3.69 1.42 3.69 1.87 7.32 1.87 7.32 0.78 7.55 0.78 7.55 2.9 7.32 2.9 7.32 2.1 3.46 2.1  ;
        POLYGON 3.23 2.33 7.04 2.33 7.04 3.16 8.56 3.16 8.56 1.82 8.79 1.82 8.79 3.39 6.81 3.39 6.81 2.56 4.04 2.56 4.04 3.125 3.81 3.125 3.81 2.56 3 2.56 3 0.845 3.89 0.845 3.89 1.075 3.23 1.075  ;
        POLYGON 8.04 0.78 8.27 0.78 8.27 1.34 9.91 1.34 9.91 1.575 8.27 1.575 8.27 2.9 8.04 2.9  ;
        POLYGON 11.09 2.26 12.01 2.26 12.01 2.93 11.78 2.93 11.78 2.495 10.86 2.495 10.86 0.53 11.975 0.53 11.975 0.76 11.09 0.76  ;
        POLYGON 10.18 0.78 10.51 0.78 10.51 3.16 12.34 3.16 12.34 1.91 13.63 1.91 13.63 2.14 12.57 2.14 12.57 3.39 10.18 3.39  ;
        POLYGON 13.785 0.53 14.57 0.53 14.57 0.99 14.79 0.99 14.79 1.79 16.07 1.79 16.07 2.13 14.79 2.13 14.79 3.18 14.56 3.18 14.56 1.22 14.34 1.22 14.34 0.76 13.785 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtn_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__icgtn_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtn_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 18.48 BY 3.92 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.725 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.81 1.21 14.215 1.21 14.215 2.25 13.985 2.25 13.985 1.59 11.81 1.59  ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.865 1.77 2.75 1.77 2.75 3.37 2.34 3.37 2.34 2.15 1.865 2.15  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.29 1.77 1.59 1.77 1.59 2.15 0.29 2.15  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.962 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.455 2.37 17.19 2.37 17.45 2.37 17.45 1.415 16.75 1.415 16.75 0.6 17.22 0.6 17.22 1.145 17.83 1.145 17.83 2.71 17.19 2.71 16.795 2.71 16.795 3.305 16.455 3.305  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.48 0.575 2.48 0.575 3.62 2.77 3.62 6.3 3.62 6.3 2.79 6.53 2.79 6.53 3.62 8.79 3.62 9.11 3.62 9.11 2.47 9.34 2.47 9.34 3.62 9.91 3.62 12.8 3.62 12.8 2.695 13.03 2.695 13.03 3.62 13.63 3.62 15.49 3.62 15.49 2.61 15.72 2.61 15.72 3.62 17.19 3.62 17.53 3.62 17.53 3.02 17.76 3.02 17.76 3.62 18.48 3.62 18.48 4.22 17.19 4.22 13.63 4.22 9.91 4.22 8.79 4.22 2.77 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 18.48 -0.3 18.48 0.3 18.15 0.3 18.15 0.915 17.92 0.915 17.92 0.3 15.91 0.3 15.91 1.09 15.68 1.09 15.68 0.3 15.245 0.3 15.245 0.76 14.905 0.76 14.905 0.3 13.005 0.3 13.005 0.76 12.665 0.76 12.665 0.3 9.445 0.3 9.445 1.075 9.105 1.075 9.105 0.3 6.405 0.3 6.405 1.075 6.065 1.075 6.065 0.3 1.65 0.3 1.65 1.06 1.31 1.06 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.845 0.53 0.845 0.53 1.29 1.885 1.29 1.885 0.845 2.77 0.845 2.77 1.075 2.115 1.075 2.115 1.52 0.19 1.52  ;
        POLYGON 3.46 1.42 3.69 1.42 3.69 1.87 7.32 1.87 7.32 0.78 7.55 0.78 7.55 2.9 7.32 2.9 7.32 2.1 3.46 2.1  ;
        POLYGON 3.23 2.33 7.04 2.33 7.04 3.16 8.56 3.16 8.56 1.82 8.79 1.82 8.79 3.39 6.81 3.39 6.81 2.56 4.04 2.56 4.04 3.265 3.81 3.265 3.81 2.56 3 2.56 3 0.845 3.89 0.845 3.89 1.075 3.23 1.075  ;
        POLYGON 8.04 0.78 8.27 0.78 8.27 1.34 9.91 1.34 9.91 1.575 8.27 1.575 8.27 2.9 8.04 2.9  ;
        POLYGON 11.09 2.26 12.01 2.26 12.01 2.93 11.78 2.93 11.78 2.495 10.86 2.495 10.86 0.53 11.885 0.53 11.885 0.76 11.09 0.76  ;
        POLYGON 10.18 0.78 10.51 0.78 10.51 3.16 12.34 3.16 12.34 1.91 13.63 1.91 13.63 2.14 12.57 2.14 12.57 3.39 10.18 3.39  ;
        POLYGON 13.785 0.53 14.675 0.53 14.675 0.99 14.79 0.99 14.79 1.79 17.19 1.79 17.19 2.14 14.79 2.14 14.79 3.18 14.56 3.18 14.56 2.13 14.445 2.13 14.445 0.76 13.785 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtn_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__icgtn_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtn_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.72 BY 3.92 ;
  PIN CLKN
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.725 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.81 1.21 13.865 1.21 13.865 1.45 14.255 1.45 14.255 2.195 14.025 2.195 14.025 1.68 13.57 1.68 13.57 1.59 11.81 1.59  ;
    END
  END CLKN
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.865 1.8 2.75 1.8 2.75 3.37 2.34 3.37 2.34 2.12 1.865 2.12  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.29 1.8 1.59 1.8 1.59 2.12 0.29 2.12  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.924 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.51 2.37 19.28 2.37 19.69 2.37 19.69 1.535 16.75 1.535 16.75 0.6 17.22 0.6 17.22 1.265 19.04 1.265 19.04 0.6 19.47 0.6 19.47 1.265 20.07 1.265 20.07 2.71 19.28 2.71 18.78 2.71 18.78 3.18 18.55 3.18 18.55 2.71 16.74 2.71 16.74 3.18 16.51 3.18  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.48 0.575 2.48 0.575 3.62 2.77 3.62 6.3 3.62 6.3 2.79 6.53 2.79 6.53 3.62 8.79 3.62 9.11 3.62 9.11 2.47 9.34 2.47 9.34 3.62 9.91 3.62 12.8 3.62 12.8 2.645 13.03 2.645 13.03 3.62 13.63 3.62 15.49 3.62 15.49 2.645 15.72 2.645 15.72 3.62 17.53 3.62 17.53 3.02 17.76 3.02 17.76 3.62 19.28 3.62 19.57 3.62 19.57 3.02 19.8 3.02 19.8 3.62 20.72 3.62 20.72 4.22 19.28 4.22 13.63 4.22 9.91 4.22 8.79 4.22 2.77 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.72 -0.3 20.72 0.3 20.39 0.3 20.39 0.975 20.16 0.975 20.16 0.3 18.15 0.3 18.15 0.975 17.92 0.975 17.92 0.3 15.91 0.3 15.91 1.09 15.68 1.09 15.68 0.3 15.245 0.3 15.245 0.76 14.905 0.76 14.905 0.3 13.005 0.3 13.005 0.76 12.665 0.76 12.665 0.3 9.445 0.3 9.445 1.075 9.105 1.075 9.105 0.3 6.405 0.3 6.405 1.075 6.065 1.075 6.065 0.3 1.65 0.3 1.65 1.06 1.31 1.06 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.845 0.53 0.845 0.53 1.305 1.885 1.305 1.885 0.845 2.77 0.845 2.77 1.075 2.115 1.075 2.115 1.54 0.19 1.54  ;
        POLYGON 3.46 1.42 3.69 1.42 3.69 1.87 7.32 1.87 7.32 0.78 7.55 0.78 7.55 2.9 7.32 2.9 7.32 2.1 3.46 2.1  ;
        POLYGON 3.23 2.33 7.04 2.33 7.04 3.16 8.56 3.16 8.56 1.82 8.79 1.82 8.79 3.39 6.81 3.39 6.81 2.56 4.04 2.56 4.04 3.265 3.81 3.265 3.81 2.56 3 2.56 3 0.845 3.89 0.845 3.89 1.075 3.23 1.075  ;
        POLYGON 8.04 0.78 8.27 0.78 8.27 1.34 9.91 1.34 9.91 1.575 8.27 1.575 8.27 2.9 8.04 2.9  ;
        POLYGON 11.09 2.26 12.01 2.26 12.01 2.93 11.78 2.93 11.78 2.495 10.86 2.495 10.86 0.53 11.975 0.53 11.975 0.76 11.09 0.76  ;
        POLYGON 10.18 0.78 10.51 0.78 10.51 3.16 12.34 3.16 12.34 1.91 13.63 1.91 13.63 2.14 12.57 2.14 12.57 3.39 10.18 3.39  ;
        POLYGON 13.785 0.53 14.57 0.53 14.57 0.99 14.79 0.99 14.79 1.79 19.28 1.79 19.28 2.14 14.79 2.14 14.79 3.18 14.56 3.18 14.56 1.22 14.34 1.22 14.34 0.76 13.785 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtn_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__icgtp_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtp_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.68 BY 3.92 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.388 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.215 1.535 10.785 1.535 10.785 1.21 11.235 1.21 12.755 1.21 12.755 1.59 11.235 1.59 11.065 1.59 11.065 1.765 10.215 1.765  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.865 1.77 2.75 1.77 2.75 3.37 2.34 3.37 2.34 2.15 1.865 2.15  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.29 1.77 1.59 1.77 1.59 2.15 0.29 2.15  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.814 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.16 2.33 14.55 2.33 14.78 2.33 14.78 1.12 14.7 1.12 14.7 0.56 15.23 0.56 15.23 3.27 14.55 3.27 14.16 3.27  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.48 0.575 2.48 0.575 3.62 2.77 3.62 6.245 3.62 6.245 2.845 6.585 2.845 6.585 3.62 9.69 3.62 9.69 2.92 9.92 2.92 9.92 3.62 11.635 3.62 11.635 2.46 11.865 2.46 11.865 3.62 13.7 3.62 13.7 2.9 13.93 2.9 13.93 3.62 14.55 3.62 15.68 3.62 15.68 4.22 14.55 4.22 2.77 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 15.68 -0.3 15.68 0.3 13.93 0.3 13.93 0.805 13.7 0.805 13.7 0.3 10.05 0.3 10.05 0.845 9.82 0.845 9.82 0.3 6.405 0.3 6.405 1.075 6.065 1.075 6.065 0.3 1.65 0.3 1.65 0.995 1.31 0.995 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.765 0.53 0.765 0.53 1.225 1.885 1.225 1.885 0.765 2.77 0.765 2.77 0.995 2.115 0.995 2.115 1.46 0.19 1.46  ;
        POLYGON 3.46 1.445 3.69 1.445 3.69 1.87 4.935 1.87 4.935 2.1 3.46 2.1  ;
        POLYGON 3.23 2.33 5.205 2.33 5.205 1.34 7.08 1.34 7.08 1.575 5.435 1.575 5.435 2.56 4.04 2.56 4.04 3.125 3.81 3.125 3.81 2.56 3 2.56 3 0.765 3.89 0.765 3.89 0.995 3.23 0.995  ;
        POLYGON 7.915 0.53 9.075 0.53 9.075 0.76 8.275 0.76 8.275 1.805 8.93 1.805 8.93 2.85 8.645 2.85 8.645 2.035 7.915 2.035  ;
        POLYGON 9.245 1.075 10.28 1.075 10.28 0.53 11.235 0.53 11.235 0.76 10.51 0.76 10.51 1.305 9.485 1.305 9.485 1.995 10.945 1.995 10.945 2.85 10.715 2.85 10.715 2.225 9.245 2.225  ;
        POLYGON 5.685 1.805 7.32 1.805 7.32 0.78 7.55 0.78 7.55 3.16 9.165 3.16 9.165 2.455 10.43 2.455 10.43 3.16 11.175 3.16 11.175 1.995 12.01 1.995 12.01 1.965 13.415 1.965 13.415 2.21 12.265 2.21 12.265 2.225 11.405 2.225 11.405 3.39 10.2 3.39 10.2 2.69 9.395 2.69 9.395 3.39 7.32 3.39 7.32 2.035 5.685 2.035  ;
        POLYGON 12.68 2.44 13.645 2.44 13.645 1.535 13.01 1.535 13.01 0.76 11.595 0.76 11.595 0.53 13.24 0.53 13.24 1.265 13.875 1.265 13.875 1.685 14.55 1.685 14.55 2.025 13.875 2.025 13.875 2.67 12.91 2.67 12.91 3.25 12.68 3.25  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtp_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__icgtp_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtp_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 16.8 BY 3.92 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.679 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.11 1.535 10.74 1.535 10.74 1.21 11.235 1.21 12.755 1.21 12.755 1.59 11.235 1.59 10.97 1.59 10.97 1.765 10.11 1.765  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.865 1.8 2.75 1.8 2.75 3.37 2.34 3.37 2.34 2.12 1.865 2.12  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.29 1.8 1.59 1.8 1.59 2.12 0.29 2.12  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.118 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.66 2.4 14.97 2.4 15.22 2.4 15.22 1.08 14.555 1.08 14.555 0.6 15.58 0.6 15.58 2.74 15.02 2.74 15.02 3.38 14.97 3.38 14.66 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.29 3.62 0.29 2.535 0.63 2.535 0.63 3.62 2.77 3.62 6.28 3.62 6.28 2.505 6.51 2.505 6.51 3.62 9.69 3.62 9.69 2.92 9.92 2.92 9.92 3.62 11.635 3.62 11.635 2.57 11.865 2.57 11.865 3.62 13.645 3.62 13.645 2.815 13.985 2.815 13.985 3.62 14.97 3.62 15.87 3.62 15.87 2.53 16.1 2.53 16.1 3.62 16.8 3.62 16.8 4.22 14.97 4.22 2.77 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 16.8 -0.3 16.8 0.3 16.235 0.3 16.235 0.75 15.885 0.75 15.885 0.3 13.93 0.3 13.93 0.845 13.7 0.845 13.7 0.3 10.05 0.3 10.05 0.845 9.82 0.845 9.82 0.3 6.405 0.3 6.405 1.075 6.065 1.075 6.065 0.3 1.65 0.3 1.65 0.995 1.31 0.995 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.765 0.53 0.765 0.53 1.225 1.885 1.225 1.885 0.765 2.77 0.765 2.77 0.995 2.115 0.995 2.115 1.46 0.19 1.46  ;
        POLYGON 3.46 1.445 3.69 1.445 3.69 1.87 4.935 1.87 4.935 2.1 3.46 2.1  ;
        POLYGON 3.23 2.33 5.205 2.33 5.205 1.34 7.08 1.34 7.08 1.575 5.435 1.575 5.435 2.56 4.04 2.56 4.04 3.265 3.81 3.265 3.81 2.56 3 2.56 3 0.765 3.89 0.765 3.89 0.995 3.23 0.995  ;
        POLYGON 7.915 0.53 9.075 0.53 9.075 0.76 8.275 0.76 8.275 1.805 8.93 1.805 8.93 2.85 8.645 2.85 8.645 2.035 7.915 2.035  ;
        POLYGON 9.175 1.075 10.28 1.075 10.28 0.53 11.235 0.53 11.235 0.76 10.51 0.76 10.51 1.305 9.415 1.305 9.415 1.995 10.945 1.995 10.945 2.85 10.715 2.85 10.715 2.225 9.175 2.225  ;
        POLYGON 5.685 1.805 7.32 1.805 7.32 0.78 7.55 0.78 7.55 3.16 9.165 3.16 9.165 2.455 10.43 2.455 10.43 3.16 11.175 3.16 11.175 1.895 13.415 1.895 13.415 2.125 11.405 2.125 11.405 3.39 10.2 3.39 10.2 2.69 9.395 2.69 9.395 3.39 7.32 3.39 7.32 2.035 5.685 2.035  ;
        POLYGON 12.68 2.355 13.645 2.355 13.645 1.535 13.01 1.535 13.01 0.76 11.595 0.76 11.595 0.53 13.24 0.53 13.24 1.265 13.875 1.265 13.875 1.595 14.97 1.595 14.97 1.825 13.875 1.825 13.875 2.585 12.91 2.585 12.91 3.38 12.68 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtp_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__icgtp_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__icgtp_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.685 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.105 1.535 10.785 1.535 10.785 1.21 11.235 1.21 12.755 1.21 12.755 1.59 11.235 1.59 11.065 1.59 11.065 1.765 10.105 1.765  ;
    END
  END CLK
  PIN E
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.865 1.77 2.71 1.77 2.71 3.27 2.33 3.27 2.33 2.15 1.865 2.15  ;
    END
  END E
  PIN TE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.6995 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.29 1.77 1.59 1.77 1.59 2.15 0.29 2.15  ;
    END
  END TE
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.924 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.7 2.33 17.57 2.33 18.01 2.33 18.01 1.535 14.82 1.535 14.82 0.705 15.05 0.705 15.05 1.265 17.06 1.265 17.06 0.705 17.29 0.705 17.29 1.265 18.39 1.265 18.39 2.71 17.57 2.71 16.99 2.71 16.99 3.195 16.76 3.195 16.76 2.71 14.975 2.71 14.975 3.195 14.7 3.195  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.48 0.575 2.48 0.575 3.62 2.77 3.62 6.28 3.62 6.28 2.605 6.51 2.605 6.51 3.62 9.69 3.62 9.69 2.92 9.92 2.92 9.92 3.62 11.635 3.62 11.635 2.76 11.865 2.76 11.865 3.62 13.7 3.62 13.7 3.04 13.93 3.04 13.93 3.62 15.74 3.62 15.74 3.04 15.97 3.04 15.97 3.62 17.57 3.62 17.78 3.62 17.78 3.045 18.01 3.045 18.01 3.62 19.04 3.62 19.04 4.22 17.57 4.22 2.77 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 18.41 0.3 18.41 0.805 18.18 0.805 18.18 0.3 16.17 0.3 16.17 0.805 15.94 0.805 15.94 0.3 13.93 0.3 13.93 0.805 13.7 0.805 13.7 0.3 10.05 0.3 10.05 0.845 9.82 0.845 9.82 0.3 6.405 0.3 6.405 1.075 6.065 1.075 6.065 0.3 1.65 0.3 1.65 0.995 1.31 0.995 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.765 0.53 0.765 0.53 1.225 1.885 1.225 1.885 0.765 2.77 0.765 2.77 0.995 2.115 0.995 2.115 1.46 0.19 1.46  ;
        POLYGON 3.46 1.445 3.69 1.445 3.69 1.87 4.935 1.87 4.935 2.1 3.46 2.1  ;
        POLYGON 3.23 2.33 5.205 2.33 5.205 1.34 7.08 1.34 7.08 1.575 5.435 1.575 5.435 2.56 4.04 2.56 4.04 3.125 3.81 3.125 3.81 2.56 3 2.56 3 0.765 3.89 0.765 3.89 0.995 3.23 0.995  ;
        POLYGON 7.915 0.53 9.075 0.53 9.075 0.76 8.275 0.76 8.275 1.805 8.93 1.805 8.93 2.85 8.645 2.85 8.645 2.035 7.915 2.035  ;
        POLYGON 9.175 1.075 10.28 1.075 10.28 0.53 11.235 0.53 11.235 0.76 10.51 0.76 10.51 1.305 9.415 1.305 9.415 1.995 10.945 1.995 10.945 2.85 10.715 2.85 10.715 2.225 9.175 2.225  ;
        POLYGON 5.685 1.805 7.32 1.805 7.32 0.78 7.55 0.78 7.55 3.16 9.165 3.16 9.165 2.455 10.43 2.455 10.43 3.16 11.175 3.16 11.175 1.995 13.075 1.995 13.075 1.965 13.415 1.965 13.415 2.225 11.405 2.225 11.405 3.39 10.2 3.39 10.2 2.69 9.395 2.69 9.395 3.39 7.32 3.39 7.32 2.035 5.685 2.035  ;
        POLYGON 12.68 2.455 13.7 2.455 13.7 1.535 13.105 1.535 13.105 0.76 11.595 0.76 11.595 0.53 13.335 0.53 13.335 1.265 13.93 1.265 13.93 1.825 17.57 1.825 17.57 2.095 13.93 2.095 13.93 2.685 12.91 2.685 12.91 3.265 12.68 3.265  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__icgtp_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 2.24 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 1.2 1.035 1.2 1.035 2.2 0.71 2.2  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 0.53 1.595 0.53 1.595 3.39 1.265 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.575 2.53 0.575 3.62 2.24 3.62 2.24 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 2.24 -0.3 2.24 0.3 0.475 0.3 0.475 1.16 0.245 1.16 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 13.224 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.64 1.765 6.155 1.765 6.155 2.15 0.64 2.15  ;
        POLYGON 7.8 1.765 13.31 1.765 13.31 2.15 7.8 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 7.0968 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.52 6.55 2.52 6.55 1.45 1.365 1.45 1.365 0.675 1.595 0.675 1.595 1.01 3.605 1.01 3.605 0.675 3.835 0.675 3.835 1.01 5.845 1.01 5.845 0.675 6.075 0.675 6.075 1.01 8.085 1.01 8.085 0.675 8.315 0.675 8.315 1.01 10.325 1.01 10.325 0.675 10.555 0.675 10.555 1.01 12.565 1.01 12.565 0.675 12.795 0.675 12.795 1.45 7.45 1.45 7.45 2.535 12.695 2.535 12.695 3.39 12.465 3.39 12.465 2.96 10.455 2.96 10.455 3.39 10.225 3.39 10.225 2.96 8.215 2.96 8.215 3.39 7.985 3.39 7.985 2.96 5.975 2.96 5.975 3.39 5.745 3.39 5.745 2.96 3.735 2.96 3.735 3.39 3.505 3.39 3.505 2.96 1.595 2.96 1.595 3.39 1.365 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.68 0.475 2.68 0.475 3.62 2.385 3.62 2.385 3.21 2.615 3.21 2.615 3.62 4.625 3.62 4.625 3.21 4.855 3.21 4.855 3.62 6.865 3.62 6.865 3.21 7.095 3.21 7.095 3.62 9.105 3.62 9.105 3.21 9.335 3.21 9.335 3.62 11.345 3.62 11.345 3.21 11.575 3.21 11.575 3.62 13.585 3.62 13.585 2.68 13.815 2.68 13.815 3.62 14.56 3.62 14.56 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 13.915 0.3 13.915 1.015 13.685 1.015 13.685 0.3 11.675 0.3 11.675 0.69 11.445 0.69 11.445 0.3 9.435 0.3 9.435 0.69 9.205 0.69 9.205 0.3 7.195 0.3 7.195 0.69 6.965 0.69 6.965 0.3 4.955 0.3 4.955 0.69 4.725 0.69 4.725 0.3 2.715 0.3 2.715 0.69 2.485 0.69 2.485 0.3 0.475 0.3 0.475 1.015 0.245 1.015 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_12

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 17.632 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.765 8.51 1.765 8.51 2.19 0.62 2.19  ;
        POLYGON 10.015 1.765 17.92 1.765 17.92 2.19 10.015 2.19  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.4624 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.42 8.79 2.42 8.79 1.445 1.365 1.445 1.365 0.675 1.625 0.675 1.625 0.865 3.605 0.865 3.605 0.675 3.835 0.675 3.835 0.865 5.845 0.865 5.845 0.675 6.075 0.675 6.075 0.865 8.085 0.865 8.085 0.675 8.315 0.675 8.315 0.865 10.325 0.865 10.325 0.675 10.555 0.675 10.555 0.865 12.565 0.865 12.565 0.675 12.795 0.675 12.795 0.865 14.805 0.865 14.805 0.675 15.035 0.675 15.035 0.865 17.045 0.865 17.045 0.675 17.275 0.675 17.275 1.445 9.69 1.445 9.69 2.42 17.175 2.42 17.175 3.39 16.945 3.39 16.945 3 14.935 3 14.935 3.39 14.705 3.39 14.705 3 12.695 3 12.695 3.39 12.465 3.39 12.465 3 10.455 3 10.455 3.39 10.225 3.39 10.225 3 8.31 3 8.31 3.39 8.08 3.39 8.08 3 5.975 3 5.975 3.39 5.745 3.39 5.745 3 3.735 3 3.735 3.39 3.505 3.39 3.505 3 1.595 3 1.595 3.39 1.365 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.68 0.475 2.68 0.475 3.62 2.385 3.62 2.385 3.23 2.615 3.23 2.615 3.62 4.625 3.62 4.625 3.23 4.855 3.23 4.855 3.62 6.865 3.62 6.865 3.23 7.095 3.23 7.095 3.62 9.105 3.62 9.105 3.23 9.335 3.23 9.335 3.62 11.345 3.62 11.345 3.23 11.575 3.23 11.575 3.62 13.585 3.62 13.585 3.23 13.815 3.23 13.815 3.62 15.825 3.62 15.825 3.23 16.055 3.23 16.055 3.62 18.065 3.62 18.065 2.68 18.295 2.68 18.295 3.62 19.04 3.62 19.04 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 18.395 0.3 18.395 1.015 18.165 1.015 18.165 0.3 16.21 0.3 16.21 0.635 15.87 0.635 15.87 0.3 13.97 0.3 13.97 0.635 13.63 0.635 13.63 0.3 11.73 0.3 11.73 0.635 11.39 0.635 11.39 0.3 9.49 0.3 9.49 0.635 9.15 0.635 9.15 0.3 7.25 0.3 7.25 0.635 6.91 0.635 6.91 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.475 0.3 0.475 1.015 0.245 1.015 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_16

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 3.36 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.705 2.15 1.705 2.15 2.12 0.63 2.12  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.366 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.22 2.36 2.38 2.36 2.38 1.475 1.395 1.475 1.395 0.53 1.625 0.53 1.625 1.22 2.68 1.22 2.68 2.68 1.67 2.68 1.67 3.39 1.22 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.64 0.475 2.64 0.475 3.62 2.515 3.62 2.515 2.93 2.745 2.93 2.745 3.62 3.36 3.62 3.36 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 3.36 -0.3 3.36 0.3 2.745 0.3 2.745 0.95 2.515 0.95 2.515 0.3 0.475 0.3 0.475 0.95 0.245 0.95 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_20
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_20 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 23.52 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 22.04 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.61 1.765 8.02 1.765 8.02 2.15 0.61 2.15  ;
        POLYGON 14.985 1.765 22.375 1.765 22.375 2.15 14.985 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 11.828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.38 8.395 2.38 8.395 2.315 11.03 2.315 11.03 1.605 8.415 1.605 8.415 1.535 1.31 1.535 1.31 0.73 1.65 0.73 1.65 0.865 3.605 0.865 3.605 0.675 3.835 0.675 3.835 0.865 5.845 0.865 5.845 0.675 6.075 0.675 6.075 0.865 8.085 0.865 8.085 0.675 8.315 0.675 8.315 0.865 10.325 0.865 10.325 0.675 10.555 0.675 10.555 0.865 12.565 0.865 12.565 0.675 12.795 0.675 12.795 0.865 14.805 0.865 14.805 0.675 15.035 0.675 15.035 0.865 17.045 0.865 17.045 0.675 17.275 0.675 17.275 0.865 19.285 0.865 19.285 0.675 19.515 0.675 19.515 0.865 21.525 0.865 21.525 0.675 21.755 0.675 21.755 1.535 14.77 1.535 14.77 1.605 11.93 1.605 11.93 2.315 14.665 2.315 14.665 2.38 21.655 2.38 21.655 3.375 21.425 3.375 21.425 3.055 19.415 3.055 19.415 3.375 19.185 3.375 19.185 3.055 17.175 3.055 17.175 3.375 16.945 3.375 16.945 3.055 14.935 3.055 14.935 3.375 14.705 3.375 14.705 3.055 12.695 3.055 12.695 3.375 12.465 3.375 12.465 3.055 10.455 3.055 10.455 3.375 10.225 3.375 10.225 3.055 8.215 3.055 8.215 3.375 7.985 3.375 7.985 3.055 5.975 3.055 5.975 3.375 5.745 3.375 5.745 3.055 3.735 3.055 3.735 3.375 3.505 3.375 3.505 3.055 1.595 3.055 1.595 3.375 1.365 3.375  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.64 0.475 2.64 0.475 3.62 2.33 3.62 2.33 3.285 2.67 3.285 2.67 3.62 4.57 3.62 4.57 3.285 4.91 3.285 4.91 3.62 6.81 3.62 6.81 3.285 7.15 3.285 7.15 3.62 9.05 3.62 9.05 3.285 9.39 3.285 9.39 3.62 11.29 3.62 11.29 3.285 11.63 3.285 11.63 3.62 13.53 3.62 13.53 3.285 13.87 3.285 13.87 3.62 15.77 3.62 15.77 3.285 16.11 3.285 16.11 3.62 18.01 3.62 18.01 3.285 18.35 3.285 18.35 3.62 20.25 3.62 20.25 3.285 20.59 3.285 20.59 3.62 22.545 3.62 22.545 2.64 22.775 2.64 22.775 3.62 23.52 3.62 23.52 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 23.52 -0.3 23.52 0.3 22.875 0.3 22.875 1.015 22.645 1.015 22.645 0.3 20.69 0.3 20.69 0.635 20.35 0.635 20.35 0.3 18.45 0.3 18.45 0.635 18.11 0.635 18.11 0.3 16.21 0.3 16.21 0.635 15.87 0.635 15.87 0.3 13.97 0.3 13.97 0.635 13.63 0.635 13.63 0.3 11.73 0.3 11.73 0.635 11.39 0.635 11.39 0.3 9.49 0.3 9.49 0.635 9.15 0.635 9.15 0.3 7.25 0.3 7.25 0.635 6.91 0.635 6.91 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.475 0.3 0.475 1.015 0.245 1.015 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_20

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.306 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 1.76 3.015 1.76 3.015 2.12 0.41 2.12  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2024 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.36 3.41 2.36 3.41 1.525 1.365 1.525 1.365 0.53 1.595 0.53 1.595 1.29 3.41 1.29 3.41 0.53 3.835 0.53 3.835 3.39 3.41 3.39 3.41 2.68 1.595 2.68 1.595 3.39 1.365 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 2.485 3.62 2.485 2.985 2.715 2.985 2.715 3.62 4.48 3.62 4.48 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 2.715 0.3 2.715 1.055 2.485 1.055 2.485 0.3 0.475 0.3 0.475 1.16 0.245 1.16 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_3

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.74 1.95 1.74 1.95 2.15 0.37 2.15  ;
        POLYGON 3.035 1.74 4.315 1.74 4.315 2.15 3.035 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.6096 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.71 2.39 3.835 2.39 3.835 3.39 3.605 3.39 3.605 2.77 1.595 2.77 1.595 3.39 1.365 3.39 1.365 2.39 2.33 2.39 2.33 1.44 1.365 1.44 1.365 0.675 1.595 0.675 1.595 1.06 3.605 1.06 3.605 0.675 3.835 0.675 3.835 1.44 2.71 1.44  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.615 0.475 2.615 0.475 3.62 2.485 3.62 2.485 3.13 2.715 3.13 2.715 3.62 4.725 3.62 4.725 2.62 4.955 2.62 4.955 3.62 5.6 3.62 5.6 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 4.955 0.3 4.955 0.975 4.725 0.975 4.725 0.3 2.715 0.3 2.715 0.775 2.485 0.775 2.485 0.3 0.475 0.3 0.475 0.97 0.245 0.97 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__inv_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__inv_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 8.816 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.63 1.765 4.26 1.765 4.26 2.12 0.63 2.12  ;
        POLYGON 5.32 1.765 8.96 1.765 8.96 2.12 5.32 2.12  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.2192 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.95 2.375 8.315 2.375 8.315 3.38 8.085 3.38 8.085 2.68 6.075 2.68 6.075 3.38 5.845 3.38 5.845 2.675 3.835 2.675 3.835 3.38 3.605 3.38 3.605 2.675 1.595 2.675 1.595 3.38 1.365 3.38 1.365 2.375 4.57 2.375 4.57 1.535 1.365 1.535 1.365 0.675 1.595 0.675 1.595 1.235 3.605 1.235 3.605 0.675 3.835 0.675 3.835 1.235 5.845 1.235 5.845 0.675 6.075 0.675 6.075 1.235 8.085 1.235 8.085 0.675 8.315 0.675 8.315 1.535 4.95 1.535  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.655 0.475 2.655 0.475 3.62 2.485 3.62 2.485 2.95 2.715 2.95 2.715 3.62 4.725 3.62 4.725 2.95 4.955 2.95 4.955 3.62 6.965 3.62 6.965 2.95 7.195 2.95 7.195 3.62 9.205 3.62 9.205 2.65 9.435 2.65 9.435 3.62 10.08 3.62 10.08 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.435 0.3 9.435 1.015 9.205 1.015 9.205 0.3 7.195 0.3 7.195 0.995 6.965 0.995 6.965 0.3 4.955 0.3 4.955 0.995 4.725 0.995 4.725 0.3 2.715 0.3 2.715 0.995 2.485 0.995 2.485 0.3 0.475 0.3 0.475 1.015 0.245 1.015 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__inv_8

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 9.52 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.052 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 1.7 2.425 1.7 2.425 2.12 0.41 2.12  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.526 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.74 1.56 9.34 1.56 9.4 1.56 9.4 2.375 9.34 2.375 7.74 2.375  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.072725 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.53 0.99 4.92 0.99 4.92 2.93 4.53 2.93  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 2.865 1.495 2.865 1.495 3.62 5.615 3.62 5.615 3 5.845 3 5.845 3.62 6.98 3.62 7.77 3.62 7.77 3.115 8 3.115 8 3.62 9.34 3.62 9.52 3.62 9.52 4.22 9.34 4.22 6.98 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 9.52 -0.3 9.52 0.3 8 0.3 8 0.815 7.77 0.815 7.77 0.3 6.16 0.3 6.16 0.905 5.93 0.905 5.93 0.3 1.65 0.3 1.65 0.76 1.31 0.76 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.405 2.71 2.405 2.71 1.225 0.18 1.225 0.18 0.53 0.54 0.53 0.54 0.995 3.01 0.995 3.01 2.635 0.475 2.635 0.475 3.39 0.245 3.39  ;
        POLYGON 2.4 0.53 5.575 0.53 5.575 1.135 6.585 1.135 6.585 0.53 6.935 0.53 6.935 1.365 5.575 1.365 5.575 1.62 5.345 1.62 5.345 0.76 3.47 0.76 3.47 2.61 3.82 2.61 3.82 2.91 3.24 2.91 3.24 0.76 2.4 0.76  ;
        POLYGON 2.285 2.865 2.515 2.865 2.515 3.16 4.05 3.16 4.05 2.38 3.77 2.38 3.77 0.99 4.11 0.99 4.11 2.15 4.28 2.15 4.28 3.16 5.15 3.16 5.15 1.9 5.38 1.9 5.38 2.535 6.98 2.535 6.98 3.375 6.75 3.375 6.75 2.77 5.385 2.77 5.385 3.39 2.285 3.39  ;
        POLYGON 7.26 1.045 8.23 1.045 8.23 0.53 9.34 0.53 9.34 0.76 8.46 0.76 8.46 1.275 7.49 1.275 7.49 2.65 9.175 2.65 9.175 3.375 8.945 3.375 8.945 2.885 7.26 2.885  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_12
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_12 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 30.24 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.77 1.59 1.77 1.59 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.1185 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.615 1.77 8.475 1.77 8.475 2.15 4.615 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.594 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.445 2.46 22.65 2.46 23.04 2.46 23.04 1.265 20.75 1.265 20.75 1.135 17.12 1.135 17.12 0.865 28.88 0.865 28.88 1.135 26.61 1.135 26.61 1.265 23.44 1.265 23.44 2.46 28.28 2.46 28.28 3.38 28.045 3.38 28.045 2.86 26.235 2.86 26.235 3.38 26.005 3.38 26.005 2.86 24.195 2.86 24.195 3.38 23.965 3.38 23.965 2.86 22.65 2.86 22.055 2.86 22.055 3.38 21.825 3.38 21.825 2.86 19.815 2.86 19.815 3.38 19.585 3.38 19.585 2.86 17.675 2.86 17.675 3.38 17.445 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.63 3.62 1.63 3.13 1.86 3.13 1.86 3.62 6.4 3.62 6.4 3.445 6.74 3.445 6.74 3.62 9.815 3.62 9.815 3.1 10.045 3.1 10.045 3.62 12.02 3.62 12.02 2.59 12.36 2.59 12.36 3.62 14.06 3.62 14.06 2.59 14.4 2.59 14.4 3.62 16.17 3.62 16.17 2.59 16.51 2.59 16.51 3.62 18.465 3.62 18.465 3.23 18.695 3.23 18.695 3.62 20.705 3.62 20.705 3.23 20.935 3.23 20.935 3.62 22.65 3.62 22.945 3.62 22.945 3.23 23.175 3.23 23.175 3.62 24.985 3.62 24.985 3.23 25.215 3.23 25.215 3.62 27.025 3.62 27.025 3.23 27.255 3.23 27.255 3.62 28.84 3.62 29.065 3.62 29.065 2.53 29.295 2.53 29.295 3.62 29.485 3.62 30.24 3.62 30.24 4.22 29.485 4.22 28.84 4.22 22.65 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 30.24 -0.3 30.24 0.3 29.945 0.3 29.945 0.915 29.715 0.915 29.715 0.3 27.76 0.3 27.76 0.635 27.225 0.635 27.225 0.3 25.52 0.3 25.52 0.635 25.18 0.635 25.18 0.3 23.28 0.3 23.28 0.635 22.94 0.635 22.94 0.3 21.04 0.3 21.04 0.635 20.7 0.635 20.7 0.3 18.8 0.3 18.8 0.635 18.46 0.635 18.46 0.3 16.505 0.3 16.505 0.93 16.275 0.93 16.275 0.3 14.265 0.3 14.265 0.93 14.035 0.93 14.035 0.3 12.025 0.3 12.025 0.93 11.795 0.93 11.795 0.3 9.63 0.3 9.63 0.475 9.27 0.475 9.27 0.3 6.51 0.3 6.51 0.475 6.15 0.475 6.15 0.3 1.645 0.3 1.645 0.76 1.415 0.76 1.415 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.61 2.57 1.935 2.57 1.935 1.225 0.295 1.225 0.295 0.715 0.525 0.715 0.525 0.99 2.165 0.99 2.165 2.09 3.375 2.09 3.375 2.32 2.165 2.32 2.165 2.865 0.84 2.865 0.84 3.38 0.61 3.38  ;
        POLYGON 5.15 2.525 8.77 2.525 8.77 1.395 4.59 1.395 4.59 0.99 4.95 0.99 4.95 1.165 7.71 1.165 7.71 0.99 8.07 0.99 8.07 1.165 9 1.165 9 1.65 15.965 1.65 15.965 1.9 9 1.9 9 2.78 7.43 2.78 7.43 2.755 5.665 2.755 5.665 2.78 5.15 2.78  ;
        POLYGON 2.535 0.53 5.92 0.53 5.92 0.705 6.925 0.705 6.925 0.53 8.785 0.53 8.785 0.705 11.285 0.705 11.285 1.19 12.915 1.19 12.915 0.58 13.145 0.58 13.145 1.19 15.155 1.19 15.155 0.58 15.385 0.58 15.385 1.19 16.505 1.19 16.505 1.365 20.475 1.365 20.475 1.595 16.275 1.595 16.275 1.42 11.055 1.42 11.055 0.935 8.555 0.935 8.555 0.76 7.155 0.76 7.155 0.935 5.69 0.935 5.69 0.76 3.255 0.76 3.255 1.63 3.9 1.63 3.9 2.89 3.67 2.89 3.67 1.86 3.025 1.86 3.025 0.885 2.535 0.885  ;
        POLYGON 2.595 3.125 4.13 3.125 4.13 1.4 3.81 1.4 3.81 0.99 4.36 0.99 4.36 3.01 5.94 3.01 5.94 2.985 7.2 2.985 7.2 3.01 9.26 3.01 9.26 2.61 11.055 2.61 11.055 2.13 16.275 2.13 16.275 1.96 22.65 1.96 22.65 2.195 16.505 2.195 16.505 2.36 15.365 2.36 15.365 3.38 15.135 3.38 15.135 2.36 13.325 2.36 13.325 3.38 13.095 3.38 13.095 2.36 11.285 2.36 11.285 3.38 11.055 3.38 11.055 2.84 9.49 2.84 9.49 3.355 6.97 3.355 6.97 3.215 6.17 3.215 6.17 3.355 2.595 3.355  ;
        POLYGON 24.405 1.96 28.84 1.96 28.84 2.195 24.405 2.195  ;
        POLYGON 26.86 1.365 29.485 1.365 29.485 1.595 26.86 1.595  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_12

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_16
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_16 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 39.2 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.77 1.59 1.77 1.59 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.77 9.85 1.77 9.85 2.15 5.13 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 9.205 ;
    PORT
      LAYER Metal1 ;
        POLYGON 29.85 2.425 37.785 2.425 37.785 3.38 37.5 3.38 37.5 3.005 35.455 3.005 35.455 3.38 35.225 3.38 35.225 3.005 33.205 3.005 33.205 3.38 32.975 3.38 32.975 3.005 30.985 3.005 30.985 3.38 30.755 3.38 30.755 3.005 28.74 3.005 28.74 3.38 28.51 3.38 28.51 3.005 28.145 3.005 26.485 3.005 26.485 3.38 26.255 3.38 26.255 3.005 24.255 3.005 24.255 3.38 24.025 3.38 24.025 3.005 22.05 3.005 22.05 3.38 21.82 3.38 21.82 2.425 28.145 2.425 28.95 2.425 28.95 1.445 25.24 1.445 25.24 1.135 21.755 1.135 21.755 0.865 37.785 0.865 37.785 1.135 34.285 1.135 34.285 1.445 29.85 1.445  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.63 3.62 1.63 3.285 1.97 3.285 1.97 3.62 5.045 3.62 5.045 3.445 5.385 3.445 5.385 3.62 8.155 3.62 8.155 3.445 8.515 3.445 8.515 3.62 11.35 3.62 11.35 2.7 11.58 2.7 11.58 3.62 13.76 3.62 13.76 2.7 13.99 2.7 13.99 3.62 15.995 3.62 15.995 2.7 16.225 2.7 16.225 3.62 18.33 3.62 18.33 2.7 18.56 2.7 18.56 3.62 20.68 3.62 20.68 2.7 20.91 2.7 20.91 3.62 22.835 3.62 22.835 3.285 23.175 3.285 23.175 3.62 25.08 3.62 25.08 3.285 25.42 3.285 25.42 3.62 27.33 3.62 27.33 3.285 27.67 3.285 27.67 3.62 28.145 3.62 29.57 3.62 29.57 3.285 29.91 3.285 29.91 3.62 31.81 3.62 31.81 3.285 32.15 3.285 32.15 3.62 34.05 3.62 34.05 3.285 34.39 3.285 34.39 3.62 36.285 3.62 36.285 3.285 36.625 3.285 36.625 3.62 38.3 3.62 38.52 3.62 38.52 2.53 38.75 2.53 38.75 3.62 39.2 3.62 39.2 4.22 38.3 4.22 28.145 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 39.2 -0.3 39.2 0.3 38.85 0.3 38.85 1.015 38.62 1.015 38.62 0.3 36.665 0.3 36.665 0.635 36.325 0.635 36.325 0.3 34.425 0.3 34.425 0.635 34.085 0.635 34.085 0.3 32.185 0.3 32.185 0.635 31.845 0.635 31.845 0.3 29.945 0.3 29.945 0.635 29.605 0.635 29.605 0.3 27.705 0.3 27.705 0.635 27.365 0.635 27.365 0.3 25.465 0.3 25.465 0.635 25.125 0.635 25.125 0.3 23.225 0.3 23.225 0.635 22.885 0.635 22.885 0.3 20.93 0.3 20.93 0.87 20.7 0.87 20.7 0.3 18.51 0.3 18.51 0.87 18.28 0.87 18.28 0.3 16.27 0.3 16.27 0.87 16.04 0.87 16.04 0.3 14.03 0.3 14.03 0.87 13.8 0.87 13.8 0.3 11.635 0.3 11.635 0.475 11.275 0.475 11.275 0.3 8.515 0.3 8.515 0.475 8.155 0.475 8.155 0.3 5.385 0.3 5.385 0.53 5.1 0.53 5.1 0.3 1.7 0.3 1.7 0.76 1.47 0.76 1.47 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.665 2.57 2.045 2.57 2.045 1.225 0.35 1.225 0.35 0.675 0.58 0.675 0.58 0.99 2.275 0.99 2.275 2.035 3.375 2.035 3.375 2.8 0.895 2.8 0.895 3.38 0.665 3.38  ;
        POLYGON 6.31 2.525 10.175 2.525 10.175 1.42 6.595 1.42 6.595 0.99 6.955 0.99 6.955 1.19 9.715 1.19 9.715 0.99 10.415 0.99 10.415 1.63 20.325 1.63 20.325 1.96 10.405 1.96 10.405 2.78 9.315 2.78 9.315 2.755 7.125 2.755 7.125 2.78 6.31 2.78  ;
        POLYGON 2.59 0.53 4.87 0.53 4.87 0.76 6.135 0.76 6.135 0.53 7.415 0.53 7.415 0.73 9.255 0.73 9.255 0.53 11.045 0.53 11.045 0.73 13.255 0.73 13.255 1.1 14.92 1.1 14.92 0.53 15.15 0.53 15.15 1.1 17.16 1.1 17.16 0.53 17.39 0.53 17.39 1.1 19.58 1.1 19.58 0.53 19.81 0.53 19.81 1.1 20.93 1.1 20.93 1.365 24.785 1.365 24.785 1.595 20.7 1.595 20.7 1.33 13.025 1.33 13.025 0.96 10.815 0.96 10.815 0.76 9.485 0.76 9.485 0.96 7.185 0.96 7.185 0.76 6.365 0.76 6.365 0.99 4.64 0.99 4.64 0.76 3.31 0.76 3.31 1.575 3.955 1.575 3.955 2.89 3.725 2.89 3.725 1.805 3.08 1.805 3.08 0.885 2.59 0.885  ;
        POLYGON 2.59 3.12 4.185 3.12 4.185 1.345 3.865 1.345 3.865 0.99 4.225 0.99 4.225 1.115 4.415 1.115 4.415 2.985 5.845 2.985 5.845 3.01 7.385 3.01 7.385 2.985 9.085 2.985 9.085 3.01 10.815 3.01 10.815 2.19 20.7 2.19 20.7 1.96 28.145 1.96 28.145 2.195 20.93 2.195 20.93 2.425 19.75 2.425 19.75 3.38 19.52 3.38 19.52 2.425 17.355 2.425 17.355 3.38 17.125 3.38 17.125 2.425 15.11 2.425 15.11 3.38 14.88 3.38 14.88 2.425 12.86 2.425 12.86 3.38 12.63 3.38 12.63 2.425 11.045 2.425 11.045 3.355 8.855 3.355 8.855 3.215 7.615 3.215 7.615 3.355 5.615 3.355 5.615 3.215 4.815 3.215 4.815 3.35 2.59 3.35  ;
        POLYGON 34.765 1.365 38.3 1.365 38.3 1.595 34.765 1.595  ;
        POLYGON 32.315 1.96 38.3 1.96 38.3 2.195 32.315 2.195  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_16

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 9.52 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 1.625 1.59 1.625 1.59 2.125 0.41 2.125  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.082 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.405 1.16 7.77 1.16 7.77 1.64 8.775 1.64 8.775 2.19 7.405 2.19  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.04 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.795 0.53 7.175 0.53 7.175 2.8 6.88 2.8 6.88 1.66 6.795 1.66  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.465 3.62 1.465 2.815 1.805 2.815 1.805 3.62 5.925 3.62 5.925 2.89 6.155 2.89 6.155 3.62 7.965 3.62 7.965 2.98 8.195 2.98 8.195 3.62 9.285 3.62 9.52 3.62 9.52 4.22 9.285 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 9.52 -0.3 9.52 0.3 8.145 0.3 8.145 0.92 7.915 0.92 7.915 0.3 5.96 0.3 5.96 0.635 5.62 0.635 5.62 0.3 1.605 0.3 1.605 0.76 1.375 0.76 1.375 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.5 2.355 1.84 2.355 1.84 1.225 0.255 1.225 0.255 0.57 0.485 0.57 0.485 0.99 2.07 0.99 2.07 2.035 3.21 2.035 3.21 2.585 0.73 2.585 0.73 3.38 0.5 3.38  ;
        POLYGON 2.495 0.53 5.39 0.53 5.39 0.865 6.565 0.865 6.565 1.64 6.335 1.64 6.335 1.095 5.16 1.095 5.16 0.76 3.215 0.76 3.215 1.575 3.79 1.575 3.79 2.89 3.555 2.89 3.555 1.805 2.985 1.805 2.985 0.885 2.495 0.885  ;
        POLYGON 2.445 3.125 4.02 3.125 4.02 1.345 3.77 1.345 3.77 0.99 4.25 0.99 4.25 1.325 6.105 1.325 6.105 1.965 6.65 1.965 6.65 2.195 5.875 2.195 5.875 1.555 4.25 1.555 4.25 3.125 4.905 3.125 4.905 2.465 5.135 2.465 5.135 3.355 2.445 3.355  ;
        POLYGON 5.415 1.915 5.645 1.915 5.645 2.425 6.615 2.425 6.615 3.07 7.505 3.07 7.505 2.52 9.02 2.52 9.02 0.58 9.285 0.58 9.285 3.38 9.02 3.38 9.02 2.75 7.735 2.75 7.735 3.3 6.385 3.3 6.385 2.66 5.415 2.66  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_3
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_3 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.88 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.65 1.6 1.65 1.6 2.15 0.66 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.53 1.79 6.11 1.79 6.11 2.125 4.53 2.125  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.92 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.41 2.425 11.365 2.425 11.87 2.425 12.265 2.425 12.265 1.1 10.025 1.1 10.025 0.615 10.255 0.615 10.255 0.865 12.265 0.865 12.265 0.61 12.76 0.61 12.76 2.75 11.87 2.75 11.79 2.75 11.79 3.165 11.45 3.165 11.45 2.66 11.365 2.66 9.75 2.66 9.75 3.165 9.41 3.165  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.565 3.62 1.565 3.065 1.795 3.065 1.795 3.62 6.085 3.62 6.085 3.285 6.425 3.285 6.425 3.62 8.335 3.62 8.335 2.76 8.565 2.76 8.565 3.62 10.485 3.62 10.485 3.165 10.715 3.165 10.715 3.62 11.365 3.62 11.87 3.62 12.88 3.62 12.88 4.22 11.87 4.22 11.365 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.88 -0.3 12.88 0.3 11.43 0.3 11.43 0.635 11.09 0.635 11.09 0.3 8.955 0.3 8.955 0.9 8.725 0.9 8.725 0.3 6.47 0.3 6.47 0.635 6.13 0.635 6.13 0.3 1.65 0.3 1.65 0.76 1.42 0.76 1.42 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.545 2.495 1.86 2.495 1.86 1.225 0.3 1.225 0.3 0.675 0.53 0.675 0.53 0.99 2.09 0.99 2.09 2.035 3.255 2.035 3.255 2.79 0.775 2.79 0.775 3.305 0.545 3.305  ;
        POLYGON 5.025 2.355 6.745 2.355 6.745 1.56 5.12 1.56 5.12 1.22 4.7 1.22 4.7 0.99 5.35 0.99 5.35 1.325 7.97 1.325 7.97 1.555 6.975 1.555 6.975 2.59 5.255 2.59 5.255 2.87 5.025 2.87  ;
        POLYGON 2.53 3.155 4.065 3.155 4.065 1.345 3.815 1.345 3.815 0.99 4.295 0.99 4.295 3.155 5.485 3.155 5.485 2.825 7.875 2.825 7.875 1.96 11.365 1.96 11.365 2.195 8.105 2.195 8.105 3.055 5.715 3.055 5.715 3.39 2.53 3.39  ;
        POLYGON 2.54 0.53 5.81 0.53 5.81 0.865 7.395 0.865 7.395 0.53 7.625 0.53 7.625 0.865 8.43 0.865 8.43 1.365 11.87 1.365 11.87 1.595 8.2 1.595 8.2 1.095 5.58 1.095 5.58 0.76 3.26 0.76 3.26 1.575 3.835 1.575 3.835 2.89 3.6 2.89 3.6 1.805 3.03 1.805 3.03 0.885 2.54 0.885  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_3

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.76 1.62 1.76 1.62 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.475 1.79 6.07 1.79 6.07 2.135 4.475 2.135  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.08 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.11 2.425 9.95 2.425 10.125 2.425 10.73 2.425 10.73 1.1 9.4 1.1 9.4 0.715 9.63 0.715 9.63 0.865 11.64 0.865 11.64 0.71 11.87 0.71 11.87 1.1 11.11 1.1 11.11 2.425 11.42 2.425 11.42 3.38 11.19 3.38 11.19 2.66 10.125 2.66 9.95 2.66 9.41 2.66 9.41 3.38 9.11 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.455 3.62 1.455 3.285 1.795 3.285 1.795 3.62 5.985 3.62 5.985 3.285 6.325 3.285 6.325 3.62 8.075 3.62 8.075 2.815 8.415 2.815 8.415 3.62 9.95 3.62 10.125 3.62 10.17 3.62 10.17 3.02 10.4 3.02 10.4 3.62 12.21 3.62 12.21 2.565 12.44 2.565 12.44 3.62 13.44 3.62 13.44 4.22 10.125 4.22 9.95 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 12.99 0.3 12.99 1.06 12.76 1.06 12.76 0.3 10.805 0.3 10.805 0.635 10.465 0.635 10.465 0.3 8.565 0.3 8.565 0.635 8.225 0.635 8.225 0.3 6.325 0.3 6.325 0.635 5.985 0.635 5.985 0.3 1.595 0.3 1.595 0.76 1.365 0.76 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.49 2.51 1.87 2.51 1.87 1.225 0.245 1.225 0.245 0.67 0.475 0.67 0.475 0.99 2.1 0.99 2.1 2.085 3.26 2.085 3.26 2.32 2.1 2.32 2.1 2.74 0.72 2.74 0.72 3.38 0.49 3.38  ;
        POLYGON 4.89 2.365 6.6 2.365 6.6 1.56 4.935 1.56 4.935 1.22 4.515 1.22 4.515 0.99 5.165 0.99 5.165 1.325 6.83 1.325 6.83 1.73 7.94 1.73 7.94 2.125 6.83 2.125 6.83 2.595 5.12 2.595 5.12 2.89 4.89 2.89  ;
        POLYGON 2.475 3.125 4.01 3.125 4.01 1.345 3.76 1.345 3.76 0.99 4.24 0.99 4.24 3.12 5.395 3.12 5.395 2.825 7.11 2.825 7.11 2.355 8.335 2.355 8.335 1.96 9.95 1.96 9.95 2.195 8.565 2.195 8.565 2.585 7.34 2.585 7.34 3.38 7.11 3.38 7.11 3.055 5.625 3.055 5.625 3.355 2.475 3.355  ;
        POLYGON 2.485 0.53 5.625 0.53 5.625 0.865 8.565 0.865 8.565 1.365 10.125 1.365 10.125 1.595 8.335 1.595 8.335 1.095 5.395 1.095 5.395 0.76 3.205 0.76 3.205 1.575 3.78 1.575 3.78 2.89 3.545 2.89 3.545 1.805 2.975 1.805 2.975 0.885 2.485 0.885  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__invz_8
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__invz_8 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.84 BY 3.92 ;
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 1.77 1.625 1.77 1.625 2.15 0.37 2.15  ;
    END
  END EN
  PIN I
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.073 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.57 1.785 7.72 1.785 7.72 2.15 4.57 2.15  ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.2676 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.505 2.53 16.325 2.53 16.85 2.53 16.85 1.155 15.74 1.155 15.74 1.135 13.51 1.135 13.51 0.63 13.74 0.63 13.74 0.865 15.75 0.865 15.75 0.635 15.98 0.635 15.98 0.865 17.99 0.865 17.99 0.635 18.22 0.635 18.22 0.865 20.23 0.865 20.23 0.635 20.46 0.635 20.46 1.135 18.315 1.135 18.315 1.155 17.34 1.155 17.34 2.53 19.91 2.53 19.91 3.38 19.68 3.38 19.68 2.83 17.87 2.83 17.87 3.38 17.64 3.38 17.64 2.83 16.325 2.83 15.83 2.83 15.83 3.38 15.6 3.38 15.6 2.83 13.745 2.83 13.745 3.38 13.505 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.535 3.62 1.535 3.285 1.88 3.285 1.88 3.62 4.955 3.62 4.955 3.445 5.295 3.445 5.295 3.62 7.555 3.62 7.555 3.445 7.915 3.445 7.915 3.62 10.1 3.62 10.1 2.665 10.33 2.665 10.33 3.62 12.34 3.62 12.34 2.665 12.57 2.665 12.57 3.62 14.58 3.62 14.58 3.23 14.81 3.23 14.81 3.62 16.325 3.62 16.62 3.62 16.62 3.23 16.85 3.23 16.85 3.62 18.66 3.62 18.66 3.23 18.89 3.23 18.89 3.62 20.46 3.62 20.7 3.62 20.7 2.53 20.93 2.53 20.93 3.62 21.14 3.62 21.84 3.62 21.84 4.22 21.14 4.22 20.46 4.22 16.325 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 21.84 -0.3 21.84 0.3 21.58 0.3 21.58 1.015 21.35 1.015 21.35 0.3 19.395 0.3 19.395 0.635 19.055 0.635 19.055 0.3 17.155 0.3 17.155 0.635 16.815 0.635 16.815 0.3 14.915 0.3 14.915 0.635 14.575 0.635 14.575 0.3 12.62 0.3 12.62 0.865 12.39 0.865 12.39 0.3 10.38 0.3 10.38 0.865 10.15 0.865 10.15 0.3 8.195 0.3 8.195 0.635 7.855 0.635 7.855 0.3 5.295 0.3 5.295 0.53 5.01 0.53 5.01 0.3 1.61 0.3 1.61 0.76 1.38 0.76 1.38 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.575 2.57 1.955 2.57 1.955 1.225 0.26 1.225 0.26 0.675 0.49 0.675 0.49 0.99 2.185 0.99 2.185 2.09 3.345 2.09 3.345 2.32 2.185 2.32 2.185 2.8 0.805 2.8 0.805 3.38 0.575 3.38  ;
        POLYGON 6.105 2.525 8.5 2.525 8.5 1.555 6.515 1.555 6.515 0.99 6.935 0.99 6.935 1.325 8.73 1.325 8.73 1.625 12.145 1.625 12.145 1.955 8.73 1.955 8.73 2.755 6.58 2.755 6.58 2.78 6.105 2.78  ;
        POLYGON 2.5 0.53 4.78 0.53 4.78 0.76 5.77 0.76 5.77 0.53 7.395 0.53 7.395 0.865 9.03 0.865 9.03 0.53 9.26 0.53 9.26 0.865 9.635 0.865 9.635 1.095 11.27 1.095 11.27 0.53 11.5 0.53 11.5 1.095 12.62 1.095 12.62 1.365 15.48 1.365 15.48 1.595 12.39 1.595 12.39 1.325 9.405 1.325 9.405 1.095 7.165 1.095 7.165 0.76 6 0.76 6 0.99 4.55 0.99 4.55 0.76 3.22 0.76 3.22 1.575 3.865 1.575 3.865 2.89 3.635 2.89 3.635 1.805 2.99 1.805 2.99 0.885 2.5 0.885  ;
        POLYGON 2.52 3.125 4.095 3.125 4.095 1.345 3.775 1.345 3.775 0.99 4.135 0.99 4.135 1.115 4.325 1.115 4.325 2.985 5.875 2.985 5.875 3.055 6.81 3.055 6.81 2.985 9.025 2.985 9.025 2.185 12.39 2.185 12.39 1.96 16.325 1.96 16.325 2.195 12.62 2.195 12.62 2.415 11.45 2.415 11.45 3.26 11.22 3.26 11.22 2.415 9.365 2.415 9.365 3.215 7.325 3.215 7.325 3.355 5.525 3.355 5.525 3.215 4.725 3.215 4.725 3.355 2.52 3.355  ;
        POLYGON 18.165 1.96 20.46 1.96 20.46 2.195 18.165 2.195  ;
        POLYGON 18.505 1.365 21.14 1.365 21.14 1.595 18.505 1.595  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__invz_8

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 11.2 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.35 1.24 4 1.24 4 0.55 4.43 0.55 4.43 1.56 3.35 1.56  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.736 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.8 2.15 1.8 2.15 2.75 1.77 2.75 1.77 2.12 0.825 2.12  ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.605 0.53 9.96 0.53 9.96 3.38 9.605 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 2.66 1.495 2.66 1.495 3.62 2.36 3.62 3.485 3.62 3.485 3.085 3.715 3.085 3.715 3.62 5.1 3.62 7.765 3.62 7.765 2.655 7.995 2.655 7.995 3.62 9.17 3.62 10.625 3.62 10.625 2.53 10.855 2.53 10.855 3.62 11.2 3.62 11.2 4.22 9.17 4.22 5.1 4.22 2.36 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 11.2 -0.3 11.2 0.3 10.955 0.3 10.955 1.16 10.725 1.16 10.725 0.3 7.995 0.3 7.995 0.895 7.765 0.895 7.765 0.3 3.615 0.3 3.615 0.825 3.385 0.825 3.385 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.16 2.36 1.16 2.36 1.39 0.53 1.39 0.53 3.39 0.19 3.39  ;
        POLYGON 3.125 2.335 5.1 2.335 5.1 2.565 3.125 2.565  ;
        POLYGON 2.61 0.53 2.95 0.53 2.95 1.855 4.785 1.855 4.785 1.01 5.015 1.01 5.015 1.855 5.985 1.855 5.985 2.81 5.755 2.81 5.755 2.085 2.895 2.085 2.895 3.39 2.61 3.39  ;
        POLYGON 5.1 3.14 6.275 3.14 6.275 0.76 5.2 0.76 5.2 0.53 6.505 0.53 6.505 1.245 8.58 1.245 8.58 1.475 6.505 1.475 6.505 3.37 5.1 3.37  ;
        POLYGON 7.025 2.075 8.83 2.075 8.83 0.53 9.17 0.53 9.17 2.305 9.035 2.305 9.035 3.225 8.785 3.225 8.785 2.305 7.025 2.305  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.35 1.24 4 1.24 4 0.55 4.43 0.55 4.43 1.56 3.35 1.56  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.736 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.8 2.15 1.8 2.15 2.75 1.77 2.75 1.77 2.12 0.825 2.12  ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.66 0.53 11.08 0.53 11.08 3.38 10.66 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3.05 1.595 3.05 1.595 3.62 2.36 3.62 3.485 3.62 3.485 3.085 3.715 3.085 3.715 3.62 5.1 3.62 7.41 3.62 7.41 2.805 7.75 2.805 7.75 3.62 9.17 3.62 9.705 3.62 9.705 2.53 9.935 2.53 9.935 3.62 11.745 3.62 11.745 2.53 11.975 2.53 11.975 3.62 12.32 3.62 12.32 4.22 9.17 4.22 5.1 4.22 2.36 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 12.075 0.3 12.075 1.055 11.845 1.055 11.845 0.3 9.835 0.3 9.835 1.055 9.605 1.055 9.605 0.3 7.995 0.3 7.995 0.895 7.765 0.895 7.765 0.3 3.615 0.3 3.615 0.825 3.385 0.825 3.385 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.575 0.53 0.575 1.16 2.36 1.16 2.36 1.39 0.575 1.39 0.575 3.39 0.19 3.39  ;
        POLYGON 3.125 2.335 5.1 2.335 5.1 2.565 3.125 2.565  ;
        POLYGON 2.61 0.53 2.95 0.53 2.95 1.855 4.785 1.855 4.785 1.01 5.015 1.01 5.015 1.855 5.985 1.855 5.985 2.81 5.755 2.81 5.755 2.085 2.895 2.085 2.895 3.39 2.61 3.39  ;
        POLYGON 5.1 3.14 6.275 3.14 6.275 0.76 5.2 0.76 5.2 0.53 6.505 0.53 6.505 1.245 8.58 1.245 8.58 1.475 6.505 1.475 6.505 3.37 5.1 3.37  ;
        POLYGON 6.82 2.075 8.83 2.075 8.83 0.53 9.17 0.53 9.17 2.305 8.715 2.305 8.715 3.225 8.485 3.225 8.485 2.305 6.82 2.305  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.68 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.35 1.24 4 1.24 4 0.55 4.43 0.55 4.43 1.56 3.35 1.56  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.736 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.8 2.15 1.8 2.15 2.75 1.8 2.75 1.8 2.12 0.825 2.12  ;
    END
  END E
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1216 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.24 0.53 11.7 0.53 11.7 1.8 13.28 1.8 13.28 0.53 13.88 0.53 13.88 3.38 13.28 3.38 13.28 2.12 11.7 2.12 11.7 3.38 11.24 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3.05 1.595 3.05 1.595 3.62 2.36 3.62 3.485 3.62 3.485 3.085 3.715 3.085 3.715 3.62 5.1 3.62 7.705 3.62 7.705 2.805 8.05 2.805 8.05 3.62 9.17 3.62 10.225 3.62 10.225 2.53 10.455 2.53 10.455 3.62 12.265 3.62 12.265 2.53 12.495 2.53 12.495 3.62 14.305 3.62 14.305 2.53 14.535 2.53 14.535 3.62 15.68 3.62 15.68 4.22 9.17 4.22 5.1 4.22 2.36 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 15.68 -0.3 15.68 0.3 14.935 0.3 14.935 1.055 14.705 1.055 14.705 0.3 12.695 0.3 12.695 1.055 12.465 1.055 12.465 0.3 10.455 0.3 10.455 1.055 10.225 1.055 10.225 0.3 7.995 0.3 7.995 0.895 7.765 0.895 7.765 0.3 3.615 0.3 3.615 0.825 3.385 0.825 3.385 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.575 0.53 0.575 1.16 2.36 1.16 2.36 1.39 0.575 1.39 0.575 3.39 0.19 3.39  ;
        POLYGON 3.125 2.335 5.1 2.335 5.1 2.565 3.125 2.565  ;
        POLYGON 2.61 0.53 2.95 0.53 2.95 1.855 4.785 1.855 4.785 1.01 5.015 1.01 5.015 1.855 5.985 1.855 5.985 2.81 5.755 2.81 5.755 2.085 2.895 2.085 2.895 3.39 2.61 3.39  ;
        POLYGON 5.1 3.14 6.275 3.14 6.275 0.76 5.2 0.76 5.2 0.53 6.505 0.53 6.505 1.245 8.58 1.245 8.58 1.475 6.505 1.475 6.505 3.37 5.1 3.37  ;
        POLYGON 7.12 2.075 8.83 2.075 8.83 0.53 9.17 0.53 9.17 2.305 9.015 2.305 9.015 3.225 8.785 3.225 8.785 2.305 7.12 2.305  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.285 1.24 3.31 1.24 3.31 1.63 2.285 1.63  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.045 1.825 1.045 1.825 0.68 3.905 0.68 3.905 1.035 5.475 1.035 5.475 2.135 5.16 2.135 5.16 1.265 3.675 1.265 3.675 1 2.055 1 2.055 1.275 0.76 1.275  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.38 2.365 4.64 2.365 5.705 2.365 5.705 1.565 7 1.565 7 1.795 5.935 1.795 5.935 2.68 4.64 2.68 4 2.68 4 2.595 2.38 2.595  ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.53 2.53 11.88 2.53 11.88 1.12 11.31 1.12 11.31 0.6 12.19 0.6 12.19 3.38 11.53 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 2.655 1.495 2.655 1.495 3.62 2.97 3.62 2.97 3.285 3.31 3.285 3.31 3.62 6.96 3.62 6.96 3.285 7.3 3.285 7.3 3.62 8.115 3.62 10.51 3.62 10.51 2.815 10.85 2.815 10.85 3.62 11.31 3.62 12.32 3.62 12.32 4.22 11.31 4.22 8.115 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 10.515 0.3 10.515 1.075 10.285 1.075 10.285 0.3 7.555 0.3 7.555 0.875 7.325 0.875 7.325 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.905 4.64 1.905 4.64 2.135 0.475 2.135 0.475 3.31 0.19 3.31  ;
        POLYGON 2.005 2.825 3.79 2.825 3.79 3.105 6.195 3.105 6.195 2.825 7.775 2.825 7.775 2.25 8.115 2.25 8.115 3.055 6.445 3.055 6.445 3.335 3.56 3.335 3.56 3.055 2.235 3.055 2.235 3.39 2.005 3.39  ;
        POLYGON 4.29 0.53 7.095 0.53 7.095 1.105 8.17 1.105 8.17 1.335 6.865 1.335 6.865 0.76 4.29 0.76  ;
        POLYGON 6.165 2.195 7.315 2.195 7.315 1.79 8.445 1.79 8.445 0.55 8.675 0.55 8.675 1.79 10.005 1.79 10.005 2.02 8.575 2.02 8.575 3.39 8.345 3.39 8.345 2.02 7.545 2.02 7.545 2.535 6.165 2.535  ;
        POLYGON 9.165 2.34 10.345 2.34 10.345 1.535 9.165 1.535 9.165 0.735 9.395 0.735 9.395 1.305 10.575 1.305 10.575 1.79 11.31 1.79 11.31 2.02 10.575 2.02 10.575 2.57 9.395 2.57 9.395 3.25 9.165 3.25  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.285 1.24 3.31 1.24 3.31 1.63 2.285 1.63  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.045 1.825 1.045 1.825 0.68 3.905 0.68 3.905 1.035 5.475 1.035 5.475 2.135 5.16 2.135 5.16 1.265 3.675 1.265 3.675 1 2.055 1 2.055 1.275 0.76 1.275  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.38 2.365 4.64 2.365 5.705 2.365 5.705 1.565 7 1.565 7 1.795 5.935 1.795 5.935 2.68 4.64 2.68 4 2.68 4 2.595 2.38 2.595  ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.53 2.53 11.65 2.53 11.9 2.53 11.9 1.12 11.31 1.12 11.31 0.6 12.22 0.6 12.22 3.38 11.65 3.38 11.53 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 2.655 1.495 2.655 1.495 3.62 2.97 3.62 2.97 3.285 3.31 3.285 3.31 3.62 6.96 3.62 6.96 3.285 7.3 3.285 7.3 3.62 8.115 3.62 10.51 3.62 10.51 2.815 10.85 2.815 10.85 3.62 11.65 3.62 12.605 3.62 12.605 2.53 12.835 2.53 12.835 3.62 13.44 3.62 13.44 4.22 11.65 4.22 8.115 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 12.935 0.3 12.935 1.075 12.705 1.075 12.705 0.3 10.515 0.3 10.515 1.075 10.285 1.075 10.285 0.3 7.555 0.3 7.555 0.875 7.325 0.875 7.325 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.905 4.64 1.905 4.64 2.135 0.475 2.135 0.475 3.31 0.19 3.31  ;
        POLYGON 2.005 2.825 3.79 2.825 3.79 3.105 6.195 3.105 6.195 2.825 7.775 2.825 7.775 2.25 8.115 2.25 8.115 3.055 6.445 3.055 6.445 3.335 3.56 3.335 3.56 3.055 2.235 3.055 2.235 3.39 2.005 3.39  ;
        POLYGON 4.29 0.53 7.095 0.53 7.095 1.105 8.17 1.105 8.17 1.335 6.865 1.335 6.865 0.76 4.29 0.76  ;
        POLYGON 6.165 2.195 7.315 2.195 7.315 1.79 8.445 1.79 8.445 0.55 8.675 0.55 8.675 1.79 9.89 1.79 9.89 2.02 8.575 2.02 8.575 3.39 8.345 3.39 8.345 2.02 7.545 2.02 7.545 2.535 6.165 2.535  ;
        POLYGON 9.165 2.34 10.345 2.34 10.345 1.545 9.165 1.545 9.165 0.735 9.395 0.735 9.395 1.315 10.575 1.315 10.575 1.69 11.65 1.69 11.65 2.03 10.575 2.03 10.575 2.57 9.395 2.57 9.395 3.25 9.165 3.25  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.36 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.285 1.24 3.31 1.24 3.31 1.63 2.285 1.63  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.045 1.825 1.045 1.825 0.68 3.905 0.68 3.905 1.035 5.475 1.035 5.475 2.135 5.16 2.135 5.16 1.265 3.675 1.265 3.675 1 2.055 1 2.055 1.275 0.76 1.275  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.38 2.365 4.64 2.365 5.705 2.365 5.705 1.565 7 1.565 7 1.795 5.935 1.795 5.935 2.68 4.64 2.68 4 2.68 4 2.595 2.38 2.595  ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1216 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.205 2.355 14.99 2.355 15.24 2.355 15.24 1.56 13.105 1.56 13.105 0.55 13.335 0.55 13.335 1.24 15.24 1.24 15.24 0.55 15.59 0.55 15.59 3.38 15.24 3.38 15.24 2.585 14.99 2.585 13.435 2.585 13.435 3.38 13.205 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 2.655 1.495 2.655 1.495 3.62 2.97 3.62 2.97 3.285 3.31 3.285 3.31 3.62 6.96 3.62 6.96 3.285 7.3 3.285 7.3 3.62 8.215 3.62 9.565 3.62 9.565 2.655 9.795 2.655 9.795 3.62 11.65 3.62 11.65 2.815 11.99 2.815 11.99 3.62 14.17 3.62 14.17 2.815 14.51 2.815 14.51 3.62 14.99 3.62 16.21 3.62 16.21 2.625 16.55 2.625 16.55 3.62 17.36 3.62 17.36 4.22 14.99 4.22 8.215 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.36 -0.3 17.36 0.3 16.695 0.3 16.695 0.93 16.465 0.93 16.465 0.3 14.455 0.3 14.455 0.89 14.225 0.89 14.225 0.3 12.035 0.3 12.035 0.89 11.805 0.89 11.805 0.3 9.795 0.3 9.795 0.89 9.565 0.89 9.565 0.3 7.555 0.3 7.555 0.875 7.325 0.875 7.325 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.905 4.64 1.905 4.64 2.135 0.475 2.135 0.475 3.31 0.19 3.31  ;
        POLYGON 4.29 0.53 7.095 0.53 7.095 1.105 8.17 1.105 8.17 1.335 6.865 1.335 6.865 0.76 4.29 0.76  ;
        POLYGON 2.005 2.825 3.79 2.825 3.79 3.105 6.195 3.105 6.195 2.825 7.875 2.825 7.875 2.25 8.215 2.25 8.215 3.055 6.445 3.055 6.445 3.335 3.56 3.335 3.56 3.055 2.235 3.055 2.235 3.39 2.005 3.39  ;
        POLYGON 6.165 2.195 7.315 2.195 7.315 1.79 8.445 1.79 8.445 0.55 8.675 0.55 8.675 1.79 11.56 1.79 11.56 2.02 8.675 2.02 8.675 3.25 8.445 3.25 8.445 2.02 7.545 2.02 7.545 2.535 6.165 2.535  ;
        POLYGON 10.685 2.315 11.805 2.315 11.805 1.51 10.685 1.51 10.685 0.55 10.915 0.55 10.915 1.28 12.035 1.28 12.035 1.805 14.99 1.805 14.99 2.035 12.035 2.035 12.035 2.545 10.915 2.545 10.915 3.29 10.685 3.29  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.285 1.24 3.31 1.24 3.31 1.63 2.285 1.63  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.045 1.825 1.045 1.825 0.68 3.905 0.68 3.905 1.035 5.475 1.035 5.475 2.135 5.16 2.135 5.16 1.265 3.675 1.265 3.675 1 2.055 1 2.055 1.275 0.76 1.275  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.38 2.365 4.64 2.365 5.705 2.365 5.705 1.565 7 1.565 7 1.795 5.935 1.795 5.935 2.68 4.64 2.68 4 2.68 4 2.595 2.38 2.595  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.01 1.085 9.4 1.085 9.4 2.355 9.01 2.355  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.65 2.53 13 2.53 13 1.12 12.43 1.12 12.43 0.6 13.31 0.6 13.31 3.38 12.65 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 2.655 1.495 2.655 1.495 3.62 2.97 3.62 2.97 3.285 3.31 3.285 3.31 3.62 6.96 3.62 6.96 3.285 7.3 3.285 7.3 3.62 8.115 3.62 9.545 3.62 9.545 2.655 9.775 2.655 9.775 3.62 11.63 3.62 11.63 2.815 11.97 2.815 11.97 3.62 12.43 3.62 13.44 3.62 13.44 4.22 12.43 4.22 8.115 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 11.635 0.3 11.635 1.075 11.405 1.075 11.405 0.3 7.555 0.3 7.555 0.875 7.325 0.875 7.325 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.905 4.64 1.905 4.64 2.135 0.475 2.135 0.475 3.31 0.19 3.31  ;
        POLYGON 4.29 0.53 7.095 0.53 7.095 1.105 8.115 1.105 8.115 1.335 6.865 1.335 6.865 0.76 4.29 0.76  ;
        POLYGON 2.005 2.825 3.79 2.825 3.79 3.105 6.195 3.105 6.195 2.825 7.775 2.825 7.775 2.25 8.115 2.25 8.115 3.055 6.445 3.055 6.445 3.335 3.56 3.335 3.56 3.055 2.235 3.055 2.235 3.39 2.005 3.39  ;
        POLYGON 6.165 2.195 7.315 2.195 7.315 1.79 8.525 1.79 8.525 0.605 9.99 0.605 9.99 1.79 11.125 1.79 11.125 2.02 9.76 2.02 9.76 0.835 8.755 0.835 8.755 3.39 8.525 3.39 8.525 2.02 7.545 2.02 7.545 2.535 6.165 2.535  ;
        POLYGON 10.285 2.34 11.465 2.34 11.465 1.535 10.285 1.535 10.285 0.735 10.515 0.735 10.515 1.305 11.695 1.305 11.695 1.79 12.43 1.79 12.43 2.02 11.695 2.02 11.695 2.57 10.515 2.57 10.515 3.25 10.285 3.25  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrsnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.285 1.24 3.31 1.24 3.31 1.63 2.285 1.63  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.045 1.825 1.045 1.825 0.68 3.905 0.68 3.905 1.035 5.475 1.035 5.475 2.135 5.16 2.135 5.16 1.265 3.675 1.265 3.675 1 2.055 1 2.055 1.275 0.76 1.275  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.38 2.365 4.64 2.365 5.705 2.365 5.705 1.565 6.78 1.565 6.78 1.795 5.935 1.795 5.935 2.68 4.64 2.68 4 2.68 4 2.595 2.38 2.595  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.84 1.085 9.4 1.085 9.4 2.355 8.84 2.355  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.38 2.15 12.745 2.15 12.98 2.15 12.98 1.365 12.38 1.365 12.38 0.545 12.76 0.545 12.76 1.135 13.34 1.135 13.34 2.38 12.76 2.38 12.76 3.38 12.745 3.38 12.38 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 2.655 1.495 2.655 1.495 3.62 2.97 3.62 2.97 3.285 3.31 3.285 3.31 3.62 6.96 3.62 6.96 3.285 7.3 3.285 7.3 3.62 7.875 3.62 9.345 3.62 9.345 2.655 9.575 2.655 9.575 3.62 11.21 3.62 11.21 2.63 11.55 2.63 11.55 3.62 12.745 3.62 13.35 3.62 13.35 2.63 13.69 2.63 13.69 3.62 14 3.62 14 4.22 12.745 4.22 7.875 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14 -0.3 14 0.3 13.735 0.3 13.735 0.885 13.505 0.885 13.505 0.3 11.495 0.3 11.495 0.885 11.265 0.885 11.265 0.3 7.555 0.3 7.555 0.875 7.325 0.875 7.325 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.905 4.64 1.905 4.64 2.135 0.475 2.135 0.475 3.31 0.19 3.31  ;
        POLYGON 2.005 2.825 3.79 2.825 3.79 3.105 6.195 3.105 6.195 2.825 7.535 2.825 7.535 2.25 7.875 2.25 7.875 3.055 6.445 3.055 6.445 3.335 3.56 3.335 3.56 3.055 2.235 3.055 2.235 3.39 2.005 3.39  ;
        POLYGON 4.29 0.53 7.095 0.53 7.095 1.105 8.095 1.105 8.095 1.335 6.865 1.335 6.865 0.76 4.29 0.76  ;
        POLYGON 6.165 2.195 7.03 2.195 7.03 1.79 8.325 1.79 8.325 0.605 9.895 0.605 9.895 1.67 10.985 1.67 10.985 1.9 9.665 1.9 9.665 0.835 8.555 0.835 8.555 3.39 8.325 3.39 8.325 2.02 7.28 2.02 7.28 2.535 6.165 2.535  ;
        POLYGON 10.245 2.15 11.325 2.15 11.325 1.365 10.145 1.365 10.145 0.545 10.375 0.545 10.375 1.135 11.555 1.135 11.555 1.67 12.745 1.67 12.745 1.9 11.555 1.9 11.555 2.38 10.475 2.38 10.475 3.38 10.245 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrsnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.36 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.285 1.24 3.31 1.24 3.31 1.63 2.285 1.63  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.045 1.825 1.045 1.825 0.68 3.905 0.68 3.905 1.035 5.475 1.035 5.475 2.135 5.16 2.135 5.16 1.265 3.675 1.265 3.675 1 2.055 1 2.055 1.275 0.76 1.275  ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.789 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.38 2.365 4.64 2.365 5.705 2.365 5.705 1.565 6.78 1.565 6.78 1.795 5.935 1.795 5.935 2.68 4.64 2.68 4 2.68 4 2.595 2.38 2.595  ;
    END
  END RN
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.84 1.085 9.4 1.085 9.4 2.355 8.84 2.355  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1216 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.54 2.34 16.05 2.34 16.35 2.34 16.35 1.465 13.505 1.465 13.505 0.545 13.735 0.545 13.735 1.16 15.745 1.16 15.745 0.545 15.975 0.545 15.975 1.16 16.68 1.16 16.68 2.57 16.14 2.57 16.14 3.38 16.05 3.38 15.645 3.38 15.645 2.57 13.9 2.57 13.9 3.38 13.54 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.265 3.62 1.265 2.655 1.495 2.655 1.495 3.62 2.97 3.62 2.97 3.285 3.31 3.285 3.31 3.62 6.96 3.62 6.96 3.285 7.3 3.285 7.3 3.62 7.875 3.62 9.345 3.62 9.345 2.655 9.575 2.655 9.575 3.62 10.245 3.62 10.245 2.53 10.475 2.53 10.475 3.62 12.38 3.62 12.38 2.815 12.72 2.815 12.72 3.62 14.57 3.62 14.57 2.815 14.91 2.815 14.91 3.62 16.05 3.62 16.61 3.62 16.61 2.815 16.95 2.815 16.95 3.62 17.36 3.62 17.36 4.22 16.05 4.22 7.875 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.36 -0.3 17.36 0.3 17.095 0.3 17.095 0.885 16.865 0.885 16.865 0.3 14.855 0.3 14.855 0.885 14.625 0.885 14.625 0.3 12.615 0.3 12.615 0.885 12.385 0.885 12.385 0.3 10.375 0.3 10.375 0.885 10.145 0.885 10.145 0.3 7.555 0.3 7.555 0.875 7.325 0.875 7.325 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.905 4.64 1.905 4.64 2.135 0.475 2.135 0.475 3.31 0.19 3.31  ;
        POLYGON 2.005 2.825 3.79 2.825 3.79 3.105 6.195 3.105 6.195 2.825 7.535 2.825 7.535 2.25 7.875 2.25 7.875 3.055 6.445 3.055 6.445 3.335 3.56 3.335 3.56 3.055 2.235 3.055 2.235 3.39 2.005 3.39  ;
        POLYGON 4.29 0.53 7.095 0.53 7.095 1.105 8.095 1.105 8.095 1.335 6.865 1.335 6.865 0.76 4.29 0.76  ;
        POLYGON 6.165 2.195 7.03 2.195 7.03 1.79 8.325 1.79 8.325 0.605 9.895 0.605 9.895 1.715 12.04 1.715 12.04 1.945 9.665 1.945 9.665 0.835 8.555 0.835 8.555 3.39 8.325 3.39 8.325 2.02 7.28 2.02 7.28 2.535 6.165 2.535  ;
        POLYGON 11.265 2.34 12.345 2.34 12.345 1.465 11.265 1.465 11.265 0.545 11.495 0.545 11.495 1.235 12.575 1.235 12.575 1.715 16.05 1.715 16.05 1.945 12.575 1.945 12.575 2.57 11.495 2.57 11.495 3.38 11.265 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latrsnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 11.76 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.965 1.79 3.27 1.79 3.27 2.12 0.965 2.12  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.78 1.24 4.045 1.24 4.045 2.795 3.5 2.795 3.5 1.56 0.78 1.56  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.04 1.8 6.53 1.8 7.38 1.8 7.38 2.12 6.53 2.12 5.04 2.12  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.895 2.53 11.32 2.53 11.32 1.065 10.75 1.065 10.75 0.6 11.63 0.6 11.63 3.38 10.895 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.21 3.62 1.21 2.815 1.55 2.815 1.55 3.62 3.16 3.62 5.365 3.62 5.365 3 5.595 3 5.595 3.62 7.63 3.62 7.63 2.815 7.97 2.815 7.97 3.62 10.005 3.62 10.005 2.53 10.235 2.53 10.235 3.62 10.75 3.62 11.76 3.62 11.76 4.22 10.75 4.22 3.16 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 11.76 -0.3 11.76 0.3 9.955 0.3 9.955 1.075 9.725 1.075 9.725 0.3 5.695 0.3 5.695 0.86 5.465 0.86 5.465 0.3 1.595 0.3 1.595 0.86 1.365 0.86 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 2.35 3.16 2.35 3.16 2.58 0.53 2.58 0.53 3.38 0.19 3.38  ;
        POLYGON 3.16 3.095 4.32 3.095 4.32 0.76 3.41 0.76 3.41 0.53 4.56 0.53 4.56 1.225 6.53 1.225 6.53 1.455 4.56 1.455 4.56 3.325 3.16 3.325  ;
        POLYGON 4.81 2.35 7.63 2.35 7.63 0.53 7.97 0.53 7.97 1.805 9.285 1.805 9.285 2.145 7.97 2.145 7.97 2.58 6.895 2.58 6.895 3.38 6.665 3.38 6.665 2.58 4.81 2.58  ;
        POLYGON 8.605 2.395 9.525 2.395 9.525 1.555 8.605 1.555 8.605 0.735 8.835 0.735 8.835 1.325 9.755 1.325 9.755 1.79 10.75 1.79 10.75 2.02 9.755 2.02 9.755 2.625 8.835 2.625 8.835 3.25 8.605 3.25  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latsnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.965 1.79 3.27 1.79 3.27 2.12 0.965 2.12  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.78 1.24 4.045 1.24 4.045 2.795 3.5 2.795 3.5 1.56 0.78 1.56  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.04 1.8 6.53 1.8 7.38 1.8 7.38 2.12 6.53 2.12 5.04 2.12  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.64 2.11 10.935 2.11 11.3 2.11 11.3 1.38 10.64 1.38 10.64 0.555 11.1 0.555 11.1 1.13 11.66 1.13 11.66 2.34 11.1 2.34 11.1 3.38 10.935 3.38 10.64 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3 1.595 3 1.595 3.62 3.16 3.62 5.365 3.62 5.365 3 5.595 3 5.595 3.62 7.63 3.62 7.63 2.815 7.97 2.815 7.97 3.62 9.525 3.62 9.525 2.57 9.755 2.57 9.755 3.62 10.935 3.62 11.665 3.62 11.665 2.57 11.895 2.57 11.895 3.62 12.32 3.62 12.32 4.22 10.935 4.22 3.16 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 11.995 0.3 11.995 0.895 11.765 0.895 11.765 0.3 9.755 0.3 9.755 0.895 9.525 0.895 9.525 0.3 5.695 0.3 5.695 0.86 5.465 0.86 5.465 0.3 1.595 0.3 1.595 0.86 1.365 0.86 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 2.35 3.16 2.35 3.16 2.58 0.575 2.58 0.575 3.38 0.19 3.38  ;
        POLYGON 3.16 3.095 4.32 3.095 4.32 0.76 3.41 0.76 3.41 0.53 4.56 0.53 4.56 1.225 6.53 1.225 6.53 1.455 4.56 1.455 4.56 3.325 3.16 3.325  ;
        POLYGON 4.81 2.35 7.63 2.35 7.63 0.53 7.97 0.53 7.97 1.63 9.245 1.63 9.245 1.86 7.97 1.86 7.97 2.58 6.895 2.58 6.895 3.38 6.665 3.38 6.665 2.58 4.81 2.58  ;
        POLYGON 8.505 2.11 9.585 2.11 9.585 1.38 8.405 1.38 8.405 0.555 8.635 0.555 8.635 1.15 9.815 1.15 9.815 1.63 10.935 1.63 10.935 1.86 9.815 1.86 9.815 2.34 8.735 2.34 8.735 3.38 8.505 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latsnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__latsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__latsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.68 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.552 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.01 1.24 2.325 1.24 2.325 0.55 2.7 0.55 2.7 1.59 2.01 1.59  ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 1.2935 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.78 1.82 2.95 1.82 2.95 1.27 3.21 1.27 3.21 1.82 4.045 1.82 4.045 2.795 3.49 2.795 3.49 2.12 0.78 2.12  ;
    END
  END E
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.04 1.8 6.53 1.8 7.39 1.8 7.39 2.12 6.53 2.12 5.04 2.12  ;
    END
  END SETN
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1216 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.86 2.11 14.37 2.11 14.67 2.11 14.67 1.39 11.825 1.39 11.825 0.545 12.055 0.545 12.055 1.16 14.065 1.16 14.065 0.545 14.295 0.545 14.295 1.16 15 1.16 15 2.34 14.46 2.34 14.46 3.38 14.37 3.38 13.965 3.38 13.965 2.34 12.22 2.34 12.22 3.38 11.86 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 3 1.595 3 1.595 3.62 3.16 3.62 5.59 3.62 5.59 2.815 5.93 2.815 5.93 3.62 7.63 3.62 7.63 2.815 7.97 2.815 7.97 3.62 8.565 3.62 8.565 2.57 8.795 2.57 8.795 3.62 10.755 3.62 10.755 2.57 10.985 2.57 10.985 3.62 12.945 3.62 12.945 2.57 13.175 2.57 13.175 3.62 14.37 3.62 14.985 3.62 14.985 2.57 15.215 2.57 15.215 3.62 15.68 3.62 15.68 4.22 14.37 4.22 3.16 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 15.68 -0.3 15.68 0.3 15.415 0.3 15.415 0.885 15.185 0.885 15.185 0.3 13.175 0.3 13.175 0.885 12.945 0.885 12.945 0.3 10.935 0.3 10.935 0.885 10.705 0.885 10.705 0.3 8.695 0.3 8.695 0.885 8.465 0.885 8.465 0.3 5.75 0.3 5.75 1.065 5.41 1.065 5.41 0.3 1.595 0.3 1.595 1.115 1.365 1.115 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.815 0.53 0.815 0.53 2.35 3.16 2.35 3.16 2.58 0.575 2.58 0.575 3.38 0.19 3.38  ;
        POLYGON 3.16 3.095 4.32 3.095 4.32 1.06 3.45 1.06 3.45 0.83 4.56 0.83 4.56 1.34 6.53 1.34 6.53 1.57 4.56 1.57 4.56 3.325 3.16 3.325  ;
        POLYGON 4.81 2.35 7.63 2.35 7.63 0.53 7.97 0.53 7.97 1.63 10.36 1.63 10.36 1.86 7.97 1.86 7.97 2.58 6.895 2.58 6.895 3.38 6.665 3.38 6.665 2.58 4.81 2.58  ;
        POLYGON 9.585 2.11 10.665 2.11 10.665 1.39 9.585 1.39 9.585 0.545 9.815 0.545 9.815 1.16 10.895 1.16 10.895 1.63 14.37 1.63 14.37 1.86 10.895 1.86 10.895 2.34 9.815 2.34 9.815 3.38 9.585 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__latsnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.28 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5235 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.01 1.77 6.07 1.77 6.07 2.12 4.01 2.12  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5235 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.33 1.21 2.71 1.21 2.71 2.71 2.33 2.71  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.047 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.94 1.445 3.295 1.445 3.295 2.36 6.09 2.36 6.09 2.785 2.94 2.785  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.13 0.65 0.575 0.65 0.575 3.27 0.13 3.27  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.365 3.62 1.365 2.76 1.595 2.76 1.595 3.62 3.89 3.62 5.31 3.62 5.31 3.105 5.65 3.105 5.65 3.62 6.815 3.62 7.28 3.62 7.28 4.22 6.815 4.22 3.89 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.28 -0.3 7.28 0.3 5.695 0.3 5.695 0.88 5.465 0.88 5.465 0.3 1.595 0.3 1.595 0.865 1.365 0.865 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.055 3.11 3.89 3.11 3.89 3.34 1.825 3.34 1.825 1.625 0.84 1.625 0.84 1.39 1.825 1.39 1.825 0.575 3.88 0.575 3.88 0.815 2.055 0.815  ;
        POLYGON 4.125 1.145 6.35 1.145 6.35 0.53 6.815 0.53 6.815 3.38 6.35 3.38 6.35 1.375 4.125 1.375  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux2_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.4 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.575 1.25 7.225 1.25 7.225 1.58 5.575 1.58  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.88 1.545 3.23 1.545 3.23 3.285 2.88 3.285  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.92 1.25 5.22 1.25 5.22 1.81 7.37 1.81 7.37 2.195 4.91 2.195 4.91 1.65 3.92 1.65  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1218 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.25 0.54 1.65 0.54 1.65 3.38 1.25 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.295 3.62 0.295 2.53 0.525 2.53 0.525 3.62 2.385 3.62 2.385 2.53 2.615 2.53 2.615 3.62 5.26 3.62 6.59 3.62 6.59 2.965 6.93 2.965 6.93 3.62 8.05 3.62 8.4 3.62 8.4 4.22 8.05 4.22 5.26 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.4 -0.3 8.4 0.3 6.875 0.3 6.875 0.835 6.645 0.835 6.645 0.3 2.715 0.3 2.715 0.835 2.485 0.835 2.485 0.3 0.475 0.3 0.475 0.835 0.245 0.835 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 3.69 2.965 5.26 2.965 5.26 3.195 3.46 3.195 3.46 1.315 2.175 1.315 2.175 1.78 1.945 1.78 1.945 1.085 3.46 1.085 3.46 0.55 4.82 0.55 4.82 0.78 3.69 0.78  ;
        POLYGON 4.32 1.96 4.66 1.96 4.66 2.49 7.71 2.49 7.71 0.54 8.05 0.54 8.05 3.39 7.665 3.39 7.665 2.725 4.32 2.725  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux2_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.64 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.89 1.25 9.54 1.25 9.54 1.58 7.89 1.58  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.15 1.545 5.5 1.545 5.5 3.285 5.15 3.285  ;
    END
  END I1
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.255 1.25 7.59 1.25 7.59 1.81 9.635 1.81 9.635 2.195 7.28 2.195 7.28 1.65 6.255 1.65  ;
    END
  END S
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3046 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.25 0.54 1.705 0.54 1.705 1.8 3.49 1.8 3.49 0.54 3.945 0.54 3.945 3.38 3.49 3.38 3.49 2.12 1.705 2.12 1.705 3.38 1.25 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.35 3.62 0.35 2.53 0.58 2.53 0.58 3.62 2.49 3.62 2.49 2.53 2.72 2.53 2.72 3.62 4.68 3.62 4.68 2.53 4.91 2.53 4.91 3.62 7.555 3.62 8.885 3.62 8.885 2.955 9.225 2.955 9.225 3.62 10.345 3.62 10.64 3.62 10.64 4.22 10.345 4.22 7.555 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.64 -0.3 10.64 0.3 9.17 0.3 9.17 0.835 8.94 0.835 8.94 0.3 5.01 0.3 5.01 0.835 4.78 0.835 4.78 0.3 2.77 0.3 2.77 0.835 2.54 0.835 2.54 0.3 0.53 0.3 0.53 0.835 0.3 0.835 0.3 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 5.985 2.965 7.555 2.965 7.555 3.195 5.755 3.195 5.755 1.315 4.47 1.315 4.47 1.78 4.24 1.78 4.24 1.085 5.755 1.085 5.755 0.55 7.115 0.55 7.115 0.78 5.985 0.78  ;
        POLYGON 6.615 1.96 6.955 1.96 6.955 2.49 10.005 2.49 10.005 0.54 10.345 0.54 10.345 3.39 9.96 3.39 9.96 2.725 6.615 2.725  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux2_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.92 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5015 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.25 1.75 15.275 1.75 16.94 1.75 16.94 2.12 15.275 2.12 15.25 2.12  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5015 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.59 1.78 12.5 1.78 12.5 2.13 10.59 2.13  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5015 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.97 1.01 0.97 1.01 2.95 0.705 2.95  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5015 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.3 1.375 4.585 1.375 4.585 1.8 5.55 1.8 5.55 2.15 4.3 2.15  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.185 1.8 3.2 1.8 3.2 1.24 3.495 1.24 3.495 2.12 2.415 2.12 2.415 2.465 2.185 2.465  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.003 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.96 1.165 8.3 1.165 8.3 1.77 8.76 1.77 9.3 1.77 9.3 2.465 9.07 2.465 9.07 2.15 8.76 2.15 7.96 2.15  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.5104 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.65 0.6 6.38 0.6 6.38 2.855 5.99 2.855 5.99 1.57 5.65 1.57  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.685 0.475 2.685 0.475 3.62 1.65 3.62 4.845 3.62 4.845 2.845 5.185 2.845 5.185 3.62 7.27 3.62 8.76 3.62 11.67 3.62 11.67 2.845 12.015 2.845 12.015 3.62 14.1 3.62 15.955 3.62 15.955 2.815 16.295 2.815 16.295 3.62 17.46 3.62 17.92 3.62 17.92 4.22 17.46 4.22 14.1 4.22 8.76 4.22 7.27 4.22 1.65 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.92 -0.3 17.92 0.3 16.34 0.3 16.34 1.145 16.11 1.145 16.11 0.3 11.86 0.3 11.86 1.145 11.63 1.145 11.63 0.3 5.08 0.3 5.08 1.16 4.85 1.16 4.85 0.3 0.475 0.3 0.475 1.13 0.245 1.13 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.26 0.845 1.65 0.845 1.65 1.075 1.495 1.075 1.495 3.025 1.26 3.025  ;
        POLYGON 3.725 0.78 4.07 0.78 4.07 2.87 3.725 2.87  ;
        POLYGON 6.86 2.665 7.27 2.665 7.27 3.005 6.86 3.005 6.86 3.39 5.52 3.39 5.52 2.615 4.53 2.615 4.53 3.33 2.635 3.33 2.635 2.97 1.725 2.97 1.725 1.34 2.04 1.34 2.04 0.845 2.77 0.845 2.77 1.075 2.29 1.075 2.29 1.57 1.955 1.57 1.955 2.74 2.975 2.74 2.975 3.1 4.3 3.1 4.3 2.38 5.75 2.38 5.75 3.155 6.63 3.155 6.63 0.79 7.27 0.79 7.27 1.13 6.86 1.13  ;
        POLYGON 7.09 1.46 7.5 1.46 7.5 0.53 8.76 0.53 8.76 1.145 8.53 1.145 8.53 0.76 7.73 0.76 7.73 2.72 8.755 2.72 8.755 2.95 7.5 2.95 7.5 1.82 7.09 1.82  ;
        POLYGON 10.35 2.575 10.84 2.575 10.84 2.925 10.11 2.925 10.11 0.795 10.84 0.795 10.84 1.145 10.35 1.145  ;
        POLYGON 12.75 0.78 12.98 0.78 12.98 2.925 12.75 2.925  ;
        POLYGON 9.65 0.78 9.88 0.78 9.88 3.16 11.125 3.16 11.125 2.38 12.495 2.38 12.495 3.16 13.77 3.16 13.77 0.78 14.1 0.78 14.1 3.39 12.265 3.39 12.265 2.615 11.355 2.615 11.355 3.39 9.65 3.39  ;
        POLYGON 14.33 0.85 15.275 0.85 15.275 1.08 14.56 1.08 14.56 2.815 15.19 2.815 15.19 3.045 14.33 3.045  ;
        POLYGON 14.79 1.685 15.02 1.685 15.02 2.355 17.23 2.355 17.23 0.78 17.46 0.78 17.46 3.14 17.125 3.14 17.125 2.585 14.79 2.585  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux4_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.04 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5165 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.485 1.78 16.51 1.78 18.175 1.78 18.175 2.12 16.51 2.12 16.485 2.12  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5165 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.835 1.78 13.735 1.78 13.735 2.13 11.835 2.13  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.97 1.01 0.97 1.01 2.95 0.705 2.95  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.505 0.55 4.935 0.55 4.935 1.8 5.755 1.8 5.755 2.15 4.505 2.15  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.651 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.255 1.8 3.3 1.8 3.3 1.24 3.7 1.24 3.7 2.25 2.255 2.25  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.17 1.305 9.535 1.305 9.535 1.77 9.95 1.77 10.535 1.77 10.535 3.32 10.165 3.32 10.165 2.15 9.95 2.15 9.17 2.15  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.7592 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.23 0.6 6.6 0.6 6.6 2.855 6.23 2.855  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.575 0.475 2.575 0.475 3.62 1.65 3.62 5.01 3.62 5.01 2.845 5.35 2.845 5.35 3.62 7.405 3.62 7.405 2.57 7.635 2.57 7.635 3.62 8.48 3.62 9.95 3.62 12.905 3.62 12.905 2.845 13.25 2.845 13.25 3.62 15.335 3.62 17.19 3.62 17.19 2.815 17.53 2.815 17.53 3.62 18.695 3.62 19.04 3.62 19.04 4.22 18.695 4.22 15.335 4.22 9.95 4.22 8.48 4.22 1.65 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.04 -0.3 19.04 0.3 17.575 0.3 17.575 1.145 17.345 1.145 17.345 0.3 13.095 0.3 13.095 1.145 12.865 1.145 12.865 0.3 7.635 0.3 7.635 1.16 7.405 1.16 7.405 0.3 5.395 0.3 5.395 1.16 5.165 1.16 5.165 0.3 0.475 0.3 0.475 1.13 0.245 1.13 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.26 0.845 1.65 0.845 1.65 1.075 1.495 1.075 1.495 2.95 1.26 2.95  ;
        POLYGON 3.93 0.78 4.275 0.78 4.275 2.87 3.93 2.87  ;
        POLYGON 8.095 2.665 8.48 2.665 8.48 3.005 7.865 3.005 7.865 2.275 7.095 2.275 7.095 3.39 5.67 3.39 5.67 2.615 4.735 2.615 4.735 3.33 2.71 3.33 2.71 2.97 1.725 2.97 1.725 1.34 2.04 1.34 2.04 0.845 2.91 0.845 2.91 1.075 2.29 1.075 2.29 1.57 1.955 1.57 1.955 2.74 3.05 2.74 3.05 3.1 4.505 3.1 4.505 2.38 5.9 2.38 5.9 3.155 6.865 3.155 6.865 2.045 7.865 2.045 7.865 0.79 8.48 0.79 8.48 1.13 8.095 1.13  ;
        POLYGON 8.325 1.46 8.71 1.46 8.71 0.845 9.95 0.845 9.95 1.075 8.94 1.075 8.94 2.72 9.88 2.72 9.88 2.95 8.71 2.95 8.71 1.82 8.325 1.82  ;
        POLYGON 11.595 2.575 12.075 2.575 12.075 2.925 11.345 2.925 11.345 0.795 12.075 0.795 12.075 1.145 11.595 1.145  ;
        POLYGON 13.985 0.78 14.215 0.78 14.215 2.925 13.985 2.925  ;
        POLYGON 10.885 0.78 11.115 0.78 11.115 3.16 12.36 3.16 12.36 2.38 13.73 2.38 13.73 3.16 15.005 3.16 15.005 0.78 15.335 0.78 15.335 3.39 13.5 3.39 13.5 2.615 12.59 2.615 12.59 3.39 10.885 3.39  ;
        POLYGON 15.565 0.85 16.51 0.85 16.51 1.08 15.795 1.08 15.795 2.815 16.425 2.815 16.425 3.045 15.565 3.045  ;
        POLYGON 16.025 1.675 16.255 1.675 16.255 2.355 18.465 2.355 18.465 0.78 18.695 0.78 18.695 3.14 18.36 3.14 18.36 2.585 16.025 2.585  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux4_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__mux4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__mux4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN I0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5165 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.725 1.78 18.75 1.78 20.415 1.78 20.415 2.12 18.75 2.12 18.725 2.12  ;
    END
  END I0
  PIN I1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.5165 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.075 1.78 15.975 1.78 15.975 2.13 14.075 2.13  ;
    END
  END I1
  PIN I2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.025 1.01 1.025 1.01 2.835 0.705 2.835  ;
    END
  END I2
  PIN I3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.618 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.505 0.55 4.935 0.55 4.935 1.8 5.755 1.8 5.755 2.15 4.505 2.15  ;
    END
  END I3
  PIN S0
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.651 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.255 1.8 3.3 1.8 3.3 1.24 3.7 1.24 3.7 2.25 2.255 2.25  ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.033 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.41 1.305 11.775 1.305 11.775 1.77 12.19 1.77 12.775 1.77 12.775 3.32 12.405 3.32 12.405 2.15 12.19 2.15 11.41 2.15  ;
    END
  END S1
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.2064 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.23 0.6 6.6 0.6 6.6 1.8 8.425 1.8 8.425 0.6 8.84 0.6 8.84 2.925 8.425 2.925 8.425 2.15 6.615 2.15 6.615 2.925 6.23 2.925  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.575 0.475 2.575 0.475 3.62 1.65 3.62 5.12 3.62 5.12 2.845 5.46 2.845 5.46 3.62 7.35 3.62 7.35 2.845 7.69 2.845 7.69 3.62 9.53 3.62 9.53 2.845 9.87 2.845 9.87 3.62 10.72 3.62 12.19 3.62 15.145 3.62 15.145 2.845 15.49 2.845 15.49 3.62 17.575 3.62 19.43 3.62 19.43 2.815 19.77 2.815 19.77 3.62 20.935 3.62 21.28 3.62 21.28 4.22 20.935 4.22 17.575 4.22 12.19 4.22 10.72 4.22 1.65 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 19.815 0.3 19.815 1.145 19.585 1.145 19.585 0.3 15.335 0.3 15.335 1.145 15.105 1.145 15.105 0.3 9.875 0.3 9.875 1.16 9.645 1.16 9.645 0.3 7.635 0.3 7.635 1.16 7.405 1.16 7.405 0.3 5.395 0.3 5.395 1.16 5.165 1.16 5.165 0.3 0.475 0.3 0.475 1.13 0.245 1.13 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.26 0.845 1.65 0.845 1.65 1.075 1.495 1.075 1.495 2.95 1.26 2.95  ;
        POLYGON 3.93 0.78 4.275 0.78 4.275 2.87 3.93 2.87  ;
        POLYGON 10.335 2.38 10.72 2.38 10.72 3.005 10.49 3.005 10.49 2.615 9.3 2.615 9.3 3.39 7.92 3.39 7.92 2.615 7.12 2.615 7.12 3.39 5.755 3.39 5.755 2.615 4.735 2.615 4.735 3.33 2.71 3.33 2.71 2.97 1.725 2.97 1.725 1.34 2.04 1.34 2.04 0.845 2.91 0.845 2.91 1.075 2.29 1.075 2.29 1.57 1.955 1.57 1.955 2.74 3.05 2.74 3.05 3.1 4.505 3.1 4.505 2.38 5.985 2.38 5.985 3.16 6.89 3.16 6.89 2.38 8.15 2.38 8.15 3.155 9.07 3.155 9.07 2.38 10.105 2.38 10.105 0.79 10.72 0.79 10.72 1.13 10.335 1.13  ;
        POLYGON 10.565 1.46 10.95 1.46 10.95 0.845 12.19 0.845 12.19 1.075 11.18 1.075 11.18 2.72 12.12 2.72 12.12 2.95 10.95 2.95 10.95 1.82 10.565 1.82  ;
        POLYGON 13.835 2.575 14.315 2.575 14.315 2.925 13.585 2.925 13.585 0.795 14.315 0.795 14.315 1.145 13.835 1.145  ;
        POLYGON 16.225 0.78 16.455 0.78 16.455 2.925 16.225 2.925  ;
        POLYGON 13.125 0.78 13.355 0.78 13.355 3.16 14.6 3.16 14.6 2.38 15.97 2.38 15.97 3.16 17.245 3.16 17.245 0.78 17.575 0.78 17.575 3.39 15.74 3.39 15.74 2.615 14.83 2.615 14.83 3.39 13.125 3.39  ;
        POLYGON 17.805 0.85 18.75 0.85 18.75 1.08 18.035 1.08 18.035 2.815 18.665 2.815 18.665 3.045 17.805 3.045  ;
        POLYGON 18.265 1.675 18.495 1.675 18.495 2.355 20.705 2.355 20.705 0.78 20.935 0.78 20.935 3.14 20.6 3.14 20.6 2.585 18.265 2.585  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__mux4_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 2.8 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.24 0.555 1.605 0.555 1.605 1.44 2.055 1.44 2.055 1.82 1.24 1.82  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.635 1.06 1 1.06 1 2.19 0.635 2.19  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.9484 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.27 2.07 2.29 2.07 2.29 0.53 2.68 0.53 2.68 2.3 1.5 2.3 1.5 3.38 1.27 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.25 3.62 0.25 2.53 0.48 2.53 0.48 3.62 2.29 3.62 2.29 2.53 2.52 2.53 2.52 3.62 2.8 3.62 2.8 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 2.8 -0.3 2.8 0.3 0.48 0.3 0.48 0.805 0.25 0.805 0.25 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand2_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.04 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.114 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.24 3.16 1.24 3.16 1.56 0.62 1.56  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.114 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.8 4.03 1.8 4.03 2.12 0.62 2.12  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6016 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.22 2.36 4.26 2.36 4.26 1.535 3.46 1.535 3.46 1 2.15 1 2.15 0.68 3.82 0.68 3.82 1.265 4.49 1.265 4.49 2.68 3.535 2.68 3.535 3.38 3.305 3.38 3.305 2.68 1.58 2.68 1.58 3.38 1.22 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.64 0.475 2.64 0.475 3.62 2.285 3.62 2.285 3.085 2.515 3.085 2.515 3.62 4.325 3.62 4.325 3.085 4.555 3.085 4.555 3.62 5.04 3.62 5.04 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.04 -0.3 5.04 0.3 4.62 0.3 4.62 0.635 4.26 0.635 4.26 0.3 0.475 0.3 0.475 0.905 0.245 0.905 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand2_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.96 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.228 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.45 1.8 7.175 1.8 7.175 2.13 0.45 2.13  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.228 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.61 1.24 3.545 1.24 3.545 1.325 5.265 1.325 5.265 1.24 7.635 1.24 7.635 1.825 8.11 1.825 8.11 2.095 7.405 2.095 7.405 1.57 0.61 1.57  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.2401 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.36 8.34 2.36 8.34 1.575 7.885 1.575 7.885 1.01 5.035 1.01 5.035 1.095 3.775 1.095 3.775 1.01 2.14 1.01 2.14 0.68 4.005 0.68 4.005 0.865 4.805 0.865 4.805 0.68 8.115 0.68 8.115 1.345 8.57 1.345 8.57 2.68 7.615 2.68 7.615 3.39 7.385 3.39 7.385 2.68 5.575 2.68 5.575 3.39 5.345 3.39 5.345 2.68 3.535 2.68 3.535 3.39 3.305 3.39 3.305 2.68 1.495 2.68 1.495 3.39 1.265 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.64 0.475 2.64 0.475 3.62 2.285 3.62 2.285 2.93 2.515 2.93 2.515 3.62 4.325 3.62 4.325 2.93 4.555 2.93 4.555 3.62 6.365 3.62 6.365 2.93 6.595 2.93 6.595 3.62 8.405 3.62 8.405 2.93 8.635 2.93 8.635 3.62 8.96 3.62 8.96 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.96 -0.3 8.96 0.3 8.69 0.3 8.69 0.635 8.35 0.635 8.35 0.3 4.575 0.3 4.575 0.635 4.235 0.635 4.235 0.3 0.555 0.3 0.555 0.905 0.325 0.905 0.325 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand2_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 3.92 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9845 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.9 0.55 3.21 0.55 3.21 1.96 2.9 1.96  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9845 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 0.55 2.14 0.55 2.14 1.96 1.78 1.96  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9845 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.12 1.76 0.66 1.76 0.66 1.055 1.065 1.055 1.065 2.15 0.12 2.15  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.3064 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 2.36 3.44 2.36 3.44 0.655 3.67 0.655 3.67 3.38 3.38 3.38 3.38 2.78 1.63 2.78 1.63 3.38 1.4 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.38 3.62 0.38 2.53 0.61 2.53 0.61 3.62 2.365 3.62 2.365 3.13 2.705 3.13 2.705 3.62 3.92 3.62 3.92 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 3.92 -0.3 3.92 0.3 0.61 0.3 0.61 0.805 0.38 0.805 0.38 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand3_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.28 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.95 1.265 4.2 1.265 4.2 1.555 1.95 1.555  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.77 1.785 4.53 1.785 4.53 1.26 6.245 1.26 6.245 1.535 5.05 1.535 5.05 2.02 1.77 2.02  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.78 1.77 1.54 1.77 1.54 2.25 5.69 2.25 5.69 1.785 6.67 1.785 6.67 2.15 6.175 2.15 6.175 2.485 1.265 2.485 1.265 2.15 0.78 2.15  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.963 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.43 2.715 5.725 2.715 5.725 2.95 0.13 2.95 0.13 0.865 1.04 0.865 1.04 0.705 3.995 0.705 3.995 0.975 1.37 0.975 1.37 1.1 0.43 1.1  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.265 3.62 0.265 3.18 0.495 3.18 0.495 3.62 2.305 3.62 2.305 3.18 2.535 3.18 2.535 3.62 4.345 3.62 4.345 3.18 4.575 3.18 4.575 3.62 6.385 3.62 6.385 2.64 6.615 2.64 6.615 3.62 7.28 3.62 7.28 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.28 -0.3 7.28 0.3 6.615 0.3 6.615 0.9 6.385 0.9 6.385 0.3 0.69 0.3 0.69 0.635 0.35 0.635 0.35 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand3_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.05 1.79 12.67 1.79 12.67 2.13 9.05 2.13  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.65 1.79 8.53 1.79 8.53 2.15 0.65 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.71 1.33 3.45 1.33 3.45 1.21 5.66 1.21 5.66 1.33 7.54 1.33 7.54 1.56 1.71 1.56  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.8014 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 2.38 12.97 2.38 12.97 1.22 9.68 1.22 9.68 0.99 13.35 0.99 13.35 3.36 12.66 3.36 12.66 2.755 10.33 2.755 10.33 3.36 9.99 3.36 9.99 2.755 7.97 2.755 7.97 3.36 7.63 3.36 7.63 2.755 5.83 2.755 5.83 3.36 5.49 3.36 5.49 2.755 3.69 2.755 3.69 3.36 3.35 3.36 3.35 2.755 1.55 2.755 1.55 3.36 1.21 3.36  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.76 0.475 2.76 0.475 3.62 2.285 3.62 2.285 2.985 2.515 2.985 2.515 3.62 4.425 3.62 4.425 2.985 4.655 2.985 4.655 3.62 6.565 3.62 6.565 2.985 6.795 2.985 6.795 3.62 8.705 3.62 8.705 2.985 8.935 2.985 8.935 3.62 11.285 3.62 11.285 2.985 11.515 2.985 11.515 3.62 13.965 3.62 13.965 2.76 14.195 2.76 14.195 3.62 14.36 3.62 14.56 3.62 14.56 4.22 14.36 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 6.96 0.3 6.96 0.635 6.6 0.635 6.6 0.3 2.68 0.3 2.68 0.635 2.32 0.635 2.32 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.865 2.945 0.865 2.945 0.53 6.365 0.53 6.365 0.865 7.75 0.865 7.75 0.53 14.36 0.53 14.36 0.76 7.98 0.76 7.98 1.1 6.135 1.1 6.135 0.76 3.175 0.76 3.175 1.095 0.18 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nand3_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.04 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.02 1.21 4.37 1.21 4.37 2.19 4.02 2.19  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.9 0.61 3.24 0.61 3.24 2.19 2.9 2.19  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.61 2.14 0.61 2.14 2.19 1.8 2.19  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9145 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.21 1.02 1.21 1.02 1.89 1.4 1.89 1.4 2.19 0.66 2.19  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.2396 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.26 2.715 4.6 2.715 4.6 0.98 3.775 0.98 3.775 0.53 4.91 0.53 4.91 2.95 3.77 2.95 3.77 3.39 3.46 3.39 3.46 2.945 1.65 2.945 1.65 3.39 1.26 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.4 3.62 0.4 3.18 0.63 3.18 0.63 3.62 2.44 3.62 2.44 3.18 2.67 3.18 2.67 3.62 4.48 3.62 4.48 3.18 4.71 3.18 4.71 3.62 5.04 3.62 5.04 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.04 -0.3 5.04 0.3 0.63 0.3 0.63 0.98 0.4 0.98 0.4 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand4_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.96 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.829 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.61 1.82 2.35 1.82 2.35 1.445 4.03 1.445 4.03 1.675 2.58 1.675 2.58 2.1 0.61 2.1  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.829 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.81 1.905 4.455 1.905 4.455 1.75 5.5 1.75 5.5 1.465 6.15 1.465 6.15 1.695 5.775 1.695 5.775 2.135 2.81 2.135  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.829 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.61 1.21 1.755 1.21 1.755 0.985 4.13 0.985 4.13 0.99 7.19 0.99 7.19 1.555 6.81 1.555 6.81 1.22 4.08 1.22 4.08 1.215 2.095 1.215 2.095 1.59 0.61 1.59  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.829 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.69 2.34 1.845 2.34 1.845 2.365 6.38 2.365 6.38 1.825 8.19 1.825 8.19 2.26 6.66 2.26 6.66 2.595 0.69 2.595  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.4882 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.18 2.825 6.91 2.825 6.91 2.525 8.495 2.525 8.495 1.535 7.425 1.535 7.425 0.76 4.18 0.76 4.18 0.53 7.695 0.53 7.695 1.265 8.815 1.265 8.815 3.39 8.405 3.39 8.405 2.76 7.14 2.76 7.14 3.31 6.055 3.31 6.055 3.055 4.9 3.055 4.9 3.31 3.935 3.31 3.935 3.055 3.02 3.055 3.02 3.31 1.81 3.31 1.81 3.055 0.98 3.055 0.98 3.31 0.18 3.31  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.21 3.62 1.21 3.285 1.55 3.285 1.55 3.62 3.25 3.62 3.25 3.285 3.59 3.285 3.59 3.62 5.29 3.62 5.29 3.285 5.63 3.285 5.63 3.62 7.385 3.62 7.385 3 7.615 3 7.615 3.62 8.96 3.62 8.96 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.96 -0.3 8.96 0.3 8.635 0.3 8.635 0.83 8.405 0.83 8.405 0.3 0.475 0.3 0.475 0.83 0.245 0.83 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nand4_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nand4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nand4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.92 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.658 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.45 1.265 10.3 1.265 10.3 1.45 16.155 1.45 16.155 1.68 9.95 1.68 9.95 1.535 8.45 1.535  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.658 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.45 1.825 9.47 1.825 9.47 1.91 16.385 1.91 16.385 1.75 17.27 1.75 17.27 2.15 8.45 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.658 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.825 8.2 1.825 8.2 2.095 0.62 2.095  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.658 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.73 1.325 3.345 1.325 3.345 1.21 5.51 1.21 5.51 1.325 7.18 1.325 7.18 1.555 1.73 1.555  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.1796 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 2.38 17.505 2.38 17.505 1.22 10.6 1.22 10.6 0.99 17.73 0.99 17.775 0.99 17.775 2.655 17.73 2.655 16.655 2.655 16.655 3.31 16.425 3.31 16.425 2.655 14.175 2.655 14.175 3.31 13.945 3.31 13.945 2.655 12.135 2.655 12.135 3.31 11.905 3.31 11.905 2.655 9.655 2.655 9.655 3.31 9.425 3.31 9.425 2.655 7.615 2.655 7.615 3.31 7.385 3.31 7.385 2.655 5.575 2.655 5.575 3.31 5.345 3.31 5.345 2.655 3.535 2.655 3.535 3.31 3.305 3.31 3.305 2.655 1.495 2.655 1.495 3.31 1.265 3.31  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.84 0.475 2.84 0.475 3.62 2.285 3.62 2.285 2.935 2.515 2.935 2.515 3.62 4.325 3.62 4.325 2.935 4.555 2.935 4.555 3.62 6.365 3.62 6.365 2.935 6.595 2.935 6.595 3.62 8.405 3.62 8.405 2.935 8.635 2.935 8.635 3.62 10.885 3.62 10.885 2.935 11.115 2.935 11.115 3.62 12.925 3.62 12.925 2.935 13.155 2.935 13.155 3.62 15.405 3.62 15.405 2.935 15.635 2.935 15.635 3.62 17.445 3.62 17.445 2.935 17.675 2.935 17.675 3.62 17.73 3.62 17.92 3.62 17.92 4.22 17.73 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.92 -0.3 17.92 0.3 6.66 0.3 6.66 0.635 6.3 0.635 6.3 0.3 2.58 0.3 2.58 0.635 2.22 0.635 2.22 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.865 2.81 0.865 2.81 0.69 6.07 0.69 6.07 0.865 7.405 0.865 7.405 0.53 17.73 0.53 17.73 0.76 7.635 0.76 7.635 1.095 5.84 1.095 5.84 0.98 3.04 0.98 3.04 1.095 0.18 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nand4_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 3.36 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.949 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.6 2.13 0.6 2.13 1.79 2.855 1.79 2.855 2.13 1.825 2.13  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.949 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.18 1.01 1.18 1.01 3.32 0.705 3.32  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8306 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.24 0.6 1.595 0.6 1.595 2.36 2.665 2.36 2.665 3.38 2.385 3.38 2.385 2.68 1.24 2.68  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 3.36 3.62 3.36 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 3.36 -0.3 3.36 0.3 2.715 0.3 2.715 1.09 2.485 1.09 2.485 0.3 0.475 0.3 0.475 0.945 0.245 0.945 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor2_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.48 1.77 3.22 1.77 3.22 2.15 1.48 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.898 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.81 1.58 1.06 1.58 1.06 2.38 3.48 2.38 3.48 1.77 4.39 1.77 4.39 2.15 3.78 2.15 3.78 2.7 0.81 2.7  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.283 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.39 3.14 4.095 3.14 4.095 2.8 4.625 2.8 4.625 1.32 1.365 1.32 1.365 0.53 1.595 0.53 1.595 1.05 3.605 1.05 3.605 0.53 3.835 0.53 3.835 1.05 4.895 1.05 4.895 3.035 4.325 3.035 4.325 3.37 2.39 3.37  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.295 3.62 0.295 2.625 0.525 2.625 0.525 3.62 4.61 3.62 4.61 3.285 4.97 3.285 4.97 3.62 5.6 3.62 5.6 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 5.02 0.3 5.02 0.82 4.66 0.82 4.66 0.3 2.78 0.3 2.78 0.82 2.42 0.82 2.42 0.3 0.54 0.3 0.54 0.82 0.18 0.82 0.18 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor2_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.796 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.65 1.8 8.415 1.8 8.415 2.12 1.65 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.796 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.795 1.325 8.04 1.325 8.04 1.22 9.42 1.22 9.42 2.255 9.06 2.255 9.06 1.56 0.795 1.56  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.932 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.13 0.865 1.365 0.865 1.365 0.53 1.595 0.53 1.595 0.865 3.605 0.865 3.605 0.53 3.835 0.53 3.835 0.865 5.845 0.865 5.845 0.53 6.075 0.53 6.075 0.865 7.5 0.865 7.5 0.53 8.41 0.53 8.41 0.76 7.73 0.76 7.73 1.095 0.43 1.095 0.43 2.35 7.195 2.35 7.195 3.38 6.965 3.38 6.965 2.7 5.65 2.7 5.65 2.585 3.87 2.585 3.87 2.7 2.715 2.7 2.715 3.38 2.485 3.38 2.485 2.7 1.17 2.7 1.17 2.585 0.13 2.585  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.24 3.62 0.24 2.815 0.58 2.815 0.58 3.62 4.67 3.62 4.67 2.815 5.01 2.815 5.01 3.62 9.1 3.62 9.1 2.815 9.44 2.815 9.44 3.62 10.08 3.62 10.08 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.5 0.3 9.5 0.635 9.14 0.635 9.14 0.3 7.25 0.3 7.25 0.635 6.91 0.635 6.91 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.54 0.3 0.54 0.635 0.18 0.635 0.18 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor2_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.91 1.575 3.25 1.575 3.25 3.39 2.91 3.39  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.79 1.575 2.13 1.575 2.13 3.39 1.79 3.39  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.49 1.76 1.56 1.76 1.56 3.39 1.22 3.39 1.22 2.19 0.49 2.19  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.9832 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.31 0.695 1.65 0.695 1.65 1.05 3.55 1.05 3.55 0.695 3.89 0.695 3.89 3.39 3.49 3.39 3.49 1.285 1.31 1.285  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.575 2.53 0.575 3.62 4.48 3.62 4.48 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 2.77 0.3 2.77 0.82 2.43 0.82 2.43 0.3 0.53 0.3 0.53 0.82 0.19 0.82 0.19 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor3_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.84 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.955 1.825 4.39 1.825 4.39 2.095 2.955 2.095  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.935 1.77 2.385 1.77 2.385 1.36 4.895 1.36 4.895 1.77 5.65 1.77 5.65 2.15 4.625 2.15 4.625 1.59 2.71 1.59 2.71 2.095 1.935 2.095  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.39 1.58 1.39 1.58 2.38 6.25 2.38 6.25 1.73 6.63 1.73 6.63 2.655 1.305 2.655 1.305 1.665 0.705 1.665  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.6492 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.145 0.53 0.53 0.53 0.53 0.885 1.89 0.885 1.89 0.53 3.31 0.53 3.31 0.885 4.13 0.885 4.13 0.53 5.55 0.53 5.55 0.885 6.905 0.885 6.905 0.53 7.25 0.53 7.25 1.115 0.42 1.115 0.42 2.02 1.055 2.02 1.055 2.94 3.84 2.94 3.84 3.235 0.825 3.235 0.825 2.25 0.145 2.25  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.59 0.575 2.59 0.575 3.62 6.865 3.62 6.865 2.63 7.095 2.63 7.095 3.62 7.84 3.62 7.84 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.84 -0.3 7.84 0.3 6.14 0.3 6.14 0.655 5.78 0.655 5.78 0.3 3.9 0.3 3.9 0.655 3.54 0.655 3.54 0.3 1.66 0.3 1.66 0.655 1.3 0.655 1.3 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor3_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.55 1.41 12.18 1.41 12.18 1.64 9.96 1.64 9.96 2.85 9.55 2.85  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.405 1.75 1.57 1.75 1.57 1.87 7.97 1.87 7.97 1.75 9.03 1.75 9.03 2.15 0.405 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.556 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.79 1.41 3.47 1.41 3.47 1.01 3.91 1.01 3.91 1.41 5.7 1.41 5.7 1.01 6.15 1.01 6.15 1.41 7.735 1.41 7.735 1.64 1.79 1.64  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.9636 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.19 1.875 12.42 1.875 12.42 1.18 6.45 1.18 6.45 0.76 5.47 0.76 5.47 1.18 4.21 1.18 4.21 0.76 3.23 0.76 3.23 1.18 1.255 1.18 1.255 0.53 1.65 0.53 1.65 0.945 3 0.945 3 0.53 4.44 0.53 4.44 0.945 5.24 0.945 5.24 0.53 6.68 0.53 6.68 0.945 7.95 0.945 7.95 0.53 8.82 0.53 8.82 0.945 9.72 0.945 9.72 0.53 11.16 0.53 11.16 0.945 12.46 0.945 12.46 0.53 12.85 0.53 12.85 2.91 12.46 2.91 12.46 2.11 10.555 2.11 10.555 2.91 10.19 2.91  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.385 3.62 2.385 3.155 2.615 3.155 2.615 3.62 6.865 3.62 6.865 3.155 7.095 3.155 7.095 3.62 13.815 3.62 14.56 3.62 14.56 4.22 13.815 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 13.97 0.3 13.97 0.655 13.63 0.655 13.63 0.3 11.73 0.3 11.73 0.655 11.39 0.655 11.39 0.3 9.49 0.3 9.49 0.655 9.15 0.655 9.15 0.3 7.25 0.3 7.25 0.655 6.91 0.655 6.91 0.3 5.01 0.3 5.01 0.655 4.67 0.655 4.67 0.3 2.77 0.3 2.77 0.655 2.43 0.655 2.43 0.3 0.53 0.3 0.53 0.655 0.19 0.655 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 2.57 8.22 2.57 8.22 3.16 11.345 3.16 11.345 2.53 11.575 2.53 11.575 3.16 13.585 3.16 13.585 2.53 13.815 2.53 13.815 3.39 7.99 3.39 7.99 2.8 4.855 2.8 4.855 3.38 4.625 3.38 4.625 2.8 0.475 2.8 0.475 3.38 0.245 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nor3_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.826 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.03 1.685 4.37 1.685 4.37 3.38 4.03 3.38  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.826 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.91 1.685 3.25 1.685 3.25 3.38 2.91 3.38  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.826 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.79 1.685 2.13 1.685 2.13 3.38 1.79 3.38  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.826 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.585 1.685 1.56 1.685 1.56 3.38 1.22 3.38 1.22 2.195 0.585 2.195  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.9112 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.255 0.53 1.65 0.53 1.65 1.07 3.505 1.07 3.505 0.53 3.89 0.53 3.89 1.07 4.91 1.07 4.91 2.38 4.905 2.38 4.905 3.38 4.61 3.38 4.61 1.305 1.255 1.305  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.575 2.53 0.575 3.62 5.6 3.62 5.6 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 4.955 0.3 4.955 0.84 4.725 0.84 4.725 0.3 2.715 0.3 2.715 0.84 2.485 0.84 2.485 0.3 0.475 0.3 0.475 0.84 0.245 0.84 0.245 0.3 0 0.3  ;
    END
  END VSS
END gf180mcu_fd_sc_mcu7t5v0__nor4_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.835 1.465 8.47 1.465 8.47 1.24 9.63 1.24 9.63 1.56 8.745 1.56 8.745 1.695 6.835 1.695  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.69 1.75 6.605 1.75 6.605 1.93 8.975 1.93 8.975 1.8 9.63 1.8 9.63 2.16 5.69 2.16  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 1.825 1.275 1.825 1.275 1.93 3.45 1.93 3.45 1.825 4.615 1.825 4.615 2.16 0.385 2.16  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.652 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 1.265 1.735 1.265 1.735 1.465 3.22 1.465 3.22 1.695 1.505 1.695 1.505 1.565 0.385 1.565  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.631 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.17 0.53 2.205 0.53 2.205 1.005 3.005 1.005 3.005 0.53 4.625 0.53 4.625 1.005 5.425 1.005 5.425 0.53 7.045 0.53 7.045 1.005 7.845 1.005 7.845 0.53 8.95 0.53 8.95 0.975 8.145 0.975 8.145 1.235 6.815 1.235 6.815 0.975 5.655 0.975 5.655 1.235 5.46 1.235 5.46 2.39 7.79 2.39 7.79 2.665 5.13 2.665 5.13 1.235 4.395 1.235 4.395 0.975 3.235 0.975 3.235 1.235 1.975 1.235 1.975 0.975 1.17 0.975  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.44 3.62 2.44 2.935 2.67 2.935 2.67 3.62 9.7 3.62 10.08 3.62 10.08 4.22 9.7 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.855 0.3 9.855 0.775 9.515 0.775 9.515 0.3 7.615 0.3 7.615 0.775 7.275 0.775 7.275 0.3 5.195 0.3 5.195 0.775 4.855 0.775 4.855 0.3 2.775 0.3 2.775 0.775 2.435 0.775 2.435 0.3 0.535 0.3 0.535 0.775 0.195 0.775 0.195 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.35 2.39 4.615 2.39 4.615 2.965 9.47 2.965 9.47 2.53 9.7 2.53 9.7 3.38 9.47 3.38 9.47 3.195 4.385 3.195 4.385 2.625 0.58 2.625 0.58 3.38 0.35 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nor4_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__nor4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__nor4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 20.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.294 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.855 1.45 13.545 1.45 13.545 1.17 13.89 1.17 13.89 1.45 16.325 1.45 16.325 1.17 16.685 1.17 16.685 1.45 18.66 1.45 18.66 1.265 20.11 1.265 20.11 1.535 18.89 1.535 18.89 1.68 11.855 1.68  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.294 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.51 1.77 11.625 1.77 11.625 1.91 19.14 1.91 19.14 1.77 20.11 1.77 20.11 2.15 10.51 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.294 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.61 1.82 1.295 1.82 1.295 1.91 8.46 1.91 8.46 1.73 9.395 1.73 9.395 2.15 0.61 2.15  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.294 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.61 1.265 1.76 1.265 1.76 1.45 3.51 1.45 3.51 1.17 3.85 1.17 3.85 1.45 6.24 1.45 6.24 1.17 6.585 1.17 6.585 1.45 8.21 1.45 8.21 1.68 1.54 1.68 1.54 1.535 0.61 1.535  ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.8304 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.17 0.53 2.25 0.53 2.25 0.99 3.05 0.99 3.05 0.53 4.67 0.53 4.67 0.99 5.47 0.99 5.47 0.53 7.09 0.53 7.09 0.99 7.89 0.99 7.89 0.53 9.51 0.53 9.51 0.99 10.405 0.99 10.405 0.53 12.21 0.53 12.21 0.99 13.01 0.99 13.01 0.53 14.8 0.53 14.8 0.99 15.6 0.99 15.6 0.53 17.39 0.53 17.39 0.99 18.2 0.99 18.2 0.53 19.55 0.53 19.55 0.975 18.43 0.975 18.43 1.22 17.16 1.22 17.16 0.92 15.83 0.92 15.83 1.22 14.57 1.22 14.57 0.92 13.24 0.92 13.24 1.22 11.07 1.22 11.07 1.52 10.24 1.52 10.24 2.38 18.07 2.38 18.07 2.835 17.215 2.835 17.215 2.655 12.91 2.655 12.91 2.84 12.57 2.84 12.57 2.665 9.66 2.665 9.66 1.48 8.535 1.48 8.535 0.975 8.12 0.975 8.12 1.22 6.86 1.22 6.86 0.92 5.7 0.92 5.7 1.22 4.44 1.22 4.44 0.92 3.28 0.92 3.28 1.22 2.02 1.22 2.02 0.975 1.17 0.975  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.485 3.62 2.485 2.95 2.715 2.95 2.715 3.62 7.325 3.62 7.325 2.95 7.555 2.95 7.555 3.62 20.38 3.62 20.72 3.62 20.72 4.22 20.38 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 20.72 -0.3 20.72 0.3 20.48 0.3 20.48 0.76 20.14 0.76 20.14 0.3 17.97 0.3 17.97 0.76 17.63 0.76 17.63 0.3 15.37 0.3 15.37 0.76 15.03 0.76 15.03 0.3 12.78 0.3 12.78 0.76 12.44 0.76 12.44 0.3 10.175 0.3 10.175 0.76 9.835 0.76 9.835 0.3 7.66 0.3 7.66 0.76 7.32 0.76 7.32 0.3 5.24 0.3 5.24 0.76 4.9 0.76 4.9 0.3 2.82 0.3 2.82 0.76 2.48 0.76 2.48 0.3 0.58 0.3 0.58 0.76 0.24 0.76 0.24 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.395 2.415 8.74 2.415 8.74 3.15 14.89 3.15 14.89 2.945 15.23 2.945 15.23 3.15 20.04 3.15 20.04 2.53 20.38 2.53 20.38 3.385 8.51 3.385 8.51 2.65 5.135 2.65 5.135 3.39 4.905 3.39 4.905 2.65 0.625 2.65 0.625 3.38 0.395 3.38  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__nor4_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai21_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai21_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.55 2.16 0.55 2.16 2.32 1.825 2.32  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.55 1 0.55 1 2.23 0.705 2.23  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 0.55 3.28 0.55 3.28 1.6 4.35 1.6 4.35 2.15 3.375 2.15 3.375 1.9 2.945 1.9  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.276 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.23 0.55 1.595 0.55 1.595 2.59 2.615 2.59 2.615 2.93 1.23 2.93  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.295 3.62 0.295 2.92 0.525 2.92 0.525 3.62 3.075 3.62 3.605 3.62 3.605 2.92 3.835 2.92 3.835 3.62 4.48 3.62 4.48 4.22 3.075 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 3.835 0.3 3.835 0.93 3.605 0.93 3.605 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.55 0.475 0.55 0.475 1.16 0.475 2.46 0.985 2.46 0.985 3.16 2.845 3.16 2.845 2.36 2.485 2.36 2.485 0.55 2.715 0.55 2.715 2.13 3.075 2.13 3.075 3.39 0.755 3.39 0.755 2.69 0.245 2.69 0.245 1.16  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai21_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai21_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai21_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.4 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.97 1.79 6.08 1.79 6.08 2.12 3.97 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.98 1.83 3.655 1.83 3.655 2.35 6.355 2.35 6.355 1.79 7.25 1.79 7.25 2.195 6.615 2.195 6.615 2.68 3.395 2.68 3.395 2.09 2.98 2.09  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.939 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.785 2.75 1.785 2.75 2.12 0.28 2.12  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3096 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.45 3.095 2.45 3.095 3.05 6.845 3.05 6.845 2.445 7.5 2.445 7.5 1.56 3.77 1.56 3.77 0.99 4.11 0.99 4.11 1.22 6.01 1.22 6.01 0.99 6.35 0.99 6.35 1.22 7.7 1.22 7.73 1.22 7.73 2.675 7.7 2.675 7.075 2.675 7.075 3.28 2.865 3.28 2.865 2.68 1.595 2.68 1.595 3.335 1.365 3.335  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.995 0.575 2.995 0.575 3.62 2.385 3.62 2.385 2.995 2.615 2.995 2.615 3.62 7.305 3.62 7.305 2.995 7.535 2.995 7.535 3.62 7.7 3.62 8.4 3.62 8.4 4.22 7.7 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.4 -0.3 8.4 0.3 1.595 0.3 1.595 1.015 1.365 1.015 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.635 0.475 0.635 0.475 1.31 2.485 1.31 2.485 0.53 7.7 0.53 7.7 0.76 2.715 0.76 2.715 1.545 0.245 1.545  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai21_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai21_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai21_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.12 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.53 1.8 3.35 1.8 3.35 1.45 8.07 1.45 8.07 1.68 3.58 1.68 3.58 2.12 1.53 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.68 1.695 1 1.695 1 2.36 3.87 2.36 3.87 1.91 9.14 1.91 9.14 2.14 4.1 2.14 4.1 2.68 0.68 2.68  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.878 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.02 1.8 14.355 1.8 14.55 1.8 14.55 2.12 14.355 2.12 10.02 2.12  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.0305 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.085 2.92 4.41 2.92 4.41 2.825 5.71 2.825 5.71 2.92 9.385 2.92 9.385 1.22 1.52 1.22 1.52 0.99 9.615 0.99 9.615 2.36 13.135 2.36 13.135 3.25 12.905 3.25 12.905 2.68 11.095 2.68 11.095 3.25 10.865 3.25 10.865 2.68 9.615 2.68 9.615 3.24 5.48 3.24 5.48 3.055 4.64 3.055 4.64 3.24 1.085 3.24  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.91 0.475 2.91 0.475 3.62 4.89 3.62 4.89 3.285 5.23 3.285 5.23 3.62 9.845 3.62 9.845 2.91 10.075 2.91 10.075 3.62 11.885 3.62 11.885 2.91 12.115 2.91 12.115 3.62 13.925 3.62 13.925 2.91 14.155 2.91 14.155 3.62 14.355 3.62 15.12 3.62 15.12 4.22 14.355 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 15.12 -0.3 15.12 0.3 13.235 0.3 13.235 0.91 13.005 0.91 13.005 0.3 10.995 0.3 10.995 0.91 10.765 0.91 10.765 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.53 10.38 0.53 10.38 1.16 11.885 1.16 11.885 0.57 12.115 0.57 12.115 1.16 14.125 1.16 14.125 0.57 14.355 0.57 14.355 1.39 10.15 1.39 10.15 0.76 0.18 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai21_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai211_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai211_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.55 2.12 0.55 2.12 2.135 1.825 2.135  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.55 1 0.55 1 2.23 0.705 2.23  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9845 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.36 1.16 2.66 1.16 2.66 1.8 3.37 1.8 3.37 2.12 2.36 2.12  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9845 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.24 3.94 1.24 3.94 1.8 4.97 1.8 4.97 2.12 3.65 2.12 3.65 1.56 2.89 1.56  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.67285 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.24 0.55 1.595 0.55 1.595 2.365 4.92 2.365 4.92 2.93 4.58 2.93 4.58 2.595 2.77 2.595 2.77 2.93 2.43 2.93 2.43 2.7 1.24 2.7  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.295 3.62 0.295 2.92 0.525 2.92 0.525 3.62 3.55 3.62 3.55 3.285 3.89 3.285 3.89 3.62 5.45 3.62 5.6 3.62 5.6 4.22 5.45 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 4.955 0.3 4.955 0.89 4.725 0.89 4.725 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.55 0.475 0.55 0.475 2.46 0.985 2.46 0.985 3.16 3.06 3.16 3.06 2.825 4.35 2.825 4.35 3.16 5.22 3.16 5.22 1.37 4.24 1.37 4.24 0.835 2.43 0.835 2.43 0.605 4.24 0.605 4.24 0.6 4.47 0.6 4.47 1.14 5.45 1.14 5.45 3.39 4.12 3.39 4.12 3.055 3.29 3.055 3.29 3.39 0.755 3.39 0.755 2.69 0.245 2.69  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai211_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai211_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai211_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.56 1.79 3.87 1.79 3.87 2.12 1.56 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.16 1.145 1.16 1.145 2.35 4.12 2.35 4.12 1.79 4.9 1.79 4.9 2.12 4.38 2.12 4.38 2.68 0.825 2.68  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.72 1.19 6.485 1.19 6.485 1.325 8.38 1.325 8.38 1.19 9.42 1.19 9.42 2.19 8.865 2.19 8.865 1.555 6.04 1.555 6.04 2.15 5.72 2.15  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.28 1.8 8.32 1.8 8.32 2.14 6.28 2.14  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.8374 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.13 2.92 4.63 2.92 4.63 2.37 5.15 2.37 5.15 1.56 1.53 1.56 1.53 0.99 1.87 0.99 1.87 1.22 3.77 1.22 3.77 0.99 4.11 0.99 4.11 1.22 5.48 1.22 5.48 2.38 8.56 2.38 8.56 3.275 8.33 3.275 8.33 2.68 6.52 2.68 6.52 3.275 6.29 3.275 6.29 2.68 4.86 2.68 4.86 3.28 2.13 3.28  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.485 0.575 2.485 0.575 3.62 5.115 3.62 5.115 3.205 5.455 3.205 5.455 3.62 7.255 3.62 7.255 3.205 7.595 3.205 7.595 3.62 9.35 3.62 9.35 2.595 9.58 2.595 9.58 3.62 9.645 3.62 10.08 3.62 10.08 4.22 9.645 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 7.595 0.3 7.595 0.635 7.255 0.635 7.255 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.53 6.965 0.53 6.965 0.865 7.85 0.865 7.85 0.53 9.645 0.53 9.645 0.76 8.08 0.76 8.08 1.095 6.735 1.095 6.735 0.76 0.18 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai211_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai211_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai211_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 18.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.96 1.45 6.79 1.45 6.79 1.77 8.31 1.77 8.31 2.12 6.54 2.12 6.54 1.68 1.96 1.68  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.91 6.205 1.91 6.205 2.36 8.54 2.36 8.54 1.77 9.41 1.77 9.41 2.12 8.88 2.12 8.88 2.68 5.955 2.68 5.955 2.14 0.62 2.14  ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.2 1.325 12.93 1.325 12.93 1.22 15.08 1.22 15.08 1.325 17.76 1.325 17.76 1.555 10.52 1.555 10.52 2.425 10.2 2.425  ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.938 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.75 1.8 16.84 1.8 16.84 2.12 10.75 2.12  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.279 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.65 2.475 2.99 2.475 2.99 2.92 4.39 2.92 4.39 2.795 5.725 2.795 5.725 2.92 9.09 2.92 9.09 2.795 9.64 2.795 9.64 1.22 1.52 1.22 1.52 0.99 9.96 0.99 9.96 2.795 17.45 2.795 17.45 3.24 16.4 3.24 16.4 3.055 15.56 3.055 15.56 3.24 14.36 3.24 14.36 3.055 13.52 3.055 13.52 3.24 12.32 3.24 12.32 3.055 11.48 3.055 11.48 3.24 10.175 3.24 10.175 3.025 9.34 3.025 9.34 3.24 5.475 3.24 5.475 3.025 4.64 3.025 4.64 3.24 2.99 3.24 2.99 3.325 2.65 3.325  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.575 2.53 0.575 3.62 4.89 3.62 4.89 3.285 5.23 3.285 5.23 3.62 9.59 3.62 9.59 3.285 9.93 3.285 9.93 3.62 11.73 3.62 11.73 3.285 12.07 3.285 12.07 3.62 13.77 3.62 13.77 3.285 14.11 3.285 14.11 3.62 15.81 3.62 15.81 3.285 16.15 3.285 16.15 3.62 17.905 3.62 17.905 2.595 18.135 2.595 18.135 3.62 18.2 3.62 18.48 3.62 18.48 4.22 18.2 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 18.48 -0.3 18.48 0.3 16.15 0.3 16.15 0.635 15.81 0.635 15.81 0.3 12.07 0.3 12.07 0.635 11.73 0.635 11.73 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.53 10.885 0.53 10.885 0.865 12.32 0.865 12.32 0.53 15.56 0.53 15.56 0.865 18.2 0.865 18.2 1.095 15.33 1.095 15.33 0.76 12.55 0.76 12.55 1.095 10.655 1.095 10.655 0.76 0.18 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai211_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai22_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai22_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.945 0.55 3.24 0.55 3.24 2.22 2.945 2.22  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.065 0.55 4.38 0.55 4.38 2.22 4.065 2.22  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.685 2.715 1.685 2.715 2.19 2.16 2.19 2.16 2.845 1.8 2.845  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.61 1.03 1.61 1.03 3.32 0.705 3.32  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.44 2.68 3.48 2.68 3.48 0.55 3.835 0.55 3.835 2.91 2.44 2.91  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.59 0.475 2.59 0.475 3.62 4.625 3.62 4.625 2.96 4.855 2.96 4.855 3.62 4.955 3.62 5.6 3.62 5.6 4.22 4.955 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.55 3.14 4.135 3.14 4.135 2.45 4.725 2.45 4.725 0.55 4.955 0.55 4.955 2.68 4.365 2.68 4.365 3.37 1.32 3.37 1.32 1.095 0.245 1.095 0.245 0.55 0.475 0.55 0.475 0.865 2.485 0.865 2.485 0.55 2.715 0.55 2.715 1.095 1.55 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai22_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai22_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai22_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.64 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.25 1.8 8.715 1.8 8.715 2.12 6.25 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.27 1.8 6.02 1.8 6.02 2.36 8.955 2.36 8.955 1.585 9.295 1.585 9.295 2.68 5.69 2.68 5.69 2.12 5.27 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.475 1.785 3.27 1.785 3.27 2.12 1.475 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.585 1.165 1.585 1.165 2.36 3.5 2.36 3.5 1.77 4.48 1.77 4.48 2.125 3.82 2.125 3.82 2.68 0.825 2.68  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3774 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.175 2.92 4.11 2.92 4.11 2.36 4.755 2.36 4.755 1.24 6.01 1.24 6.01 0.99 6.35 0.99 6.35 1.24 8.25 1.24 8.25 0.99 8.59 0.99 8.59 1.56 5.015 1.56 5.015 2.36 5.445 2.36 5.445 2.92 7.865 2.92 7.865 3.24 5.195 3.24 5.195 2.68 4.385 2.68 4.385 3.24 2.175 3.24  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.59 0.575 2.59 0.575 3.62 4.725 3.62 4.725 2.975 4.955 2.975 4.955 3.62 9.545 3.62 9.545 2.59 9.775 2.59 9.775 3.62 9.94 3.62 10.64 3.62 10.64 4.22 9.94 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.64 -0.3 10.64 0.3 3.835 0.3 3.835 0.815 3.605 0.815 3.605 0.3 1.595 0.3 1.595 0.815 1.365 0.815 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.53 0.53 0.53 0.53 1.045 2.43 1.045 2.43 0.53 2.77 0.53 2.77 1.045 4.225 1.045 4.225 0.53 9.94 0.53 9.94 0.76 4.455 0.76 4.455 1.275 0.19 1.275  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai22_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai22_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai22_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.73 1.785 12.29 1.785 12.29 1.45 17.12 1.45 17.12 1.68 12.54 1.68 12.54 2.12 10.73 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.61 1.8 10.5 1.8 10.5 2.36 12.875 2.36 12.875 1.91 18.46 1.91 18.46 2.14 13.125 2.14 13.125 2.68 10.2 2.68 10.2 2.12 9.61 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.53 1.785 3.11 1.785 3.11 1.405 7.94 1.405 7.94 1.635 3.36 1.635 3.36 2.12 1.53 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.585 1.145 1.585 1.145 2.36 3.69 2.36 3.69 1.865 8.85 1.865 8.85 2.095 3.94 2.095 3.94 2.68 0.825 2.68  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.369 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.73 2.92 4.17 2.92 4.17 2.795 6.91 2.795 6.91 2.57 7.25 2.57 7.25 2.795 9.08 2.795 9.08 0.99 17.56 0.99 17.56 1.22 9.38 1.22 9.38 2.795 9.99 2.795 9.99 2.92 13.355 2.92 13.355 2.795 14.69 2.795 14.69 2.92 16.145 2.92 16.145 2.485 16.375 2.485 16.375 3.38 14.44 3.38 14.44 3.025 13.605 3.025 13.605 3.24 9.74 3.24 9.74 3.025 8.905 3.025 8.905 3.38 5.255 3.38 5.255 3.025 4.42 3.025 4.42 3.24 1.73 3.24  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.59 0.575 2.59 0.575 3.62 4.67 3.62 4.67 3.255 5.01 3.255 5.01 3.62 9.15 3.62 9.15 3.255 9.49 3.255 9.49 3.62 13.85 3.62 13.85 3.255 14.19 3.255 14.19 3.62 18.505 3.62 18.505 2.59 18.735 2.59 18.735 3.62 18.9 3.62 19.6 3.62 19.6 4.22 18.9 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.6 -0.3 19.6 0.3 8.37 0.3 8.37 0.715 8.03 0.715 8.03 0.3 6.13 0.3 6.13 0.715 5.79 0.715 5.79 0.3 3.89 0.3 3.89 0.715 3.55 0.715 3.55 0.3 1.65 0.3 1.65 0.715 1.31 0.715 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.19 0.55 0.53 0.55 0.53 0.945 2.43 0.945 2.43 0.55 2.77 0.55 2.77 0.945 4.67 0.945 4.67 0.55 5.01 0.55 5.01 0.945 6.91 0.945 6.91 0.55 7.25 0.55 7.25 0.945 8.61 0.945 8.61 0.53 18.9 0.53 18.9 0.76 8.84 0.76 8.84 1.175 0.19 1.175  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai22_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai221_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai221_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.16 1.17 5.5 1.17 5.5 1.77 6.11 1.77 6.11 2.15 5.16 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.01 1.17 4.39 1.17 4.39 2.135 4.01 2.135  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.24 1.345 2.11 1.345 2.11 1.575 1.56 1.575 1.56 3.32 1.24 3.32  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.345 1 1.345 1 3.32 0.705 3.32  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9645 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.34 1.21 2.715 1.21 2.945 1.21 2.945 0.61 3.26 0.61 3.26 1.665 2.715 1.665 2.34 1.665  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7536 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.91 2.38 6.11 2.38 6.11 2.93 5.77 2.93 5.77 2.7 4.795 2.7 4.795 2.595 2.77 2.595 2.77 2.93 2.43 2.93 2.43 2.365 4.62 2.365 4.62 0.61 5.095 0.61 5.095 0.91 4.91 0.91  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 3.61 3.62 3.61 3.285 3.95 3.285 3.95 3.62 6.57 3.62 6.72 3.62 6.72 4.22 6.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.72 -0.3 6.72 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.625 0.475 0.625 0.475 0.865 1.88 0.865 1.88 0.625 2.715 0.625 2.715 0.965 2.11 0.965 2.11 1.095 0.245 1.095  ;
        POLYGON 2.18 3.16 3.13 3.16 3.13 2.825 4.52 2.825 4.52 3.16 6.34 3.16 6.34 0.91 5.87 0.91 5.87 0.68 6.57 0.68 6.57 3.39 4.29 3.39 4.29 3.055 3.36 3.055 3.36 3.39 1.95 3.39 1.95 1.905 3.54 1.905 3.54 0.68 3.95 0.68 3.95 0.91 3.77 0.91 3.77 2.135 2.18 2.135  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai221_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai221_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai221_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.88 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.16 1.77 8.82 1.77 8.82 2.365 11.34 2.365 11.34 1.77 12.59 1.77 12.59 2.15 11.57 2.15 11.57 2.595 8.55 2.595 8.55 2.15 8.16 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.05 1.8 11.11 1.8 11.11 2.12 9.05 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.53 1.8 4.71 1.8 4.71 2.12 1.53 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.625 1.16 1.69 1.16 1.69 1.34 4.455 1.34 4.455 1.57 1 1.57 1 2.275 0.625 2.275  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.969 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.105 1.8 6.865 1.8 7.33 1.8 7.33 2.12 6.865 2.12 5.105 2.12  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 3.382 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.915 2.825 12.58 2.825 12.58 3.26 10.525 3.26 10.525 3.055 9.54 3.055 9.54 3.26 7.56 3.26 7.56 2.68 6.865 2.68 5.775 2.68 5.775 3.11 5.545 3.11 5.545 2.68 2.715 2.68 2.715 3.375 2.485 3.375 2.485 2.36 6.865 2.36 7.56 2.36 7.56 0.99 11.33 0.99 11.33 1.22 7.915 1.22  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.69 0.475 2.69 0.475 3.62 4.67 3.62 4.67 3.09 5.01 3.09 5.01 3.62 6.51 3.62 6.51 3.09 6.85 3.09 6.85 3.62 6.865 3.62 9.87 3.62 9.87 3.285 10.21 3.285 10.21 3.62 12.68 3.62 12.88 3.62 12.88 4.22 12.68 4.22 6.865 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.88 -0.3 12.88 0.3 5.01 0.3 5.01 0.635 4.665 0.635 4.665 0.3 2.77 0.3 2.77 0.635 2.425 0.635 2.425 0.3 0.53 0.3 0.53 0.635 0.185 0.635 0.185 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.26 0.55 2.17 0.55 2.17 0.865 5.11 0.865 5.11 0.99 6.865 0.99 6.865 1.22 4.86 1.22 4.86 1.095 1.94 1.095 1.94 0.78 1.26 0.78  ;
        POLYGON 5.38 0.53 12.68 0.53 12.68 0.76 5.38 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai221_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai221_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai221_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 24.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.015 1.6 15.245 1.6 15.245 2.365 18.32 2.365 18.32 1.91 18.66 1.91 18.66 2.365 19.34 2.365 19.34 1.91 22.385 1.91 22.385 1.79 23.06 1.79 23.06 1.12 23.42 1.12 23.42 2.14 20.11 2.14 20.11 2.68 17.97 2.68 17.97 2.595 15.015 2.595  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.715 1.8 17.675 1.8 17.675 1.45 21.88 1.45 21.88 1.68 17.925 1.68 17.925 2.12 15.715 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.8 1.35 1.8 1.35 1.34 8.17 1.34 8.17 1.77 9.47 1.77 9.47 2.12 7.94 2.12 7.94 1.57 1.59 1.57 1.59 2.12 0.62 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.84 1.8 7.71 1.8 7.71 2.12 1.84 2.12  ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 3.838 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.115 1.8 13.57 1.8 14.16 1.8 14.16 2.12 13.57 2.12 10.115 2.12  ;
    END
  END C
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.7442 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.69 2.825 17.465 2.825 17.465 2.91 20.505 2.91 20.505 2.825 23.78 2.825 23.78 3.055 20.735 3.055 20.735 3.31 17.235 3.31 17.235 3.055 14.35 3.055 14.35 2.68 13.57 2.68 12.395 2.68 12.395 3.11 12.165 3.11 12.165 2.68 10.255 2.68 10.255 3.11 10.025 3.11 10.025 2.68 9.435 2.68 9.435 3.11 9.205 3.11 9.205 2.68 4.955 2.68 4.955 3.11 4.725 3.11 4.725 2.68 0.575 2.68 0.575 3.11 0.345 3.11 0.345 2.36 13.57 2.36 14.405 2.36 14.405 0.99 22.53 0.99 22.53 1.22 14.69 1.22  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.43 3.62 2.43 3.09 2.77 3.09 2.77 3.62 6.91 3.62 6.91 3.09 7.25 3.09 7.25 3.62 10.99 3.62 10.99 3.09 11.33 3.09 11.33 3.62 13.23 3.62 13.23 3.09 13.57 3.09 13.57 3.62 16.59 3.62 16.59 3.285 16.93 3.285 16.93 3.62 21.07 3.62 21.07 3.285 21.41 3.285 21.41 3.62 23.88 3.62 24.08 3.62 24.08 4.22 23.88 4.22 13.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 24.08 -0.3 24.08 0.3 9.49 0.3 9.49 0.635 9.145 0.635 9.145 0.3 7.25 0.3 7.25 0.635 6.905 0.635 6.905 0.3 5.01 0.3 5.01 0.635 4.665 0.635 4.665 0.3 2.77 0.3 2.77 0.635 2.425 0.635 2.425 0.3 0.53 0.3 0.53 0.635 0.19 0.635 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.22 0.865 9.035 0.865 9.035 0.99 13.57 0.99 13.57 1.22 8.785 1.22 8.785 1.095 1.22 1.095  ;
        POLYGON 9.86 0.53 23.88 0.53 23.88 0.76 9.86 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai221_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai222_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai222_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.4 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.3 1.06 7.72 1.06 7.72 1.77 8.2 1.77 8.27 1.77 8.27 2.15 8.2 2.15 7.3 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.72 1.06 6.04 1.06 6.04 1.77 6.61 1.77 6.61 2.15 5.72 2.15  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.37 1.77 4.36 1.77 4.36 2.15 2.69 2.15 2.69 3.32 2.37 3.32  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.59 1.77 4.61 1.77 5.16 1.77 5.16 1.06 5.48 1.06 5.48 2.15 4.61 2.15 4.59 2.15  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 1.52 2.14 1.52 2.14 3.32 1.78 3.32  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.16 1.02 1.16 1.02 2.71 0.66 2.71  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.5684 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.055 2.9 4.61 2.9 4.755 2.9 4.755 2.74 6.84 2.74 6.84 1.22 6.51 1.22 6.51 0.99 7.07 0.99 7.07 2.74 8.1 2.74 8.1 3.26 6.035 3.26 6.035 2.97 5.065 2.97 5.065 3.26 4.61 3.26 3.055 3.26  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.95 0.575 2.95 0.575 3.62 4.61 3.62 5.445 3.62 5.445 3.2 5.675 3.2 5.675 3.62 8.2 3.62 8.4 3.62 8.4 4.22 8.2 4.22 4.61 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.4 -0.3 8.4 0.3 2.715 0.3 2.715 0.76 2.485 0.76 2.485 0.3 0.475 0.3 0.475 0.76 0.245 0.76 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.53 1.595 0.53 1.595 0.99 4.61 0.99 4.61 1.22 1.365 1.22  ;
        POLYGON 3.15 0.53 8.2 0.53 8.2 0.76 3.15 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai222_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai222_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai222_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.12 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.525 1.645 11.06 1.645 11.06 2.365 14.005 2.365 14.005 1.16 14.46 1.16 14.46 2.69 13.285 2.69 13.285 2.595 10.525 2.595  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.29 1.8 13.39 1.8 13.39 2.12 11.29 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.07 2.365 6.04 2.365 6.04 1.79 6.3 1.79 6.3 2.365 9.09 2.365 9.1 2.365 9.1 1.77 9.68 1.77 9.68 2.15 9.38 2.15 9.38 2.595 9.09 2.595 6.74 2.595 6.74 2.69 5.07 2.69  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.77 1.8 8.87 1.8 8.87 2.12 6.77 2.12  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.335 4.38 1.335 4.38 1.8 5.015 1.8 5.015 2.12 4.01 2.12 4.01 1.57 1.02 1.57 1.02 2.19 0.66 2.19  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.53 1.8 3.46 1.8 3.46 2.12 1.53 2.12  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.265 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.16 2.825 12.95 2.825 12.95 2.92 14.82 2.92 14.82 3.24 12.72 3.24 12.72 3.055 11.775 3.055 11.775 3.24 9.09 3.24 8.445 3.24 8.445 3.055 7.34 3.055 7.34 3.24 3.125 3.24 3.125 3.055 0.28 3.055 0.28 2.825 3.42 2.825 3.42 2.92 7.09 2.92 7.09 2.825 9.09 2.825 9.93 2.825 9.93 0.99 13.57 0.99 13.57 1.22 10.16 1.22  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.43 3.62 2.43 3.285 2.77 3.285 2.77 3.62 7.63 3.62 7.63 3.285 7.97 3.285 7.97 3.62 9.09 3.62 12.11 3.62 12.11 3.285 12.45 3.285 12.45 3.62 14.92 3.62 15.12 3.62 15.12 4.22 14.92 4.22 9.09 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 15.12 -0.3 15.12 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.475 0.3 0.475 0.845 0.245 0.845 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.31 0.865 5.13 0.865 5.13 0.99 9.09 0.99 9.09 1.22 4.88 1.22 4.88 1.095 1.31 1.095  ;
        POLYGON 5.39 0.53 14.92 0.53 14.92 0.76 5.39 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai222_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai222_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai222_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 28.56 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.49 1.79 19.73 1.79 19.73 2.35 22.8 2.35 22.8 1.95 23.14 1.95 23.14 2.35 23.82 2.35 23.82 1.95 24.16 1.95 24.16 2.35 27.42 2.35 27.42 1.72 27.715 1.72 27.715 2.58 24.8 2.58 24.8 2.68 22.16 2.68 22.16 2.58 19.49 2.58  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.21 1.8 22.07 1.8 22.07 1.47 24.97 1.47 24.97 1.8 26.83 1.8 26.83 2.12 24.69 2.12 24.69 1.7 22.35 1.7 22.35 2.12 20.21 2.12  ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.63 1.77 11.09 1.77 11.09 2.35 13.84 2.35 13.84 1.95 14.18 1.95 14.18 2.35 14.86 2.35 14.86 1.95 15.2 1.95 15.2 2.35 18.05 2.35 18.22 2.35 18.22 1.95 18.56 1.95 18.56 2.58 18.05 2.58 15.84 2.58 15.84 2.68 13.2 2.68 13.2 2.58 10.86 2.58 10.86 2.15 9.63 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.32 1.8 12.93 1.8 12.93 1.47 15.85 1.47 15.85 1.8 17.87 1.8 17.87 2.12 15.62 2.12 15.62 1.7 13.39 1.7 13.39 2.12 11.32 2.12  ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 1.255 1.77 1.255 1.33 8.515 1.33 8.515 1.77 9.4 1.77 9.4 2.15 8.2 2.15 8.2 1.56 1.57 1.56 1.57 2.15 0.28 2.15  ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.92 1.8 7.84 1.8 7.84 2.12 1.92 2.12  ;
    END
  END C2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 6.88075 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.12 2.82 21.91 2.82 21.91 2.92 25.05 2.92 25.05 2.82 27.965 2.82 27.965 2.53 28.195 2.53 28.195 3.38 27.965 3.38 27.965 3.05 25.3 3.05 25.3 3.24 21.66 3.24 21.66 3.05 19.12 3.05 19.12 3.38 18.81 3.38 18.81 3.05 18.05 3.05 16.34 3.05 16.34 3.24 12.7 3.24 12.7 3.05 6.66 3.05 6.66 3.24 4.955 3.24 4.955 3.38 4.725 3.38 4.725 3.24 3.02 3.24 3.02 3.05 0.525 3.05 0.525 3.38 0.295 3.38 0.295 2.53 0.525 2.53 0.525 2.82 4.725 2.82 4.725 2.53 4.955 2.53 4.955 2.82 12.95 2.82 12.95 2.92 16.09 2.92 16.09 2.82 18.05 2.82 18.81 2.82 18.81 0.99 27.01 0.99 27.01 1.22 19.12 1.22  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.43 3.62 2.43 3.28 2.77 3.28 2.77 3.62 6.91 3.62 6.91 3.285 7.25 3.285 7.25 3.62 12.11 3.62 12.11 3.285 12.45 3.285 12.45 3.62 16.59 3.62 16.59 3.285 16.93 3.285 16.93 3.62 18.05 3.62 21.07 3.62 21.07 3.285 21.41 3.285 21.41 3.62 25.55 3.62 25.55 3.285 25.89 3.285 25.89 3.62 28.36 3.62 28.56 3.62 28.56 4.22 28.36 4.22 18.05 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 28.56 -0.3 28.56 0.3 9.49 0.3 9.49 0.635 9.15 0.635 9.15 0.3 7.25 0.3 7.25 0.635 6.91 0.635 6.91 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.53 0.3 0.53 0.635 0.19 0.635 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.31 0.865 9.495 0.865 9.495 0.99 18.05 0.99 18.05 1.22 9.265 1.22 9.265 1.095 1.31 1.095  ;
        POLYGON 9.86 0.53 28.36 0.53 28.36 0.76 9.86 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai222_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai31_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai31_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.16 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0365 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.23 1.75 1.79 1.75 1.79 1.16 2.13 1.16 2.13 2.15 1.23 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0365 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.47 1.47 3.81 1.47 3.81 3.32 3.47 3.32  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0365 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.59 1.47 4.935 1.47 4.935 3.32 4.59 3.32  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.054 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.16 1 1.16 1 3.32 0.705 3.32  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.9884 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.33 2.38 2.36 2.38 2.36 0.99 4.33 0.99 5.165 0.99 5.165 0.605 5.395 0.605 5.395 1.22 4.33 1.22 2.68 1.22 2.68 2.68 1.67 2.68 1.67 3.38 1.33 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 4.33 3.62 5.165 3.62 5.165 2.53 5.395 2.53 5.395 3.62 6.16 3.62 6.16 4.22 4.33 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.16 -0.3 6.16 0.3 0.475 0.3 0.475 0.945 0.245 0.945 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.31 0.53 4.33 0.53 4.33 0.76 1.31 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai31_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai31_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai31_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.64 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.42 1.665 6.745 1.665 6.745 1.45 8.97 1.45 8.97 1.21 9.94 1.21 9.98 1.21 9.98 2.28 9.94 2.28 9.62 2.28 9.62 1.68 6.975 1.68 6.975 1.985 5.42 1.985  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.03 1.77 4.99 1.77 4.99 2.235 7.67 2.235 7.67 1.91 8.35 1.91 8.35 2.69 7.255 2.69 7.255 2.465 4.46 2.465 4.46 2.15 4.03 2.15  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.97 1.77 3.8 1.77 3.8 2.695 6.85 2.695 6.85 2.92 9.01 2.92 9.01 1.91 9.24 1.91 9.24 3.26 6.6 3.26 6.6 2.93 3.47 2.93 3.47 2.12 2.97 2.12  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.064 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.77 2.13 1.77 2.13 2.15 0.28 2.15  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.796 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 2.53 2.36 2.53 2.36 0.99 8.6 0.99 8.6 1.22 2.68 1.22 2.68 2.53 3.2 2.53 3.2 3.16 6.35 3.16 6.35 3.39 2.97 3.39 2.97 2.76 1.595 2.76 1.595 3.375 1.365 3.375  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.295 3.62 0.295 2.53 0.525 2.53 0.525 3.62 2.33 3.62 2.33 3.02 2.67 3.02 2.67 3.62 9.49 3.62 9.49 2.53 9.83 2.53 9.83 3.62 9.94 3.62 10.64 3.62 10.64 4.22 9.94 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.64 -0.3 10.64 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.865 1.9 0.865 1.9 0.53 9.94 0.53 9.94 0.76 2.13 0.76 2.13 1.095 0.18 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai31_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai31_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai31_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 19.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.48 1.77 4.69 1.77 4.69 1.45 12.42 1.45 12.42 1.68 4.92 1.68 4.92 2.15 3.48 2.15  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.15 2.22 5.42 2.22 5.42 1.91 5.92 1.91 5.92 2.22 8.86 2.22 8.86 1.91 10.22 1.91 10.22 2.22 12.97 2.22 12.97 1.725 13.89 1.725 13.89 2.45 6.775 2.45 6.775 2.71 5.15 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.68 3.24 1.68 3.24 2.15 0.62 2.15  ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.89 1.785 19.15 1.785 19.15 2.12 14.89 2.12  ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.0289 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.13 2.7 14.12 2.7 14.12 1.22 1.31 1.22 1.31 0.99 14.44 0.99 14.44 2.36 18.43 2.36 18.43 2.93 7.13 2.93  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.53 3.62 1.53 3.285 1.87 3.285 1.87 3.62 3.77 3.62 3.77 3.285 4.11 3.285 4.11 3.62 14.1 3.62 14.47 3.62 14.47 3.285 14.81 3.285 14.81 3.62 16.61 3.62 16.61 3.285 16.95 3.285 16.95 3.62 18.855 3.62 18.855 2.57 19.085 2.57 19.085 3.62 19.2 3.62 19.6 3.62 19.6 4.22 19.2 4.22 14.1 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 19.6 -0.3 19.6 0.3 18.07 0.3 18.07 0.635 17.73 0.635 17.73 0.3 15.83 0.3 15.83 0.635 15.49 0.635 15.49 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.57 4.59 2.57 4.59 3.16 14.1 3.16 14.1 3.39 4.36 3.39 4.36 2.8 2.935 2.8 2.935 3.38 2.705 3.38 2.705 2.8 0.575 2.8 0.575 3.38 0.345 3.38  ;
        POLYGON 0.18 0.53 15.21 0.53 15.21 0.865 19.2 0.865 19.2 1.095 14.98 1.095 14.98 0.76 0.18 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai31_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai32_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai32_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 1.73 3.83 1.73 3.83 2.15 3.24 2.15 3.24 2.75 2.92 2.75  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.65 2.12 1.65 2.12 3.31 1.8 3.31  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.65 1 1.65 1 3.31 0.705 3.31  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.065 0.61 4.37 0.61 4.37 2.15 4.065 2.15  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.185 0.61 5.49 0.61 5.49 2.19 5.185 2.19  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.3048 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.47 2.38 4.6 2.38 4.6 0.61 4.955 0.61 4.955 2.7 3.47 2.7  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.59 0.475 2.59 0.475 3.62 5.745 3.62 5.745 3.2 5.975 3.2 5.975 3.62 6.075 3.62 6.72 3.62 6.72 4.22 6.075 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.72 -0.3 6.72 0.3 2.715 0.3 2.715 0.915 2.485 0.915 2.485 0.3 0.475 0.3 0.475 0.915 0.245 0.915 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.68 3.05 5.22 3.05 5.22 2.64 5.845 2.64 5.845 0.61 6.075 0.61 6.075 2.87 5.45 2.87 5.45 3.28 2.45 3.28 2.45 1.4 1.365 1.4 1.365 0.61 1.595 0.61 1.595 1.165 3.605 1.165 3.605 0.61 3.835 0.61 3.835 1.4 2.68 1.4  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai32_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai32_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai32_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.88 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.85 1.8 4.39 1.8 4.39 2.12 2.85 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.535 1.77 2.35 1.77 2.35 1.325 4.85 1.325 4.85 1.77 6.07 1.77 6.07 2.12 4.62 2.12 4.62 1.555 2.6 1.555 2.6 2.135 1.535 2.135  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 1.56 1.145 1.56 1.145 2.365 6.3 2.365 6.3 1.56 6.6 1.56 6.6 2.595 6.16 2.595 6.16 2.68 0.825 2.68  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.45 1.8 10.59 1.8 10.59 2.12 8.45 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.56 1.785 7.88 1.785 7.88 2.365 11.215 2.365 11.215 1.56 11.535 1.56 11.535 2.68 8.12 2.68 8.12 2.595 7.56 2.595  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3774 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 2.92 6.41 2.92 6.41 2.825 6.84 2.825 6.84 0.99 10.84 0.99 10.84 1.22 7.16 1.22 7.16 2.825 7.75 2.825 7.75 2.92 10.17 2.92 10.17 3.24 7.5 3.24 7.5 3.055 6.66 3.055 6.66 3.24 3.365 3.24  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.65 0.575 2.65 0.575 3.62 6.91 3.62 6.91 3.285 7.25 3.285 7.25 3.62 11.785 3.62 11.785 2.65 12.015 2.65 12.015 3.62 12.18 3.62 12.88 3.62 12.88 4.22 12.18 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.88 -0.3 12.88 0.3 6.13 0.3 6.13 0.635 5.79 0.635 5.79 0.3 3.89 0.3 3.89 0.635 3.55 0.635 3.55 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.865 6.37 0.865 6.37 0.53 12.18 0.53 12.18 0.76 6.6 0.76 6.6 1.095 0.18 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai32_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai32_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai32_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 24.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.57 1.8 13.88 1.8 13.88 2.12 9.57 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.055 1.76 1.295 1.76 1.295 2.35 4.365 2.35 4.365 1.825 5.725 1.825 5.725 2.35 8.895 2.35 8.895 1.76 9.135 1.76 9.135 2.58 6.365 2.58 6.365 2.69 3.73 2.69 3.73 2.58 1.055 2.58  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.73 1.8 3.64 1.8 3.64 1.345 6.44 1.345 6.44 1.8 8.35 1.8 8.35 2.12 6.21 2.12 6.21 1.575 3.87 1.575 3.87 2.12 1.73 2.12  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.005 1.8 17.64 1.8 17.64 1.45 20.44 1.45 20.44 1.8 22.35 1.8 22.35 2.12 20.21 2.12 20.21 1.68 17.87 1.68 17.87 2.12 16.005 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.65 1.8 15.775 1.8 15.775 2.36 18.325 2.36 18.325 1.91 19.685 1.91 19.685 2.36 22.965 2.36 22.965 1.76 23.225 1.76 23.225 2.68 19.945 2.68 19.945 2.595 18.05 2.595 18.05 2.68 15.545 2.68 15.545 2.12 14.65 2.12  ;
    END
  END B2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 4.1761 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.57 2.36 14.12 2.36 14.12 0.99 22.535 0.99 22.535 1.22 14.42 1.22 14.42 2.36 15.295 2.36 15.295 2.92 18.335 2.92 18.335 2.825 19.655 2.825 19.655 2.92 21.81 2.92 21.81 3.24 19.425 3.24 19.425 3.055 18.585 3.055 18.585 3.24 15.045 3.24 15.045 2.815 9.57 2.815  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.635 3.62 2.635 3.285 2.975 3.285 2.975 3.62 7.115 3.62 7.115 3.285 7.455 3.285 7.455 3.62 14.085 3.62 14.455 3.62 14.455 3.285 14.795 3.285 14.795 3.62 18.835 3.62 18.835 3.285 19.175 3.285 19.175 3.62 23.5 3.62 23.5 2.53 23.73 2.53 23.73 3.62 23.885 3.62 24.08 3.62 24.08 4.22 23.885 4.22 14.085 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 24.08 -0.3 24.08 0.3 13.055 0.3 13.055 0.635 12.715 0.635 12.715 0.3 10.815 0.3 10.815 0.635 10.475 0.635 10.475 0.3 8.575 0.3 8.575 0.635 8.235 0.635 8.235 0.3 6.335 0.3 6.335 0.635 5.995 0.635 5.995 0.3 4.095 0.3 4.095 0.635 3.755 0.635 3.755 0.3 1.855 0.3 1.855 0.635 1.515 0.635 1.515 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.5 2.53 0.73 2.53 0.73 2.825 3.48 2.825 3.48 2.94 6.615 2.94 6.615 2.825 8.42 2.825 8.42 3.14 14.085 3.14 14.085 3.37 8.19 3.37 8.19 3.055 6.865 3.055 6.865 3.17 3.23 3.17 3.23 3.055 0.73 3.055 0.73 3.38 0.5 3.38  ;
        POLYGON 0.385 0.865 13.405 0.865 13.405 0.53 23.885 0.53 23.885 0.76 13.635 0.76 13.635 1.095 0.385 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai32_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai33_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai33_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 8.4 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.04 1.525 4.36 1.525 4.36 3.32 4.04 3.32  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.16 1.77 6.04 1.77 6.04 2.14 5.48 2.14 5.48 3.32 5.16 3.32  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.28 1.77 6.57 1.77 7.87 1.77 7.87 2.14 6.6 2.14 6.6 3.32 6.57 3.32 6.28 3.32  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 1.525 3.24 1.525 3.24 3.32 2.92 3.32  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.525 2.12 1.525 2.12 3.32 1.8 3.32  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0395 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 1.525 1 1.525 1 3.32 0.705 3.32  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.8719 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.49 0.99 6.57 0.99 7.405 0.99 7.405 0.555 7.635 0.555 7.635 1.22 6.57 1.22 3.79 1.22 3.79 3.38 3.49 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.245 3.62 0.245 2.53 0.475 2.53 0.475 3.62 6.57 3.62 7.305 3.62 7.305 2.53 7.535 2.53 7.535 3.62 8.4 3.62 8.4 4.22 6.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 8.4 -0.3 8.4 0.3 2.715 0.3 2.715 0.815 2.485 0.815 2.485 0.3 0.475 0.3 0.475 0.815 0.245 0.815 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.365 0.53 1.595 0.53 1.595 1.045 2.945 1.045 2.945 0.53 6.57 0.53 6.57 0.76 3.175 0.76 3.175 1.275 1.365 1.275  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai33_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai33_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai33_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.12 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.8 1.45 13.38 1.45 13.38 1.16 14.42 1.16 14.44 1.16 14.44 2.38 14.42 2.38 14.12 2.38 14.12 1.68 9.8 1.68  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.48 1.78 9.52 1.78 9.52 1.91 12.54 1.91 12.54 2.14 8.48 2.14  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.44 1.78 8.23 1.78 8.23 2.37 13.435 2.37 13.435 1.91 13.775 1.91 13.775 2.68 8 2.68 8 2.14 7.44 2.14  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.8 4.95 1.8 4.95 2.12 2.89 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.51 1.77 2.41 1.77 2.41 1.325 5.48 1.325 5.48 2.15 5.18 2.15 5.18 1.555 2.66 1.555 2.66 2.15 1.51 2.15  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.079 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.8 1.145 1.8 1.145 2.38 5.72 2.38 5.72 1.8 6.6 1.8 6.6 2.12 6.06 2.12 6.06 2.68 0.825 2.68 0.825 2.12 0.28 2.12  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.8038 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.75 2.92 6.41 2.92 6.41 2.825 6.85 2.825 6.85 0.99 13.07 0.99 13.07 1.22 7.15 1.22 7.15 2.825 7.75 2.825 7.75 2.92 11.215 2.92 11.215 3.24 7.5 3.24 7.5 3.055 6.66 3.055 6.66 3.24 2.75 3.24  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.63 0.575 2.63 0.575 3.62 6.91 3.62 6.91 3.285 7.25 3.285 7.25 3.62 14.025 3.62 14.025 2.63 14.255 2.63 14.255 3.62 14.42 3.62 15.12 3.62 15.12 4.22 14.42 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 15.12 -0.3 15.12 0.3 6.13 0.3 6.13 0.635 5.79 0.635 5.79 0.3 3.89 0.3 3.89 0.635 3.55 0.635 3.55 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 0.865 6.38 0.865 6.38 0.53 14.42 0.53 14.42 0.76 6.61 0.76 6.61 1.095 0.18 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai33_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__oai33_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__oai33_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 28.56 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.58 1.8 18.44 1.8 18.44 2.12 14.58 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.29 1.76 19.53 1.76 19.53 2.36 22.6 2.36 22.6 1.92 23.96 1.92 23.96 2.36 27.25 2.36 27.25 1.76 27.49 1.76 27.49 2.59 24.605 2.59 24.605 2.71 21.955 2.71 21.955 2.59 19.29 2.59  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.18 1.8 21.685 1.8 21.685 1.45 24.775 1.45 24.775 1.8 26.835 1.8 26.835 2.12 24.545 2.12 24.545 1.68 21.915 1.68 21.915 2.12 20.18 2.12  ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.58 1.8 13.34 1.8 13.34 2.12 9.58 2.12  ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.775 1.53 1.095 1.53 1.095 2.36 4.16 2.36 4.16 1.92 5.52 1.92 5.52 2.36 8.58 2.36 8.58 1.76 8.84 1.76 8.84 2.595 6.16 2.595 6.16 2.7 3.52 2.7 3.52 2.595 0.775 2.595  ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 4.158 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.8 3.59 1.8 3.59 1.335 6.45 1.335 6.45 1.8 8.31 1.8 8.31 2.12 6.22 2.12 6.22 1.565 3.82 1.565 3.82 2.12 1.74 2.12  ;
    END
  END B3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 5.0289 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.58 2.36 13.57 2.36 13.57 0.99 26.82 0.99 26.82 1.22 13.87 1.22 13.87 2.36 17.89 2.36 17.89 2.795 9.58 2.795  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.43 3.62 2.43 3.285 2.77 3.285 2.77 3.62 6.91 3.62 6.91 3.285 7.25 3.285 7.25 3.62 13.87 3.62 20.87 3.62 20.87 3.285 21.21 3.285 21.21 3.62 25.35 3.62 25.35 3.285 25.69 3.285 25.69 3.62 27.995 3.62 28.16 3.62 28.56 3.62 28.56 4.22 28.16 4.22 27.995 4.22 13.87 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 28.56 -0.3 28.56 0.3 12.85 0.3 12.85 0.635 12.51 0.635 12.51 0.3 10.61 0.3 10.61 0.635 10.27 0.635 10.27 0.3 8.37 0.3 8.37 0.635 8.03 0.635 8.03 0.3 6.13 0.3 6.13 0.635 5.79 0.635 5.79 0.3 3.89 0.3 3.89 0.635 3.55 0.635 3.55 0.3 1.65 0.3 1.65 0.635 1.31 0.635 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.295 2.53 0.525 2.53 0.525 2.825 3.27 2.825 3.27 3.09 6.41 3.09 6.41 2.825 7.73 2.825 7.73 3.09 13.87 3.09 13.87 3.32 7.5 3.32 7.5 3.055 6.66 3.055 6.66 3.32 3.02 3.32 3.02 3.055 0.525 3.055 0.525 3.38 0.295 3.38  ;
        POLYGON 14.24 3.09 20.11 3.09 20.11 2.825 21.705 2.825 21.705 3.09 24.855 3.09 24.855 2.825 27.765 2.825 27.765 2.53 27.995 2.53 27.995 3.38 27.765 3.38 27.765 3.055 25.1 3.055 25.1 3.32 21.46 3.32 21.46 3.055 20.355 3.055 20.355 3.32 14.24 3.32  ;
        POLYGON 0.18 0.865 13.1 0.865 13.1 0.53 28.16 0.53 28.16 0.76 13.33 0.76 13.33 1.095 0.18 1.095  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__oai33_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 4.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4985 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.075 1.08 1.075 1.08 2.88 0.66 2.88  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.4985 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 1.74 2.14 1.74 2.14 3.345 1.78 3.345  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.5 2.29 3.535 2.29 3.8 2.29 3.8 1.04 3.365 1.04 3.365 0.61 4.13 0.61 4.13 3.345 3.535 3.345 3.5 3.345  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.78 3.62 2.78 2.53 3.01 2.53 3.01 3.62 3.535 3.62 4.48 3.62 4.48 4.22 3.535 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 4.48 -0.3 4.48 0.3 3.01 0.3 3.01 0.85 2.78 0.85 2.78 0.3 0.53 0.3 0.53 0.825 0.3 0.825 0.3 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.335 3.13 1.31 3.13 1.31 0.53 1.705 0.53 1.705 1.28 3.535 1.28 3.535 1.64 2.68 1.64 2.68 1.51 1.54 1.51 1.54 3.36 0.335 3.36  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or2_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.015 1.02 1.015 1.02 2.28 0.66 2.28  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.102 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 1.43 2.14 1.43 2.14 3.39 1.78 3.39  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1218 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.48 0.53 3.835 0.53 3.835 3.39 3.48 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.435 3.62 2.435 2.53 2.665 2.53 2.665 3.62 3.205 3.62 4.625 3.62 4.625 2.53 4.855 2.53 4.855 3.62 5.6 3.62 5.6 4.22 3.205 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 4.955 0.3 4.955 1.045 4.725 1.045 4.725 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.53 0.3 0.53 0.635 0.19 0.635 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.53 1.3 2.53 1.3 0.53 1.595 0.53 1.595 0.885 3.205 0.885 3.205 2.115 2.975 2.115 2.975 1.115 1.53 1.115 1.53 2.765 0.575 2.765 0.575 3.39 0.345 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or2_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.595 1.8 3.5 1.8 3.5 2.12 1.595 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.204 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 1.765 1.21 1.765 1.21 2.36 3.93 2.36 3.93 1.825 4.275 1.825 4.275 2.68 0.87 2.68  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3046 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.085 2.36 8.96 2.36 9.205 2.36 9.205 1.54 5.985 1.54 5.985 0.53 6.215 0.53 6.215 1.26 8.225 1.26 8.225 0.53 8.455 0.53 8.455 1.265 9.46 1.265 9.46 2.68 8.96 2.68 8.405 2.68 8.405 3.39 8.175 3.39 8.175 2.68 6.315 2.68 6.315 3.39 6.085 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.575 2.53 0.575 3.62 4.965 3.62 4.965 2.53 5.195 2.53 5.195 3.62 7.105 3.62 7.105 2.935 7.335 2.935 7.335 3.62 8.96 3.62 9.245 3.62 9.245 2.94 9.475 2.94 9.475 3.62 10.08 3.62 10.08 4.22 8.96 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.575 0.3 9.575 0.98 9.345 0.98 9.345 0.3 7.335 0.3 7.335 0.985 7.105 0.985 7.105 0.3 4.955 0.3 4.955 1.07 4.725 1.07 4.725 0.3 2.715 0.3 2.715 1.07 2.485 1.07 2.485 0.3 0.475 0.3 0.475 1.07 0.245 1.07 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 2.35 2.945 4.505 2.945 4.505 1.57 1.365 1.57 1.365 0.53 1.595 0.53 1.595 1.325 3.605 1.325 3.605 0.53 3.835 0.53 3.835 1.325 4.735 1.325 4.735 1.825 8.96 1.825 8.96 2.095 4.735 2.095 4.735 3.215 2.35 3.215  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or2_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 5.6 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.52 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.595 1.02 1.595 1.02 2.855 0.66 2.855  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.52 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 1.595 2.14 1.595 2.14 3.39 1.78 3.39  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.52 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.9 1.595 3.35 1.595 3.35 3.39 2.9 3.39  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.985 0.53 5.455 0.53 5.455 3.39 4.985 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 3.965 3.62 3.965 2.53 4.195 2.53 4.195 3.62 4.675 3.62 5.6 3.62 5.6 4.22 4.675 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 5.6 -0.3 5.6 0.3 4.07 0.3 4.07 0.735 3.73 0.735 3.73 0.3 1.65 0.3 1.65 0.735 1.31 0.735 1.31 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.18 3.16 1.285 3.16 1.285 1.2 0.19 1.2 0.19 0.53 0.53 0.53 0.53 0.965 2.43 0.965 2.43 0.53 2.77 0.53 2.77 0.965 4.675 0.965 4.675 2.22 4.445 2.22 4.445 1.2 1.515 1.2 1.515 3.39 0.18 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or3_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.009 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 1.73 1.56 1.73 1.56 3.38 1.22 3.38 1.22 2.14 0.84 2.14  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.009 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.79 1.61 2.14 1.61 2.14 3.38 1.79 3.38  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.009 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.9 1.61 3.26 1.61 3.26 3.38 2.9 3.38  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.84 2.38 5.515 2.38 5.745 2.38 5.745 1.535 4.87 1.535 4.87 0.53 5.49 0.53 5.49 1.265 6.04 1.265 6.04 2.655 5.515 2.655 5.46 2.655 5.46 3.38 4.84 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 3.715 3.62 3.715 2.53 3.945 2.53 3.945 3.62 5.515 3.62 5.925 3.62 5.925 2.935 6.155 2.935 6.155 3.62 6.72 3.62 6.72 4.22 5.515 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.72 -0.3 6.72 0.3 6.255 0.3 6.255 0.92 6.025 0.92 6.025 0.3 3.835 0.3 3.835 0.895 3.605 0.895 3.605 0.3 1.595 0.3 1.595 0.895 1.365 0.895 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.53 0.475 0.53 0.475 1.125 2.485 1.125 2.485 0.53 2.715 0.53 2.715 1.125 4.19 1.125 4.19 1.765 5.515 1.765 5.515 1.995 3.96 1.995 3.96 1.36 0.575 1.36 0.575 3.39 0.245 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or3_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.91 1.325 3.495 1.325 3.495 1.17 3.785 1.17 3.785 1.325 5.735 1.325 5.735 1.17 6.105 1.17 6.105 1.59 2.91 1.59  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.53 1.82 5.55 1.82 5.55 2.105 1.53 2.105  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 2.018 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 1.82 1.16 1.82 1.16 2.38 5.945 2.38 5.945 1.82 6.57 1.82 6.57 2.115 6.175 2.115 6.175 2.655 0.87 2.655  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2436 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.315 2.36 11.095 2.36 11.345 2.36 11.345 1.535 8.265 1.535 8.265 0.53 8.495 0.53 8.495 1.265 10.505 1.265 10.505 0.53 10.735 0.53 10.735 1.265 11.62 1.265 11.62 2.68 11.095 2.68 10.685 2.68 10.685 3.39 10.455 3.39 10.455 2.68 8.545 2.68 8.545 3.39 8.315 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.53 0.575 2.53 0.575 3.62 6.865 3.62 6.865 3.06 7.095 3.06 7.095 3.62 9.335 3.62 9.335 3 9.565 3 9.565 3.62 11.095 3.62 11.525 3.62 11.525 3 11.755 3 11.755 3.62 12.32 3.62 12.32 4.22 11.095 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 11.855 0.3 11.855 0.97 11.625 0.97 11.625 0.3 9.615 0.3 9.615 0.9 9.385 0.9 9.385 0.3 7.25 0.3 7.25 0.635 6.91 0.635 6.91 0.3 5.01 0.3 5.01 0.635 4.67 0.635 4.67 0.3 2.77 0.3 2.77 0.635 2.43 0.635 2.43 0.3 0.475 0.3 0.475 1.005 0.245 1.005 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 3.505 2.935 6.405 2.935 6.405 2.52 6.8 2.52 6.8 1.095 6.36 1.095 6.36 0.92 5.495 0.92 5.495 1.095 4.19 1.095 4.19 0.92 3.26 0.92 3.26 1.095 1.94 1.095 1.94 0.775 1.265 0.775 1.265 0.545 2.185 0.545 2.185 0.865 3.015 0.865 3.015 0.545 4.43 0.545 4.43 0.865 5.26 0.865 5.26 0.545 6.62 0.545 6.62 0.865 7.03 0.865 7.03 1.765 11.095 1.765 11.095 1.995 7.03 1.995 7.03 2.755 6.635 2.755 6.635 3.22 3.505 3.22  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or3_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or4_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or4_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.085 1.02 1.085 1.02 2.87 0.66 2.87  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 1.58 2.26 1.58 2.26 3.28 1.78 3.28  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.9 1.58 3.38 1.58 3.38 3.28 2.9 3.28  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.496 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.02 1.58 4.5 1.58 4.5 3.28 4.02 3.28  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.07 0.63 6.575 0.63 6.575 3.38 6.07 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 5.085 3.62 5.085 2.53 5.315 2.53 5.315 3.62 5.765 3.62 6.72 3.62 6.72 4.22 5.765 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.72 -0.3 6.72 0.3 5.315 0.3 5.315 0.855 5.085 0.855 5.085 0.3 2.95 0.3 2.95 0.76 2.61 0.76 2.61 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.28 3.12 1.3 3.12 1.3 1.095 1.49 1.095 1.49 0.53 1.83 0.53 1.83 1.095 3.73 1.095 3.73 0.53 4.07 0.53 4.07 1.095 5.765 1.095 5.765 2.27 5.515 2.27 5.515 1.33 1.53 1.33 1.53 3.35 0.28 3.35  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or4_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or4_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or4_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.84 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.015 1.02 1.015 1.02 2.29 0.66 2.29  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.78 1.48 2.14 1.48 2.14 3.39 1.78 3.39  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.9 1.48 3.26 1.48 3.26 3.39 2.9 3.39  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.889 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.02 1.48 4.38 1.48 4.38 3.39 4.02 3.39  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1218 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.97 2.36 6.75 2.36 7.01 2.36 7.01 1.56 6.025 1.56 6.025 0.53 6.585 0.53 6.585 1.24 7.28 1.24 7.28 2.68 6.75 2.68 6.585 2.68 6.585 3.39 5.97 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 4.82 3.62 4.82 2.53 5.05 2.53 5.05 3.62 6.75 3.62 7.045 3.62 7.045 2.99 7.275 2.99 7.275 3.62 7.84 3.62 7.84 4.22 6.75 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.84 -0.3 7.84 0.3 7.375 0.3 7.375 0.9 7.145 0.9 7.145 0.3 5.01 0.3 5.01 0.655 4.67 0.655 4.67 0.3 2.77 0.3 2.77 0.655 2.43 0.655 2.43 0.3 0.53 0.3 0.53 0.655 0.19 0.655 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 2.53 1.31 2.53 1.31 0.53 1.65 0.53 1.65 0.945 3.55 0.945 3.55 0.53 3.89 0.53 3.89 0.945 5.26 0.945 5.26 1.845 6.75 1.845 6.75 2.075 5.03 2.075 5.03 1.18 1.54 1.18 1.54 2.76 0.575 2.76 0.575 3.39 0.345 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or4_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__or4_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__or4_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 14.56 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.405 1.205 4.025 1.205 4.025 1.545 3.405 1.545  ;
        POLYGON 5.645 1.205 6.275 1.205 6.275 1.545 5.645 1.545  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.33 1.78 6.73 1.78 6.73 2.01 3.535 2.01 3.535 2.12 2.33 2.12  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.785 1.575 2.1 1.575 2.1 2.36 3.765 2.36 3.765 2.24 7.41 2.24 7.41 1.665 7.72 1.665 7.72 2.47 3.98 2.47 3.98 2.68 1.785 2.68  ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.778 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 1.765 1.21 1.765 1.21 2.92 4.21 2.92 4.21 2.7 7.96 2.7 7.96 1.4 8.885 1.4 8.885 1.63 8.31 1.63 8.31 2.93 4.44 2.93 4.44 3.24 0.87 3.24  ;
    END
  END A4
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3046 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.49 2.36 13.47 2.36 13.73 2.36 13.73 1.56 10.505 1.56 10.505 0.615 10.735 0.615 10.735 1.24 12.745 1.24 12.745 0.615 12.975 0.615 12.975 1.24 13.97 1.24 13.97 2.68 13.47 2.68 12.875 2.68 12.875 3.38 12.645 3.38 12.645 2.68 10.75 2.68 10.75 3.38 10.49 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.555 0.575 2.555 0.575 3.62 9.38 3.62 9.38 2.53 9.61 2.53 9.61 3.62 11.575 3.62 11.575 3.04 11.805 3.04 11.805 3.62 13.47 3.62 13.765 3.62 13.765 3.04 13.995 3.04 13.995 3.62 14.56 3.62 14.56 4.22 13.47 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 14.56 -0.3 14.56 0.3 14.095 0.3 14.095 0.83 13.865 0.83 13.865 0.3 11.855 0.3 11.855 0.83 11.625 0.83 11.625 0.3 9.49 0.3 9.49 0.655 9.15 0.655 9.15 0.3 7.195 0.3 7.195 0.71 6.965 0.71 6.965 0.3 4.955 0.3 4.955 0.71 4.725 0.71 4.725 0.3 2.715 0.3 2.715 0.71 2.485 0.71 2.485 0.3 0.53 0.3 0.53 0.655 0.19 0.655 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 4.67 3.16 8.78 3.16 8.78 1.88 9.195 1.88 9.195 1.17 6.505 1.17 6.505 0.76 5.415 0.76 5.415 1.17 4.26 1.17 4.26 0.76 3.175 0.76 3.175 1.17 1.31 1.17 1.31 0.53 1.65 0.53 1.65 0.94 2.945 0.94 2.945 0.53 4.49 0.53 4.49 0.94 5.185 0.94 5.185 0.53 6.735 0.53 6.735 0.94 8.03 0.94 8.03 0.53 8.37 0.53 8.37 0.94 9.425 0.94 9.425 1.79 13.47 1.79 13.47 2.13 9.04 2.13 9.04 3.39 4.67 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__or4_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 21.28 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.795 5.085 1.795 5.085 2.215 3.41 2.215  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.739 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.465 1.795 6.63 1.795 6.63 2.2 5.465 2.2  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8932 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.79 0.615 21.15 0.615 21.15 3.365 20.79 3.365  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 2.775 3.62 5.25 3.62 5.25 3.18 5.59 3.18 5.59 3.62 7.57 3.62 7.57 3.35 7.91 3.35 7.91 3.62 10.015 3.62 12.93 3.62 12.93 2.995 13.27 2.995 13.27 3.62 16.245 3.62 17.25 3.62 17.25 2.845 17.59 2.845 17.59 3.62 18.17 3.62 19.735 3.62 19.735 2.46 19.965 2.46 19.965 3.62 20.54 3.62 21.28 3.62 21.28 4.22 20.54 4.22 18.17 4.22 16.245 4.22 10.015 4.22 2.775 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 21.28 -0.3 21.28 0.3 19.915 0.3 19.915 0.995 19.685 0.995 19.685 0.3 17.855 0.3 17.855 0.68 17.625 0.68 17.625 0.3 13.32 0.3 13.32 1.085 12.98 1.085 12.98 0.3 8.01 0.3 8.01 1.045 7.78 1.045 7.78 0.3 5.635 0.3 5.635 1.075 5.295 1.075 5.295 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.79 0.475 0.79 0.475 2.385 2.545 2.385 2.545 1.625 2.775 1.625 2.775 2.615 0.475 2.615 0.475 3.015 0.245 3.015  ;
        POLYGON 6.585 2.43 6.86 2.43 6.86 1.275 6.75 1.275 6.75 0.99 7.09 0.99 7.09 2.43 8.37 2.43 8.37 1.875 8.6 1.875 8.6 2.66 6.815 2.66 6.815 2.86 6.585 2.86  ;
        POLYGON 3.03 2.705 6.105 2.705 6.105 3.09 7.09 3.09 7.09 2.89 8.6 2.89 8.6 3.12 9.785 3.12 9.785 2.69 10.015 2.69 10.015 3.35 8.37 3.35 8.37 3.12 7.32 3.12 7.32 3.32 5.875 3.32 5.875 2.935 3.03 2.935  ;
        POLYGON 3.27 0.845 4.655 0.845 4.655 1.305 6.09 1.305 6.09 0.53 7.55 0.53 7.55 1.305 8.375 1.305 8.375 0.53 10.07 0.53 10.07 1.14 9.84 1.14 9.84 0.76 8.605 0.76 8.605 1.535 7.32 1.535 7.32 0.76 6.32 0.76 6.32 1.535 4.425 1.535 4.425 1.075 3.27 1.075  ;
        POLYGON 10.855 1.47 10.96 1.47 10.96 0.8 11.19 0.8 11.19 1.47 13.965 1.47 13.965 1.7 11.085 1.7 11.085 2.87 10.855 2.87  ;
        POLYGON 12.2 2.07 14.325 2.07 14.325 0.8 14.555 0.8 14.555 2.87 14.325 2.87 14.325 2.3 12.2 2.3  ;
        POLYGON 9.295 1.82 10.555 1.82 10.555 3.15 12.26 3.15 12.26 2.53 13.9 2.53 13.9 3.16 14.785 3.16 14.785 1.26 15.015 1.26 15.015 3.16 15.905 3.16 15.905 2.07 16.245 2.07 16.245 3.39 13.67 3.39 13.67 2.765 12.49 2.765 12.49 3.39 10.325 3.39 10.325 2.05 9.13 2.05 9.13 2.86 8.9 2.86 8.9 1.82 9.065 1.82 9.065 0.99 9.405 0.99 9.405 1.275 9.295 1.275  ;
        POLYGON 15.445 0.8 15.675 0.8 15.675 1.54 16.735 1.54 16.735 2.315 17.83 2.315 17.83 1.67 18.17 1.67 18.17 2.55 16.505 2.55 16.505 1.775 15.675 1.775 15.675 2.87 15.445 2.87  ;
        POLYGON 18.465 1.78 18.965 1.78 18.965 1.23 17.195 1.23 17.195 1.6 16.965 1.6 16.965 0.995 18.965 0.995 18.965 0.76 19.195 0.76 19.195 1.78 20.54 1.78 20.54 2.01 18.695 2.01 18.695 2.95 18.465 2.95  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 22.4 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.795 5.14 1.795 5.14 2.215 3.41 2.215  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.739 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.465 1.795 6.63 1.795 6.63 2.2 5.465 2.2  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.11635 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.76 0.615 21.18 0.615 21.18 3.39 20.76 3.39  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 2.775 3.62 5.25 3.62 5.25 3.18 5.59 3.18 5.59 3.62 7.57 3.62 7.57 3.35 7.91 3.35 7.91 3.62 10.015 3.62 12.93 3.62 12.93 2.995 13.27 2.995 13.27 3.62 16.245 3.62 17.71 3.62 17.71 2.8 18.05 2.8 18.05 3.62 18.63 3.62 19.785 3.62 19.785 2.46 20.015 2.46 20.015 3.62 20.515 3.62 21.875 3.62 21.875 2.46 22.105 2.46 22.105 3.62 22.4 3.62 22.4 4.22 20.515 4.22 18.63 4.22 16.245 4.22 10.015 4.22 2.775 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 22.4 -0.3 22.4 0.3 22.155 0.3 22.155 0.95 21.925 0.95 21.925 0.3 19.915 0.3 19.915 0.95 19.685 0.95 19.685 0.3 18.075 0.3 18.075 0.725 17.845 0.725 17.845 0.3 13.32 0.3 13.32 1.085 12.98 1.085 12.98 0.3 8.01 0.3 8.01 1.045 7.78 1.045 7.78 0.3 5.635 0.3 5.635 1.075 5.295 1.075 5.295 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.79 0.475 0.79 0.475 2.385 2.545 2.385 2.545 1.625 2.775 1.625 2.775 2.615 0.475 2.615 0.475 3.015 0.245 3.015  ;
        POLYGON 6.585 2.43 6.86 2.43 6.86 1.275 6.75 1.275 6.75 0.99 7.09 0.99 7.09 2.43 8.37 2.43 8.37 1.875 8.6 1.875 8.6 2.66 6.815 2.66 6.815 2.86 6.585 2.86  ;
        POLYGON 3.03 2.705 6.105 2.705 6.105 3.09 7.09 3.09 7.09 2.89 8.6 2.89 8.6 3.12 9.785 3.12 9.785 2.69 10.015 2.69 10.015 3.35 8.37 3.35 8.37 3.12 7.32 3.12 7.32 3.32 5.875 3.32 5.875 2.935 3.03 2.935  ;
        POLYGON 3.27 0.845 4.655 0.845 4.655 1.305 6.035 1.305 6.035 0.53 7.55 0.53 7.55 1.305 8.375 1.305 8.375 0.53 10.07 0.53 10.07 1.14 9.84 1.14 9.84 0.76 8.605 0.76 8.605 1.535 7.32 1.535 7.32 0.76 6.265 0.76 6.265 1.535 4.425 1.535 4.425 1.075 3.27 1.075  ;
        POLYGON 10.855 1.47 10.96 1.47 10.96 0.8 11.19 0.8 11.19 1.47 13.965 1.47 13.965 1.7 11.085 1.7 11.085 2.87 10.855 2.87  ;
        POLYGON 12.2 2.07 14.285 2.07 14.285 0.8 14.555 0.8 14.555 2.87 14.325 2.87 14.325 2.3 12.2 2.3  ;
        POLYGON 9.295 1.82 10.555 1.82 10.555 3.15 12.26 3.15 12.26 2.53 13.9 2.53 13.9 3.16 14.785 3.16 14.785 1.26 15.015 1.26 15.015 3.16 15.905 3.16 15.905 2.07 16.245 2.07 16.245 3.39 13.67 3.39 13.67 2.765 12.49 2.765 12.49 3.39 10.325 3.39 10.325 2.05 9.13 2.05 9.13 2.86 8.9 2.86 8.9 1.82 9.065 1.82 9.065 0.99 9.405 0.99 9.405 1.275 9.295 1.275  ;
        POLYGON 15.425 0.8 15.675 0.8 15.675 1.54 16.885 1.54 16.885 2.315 18.29 2.315 18.29 1.46 18.63 1.46 18.63 2.55 16.655 2.55 16.655 1.775 15.675 1.775 15.675 2.87 15.425 2.87  ;
        POLYGON 17.2 0.995 18.965 0.995 18.965 0.575 19.195 0.575 19.195 1.565 20.245 1.565 20.245 1.275 20.515 1.275 20.515 2.085 20.245 2.085 20.245 1.795 19.195 1.795 19.195 3.345 18.965 3.345 18.965 1.23 17.45 1.23 17.45 2.08 17.2 2.08  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 24.64 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.795 5.18 1.795 5.18 2.215 3.41 2.215  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.6 1.03 0.6 1.03 2.155 0.705 2.155  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.6 2.15 0.6 2.15 2.155 1.825 2.155  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.739 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.465 1.795 6.63 1.795 6.63 2.19 5.465 2.19  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2327 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.76 0.615 21.18 0.615 21.18 1.74 22.98 1.74 22.98 0.615 23.4 0.615 23.4 3.39 22.98 3.39 22.98 2.16 21.18 2.16 21.18 3.39 20.76 3.39  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 2.775 3.62 5.25 3.62 5.25 3.18 5.59 3.18 5.59 3.62 7.57 3.62 7.57 3.35 7.91 3.35 7.91 3.62 10.015 3.62 12.93 3.62 12.93 2.995 13.27 2.995 13.27 3.62 16.245 3.62 17.71 3.62 17.71 2.8 18.05 2.8 18.05 3.62 18.63 3.62 19.785 3.62 19.785 2.46 20.015 2.46 20.015 3.62 20.515 3.62 21.945 3.62 21.945 2.46 22.175 2.46 22.175 3.62 24.115 3.62 24.115 2.46 24.345 2.46 24.345 3.62 24.64 3.62 24.64 4.22 20.515 4.22 18.63 4.22 16.245 4.22 10.015 4.22 2.775 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 24.64 -0.3 24.64 0.3 24.395 0.3 24.395 0.95 24.165 0.95 24.165 0.3 22.155 0.3 22.155 0.95 21.925 0.95 21.925 0.3 19.915 0.3 19.915 0.95 19.685 0.95 19.685 0.3 18.075 0.3 18.075 0.725 17.845 0.725 17.845 0.3 13.32 0.3 13.32 1.085 12.98 1.085 12.98 0.3 8.01 0.3 8.01 1.045 7.78 1.045 7.78 0.3 5.635 0.3 5.635 1.075 5.295 1.075 5.295 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.79 0.475 0.79 0.475 2.385 2.545 2.385 2.545 1.625 2.775 1.625 2.775 2.615 0.475 2.615 0.475 3.015 0.245 3.015  ;
        POLYGON 6.585 2.43 6.86 2.43 6.86 1.275 6.75 1.275 6.75 0.99 7.09 0.99 7.09 2.43 8.37 2.43 8.37 1.875 8.6 1.875 8.6 2.66 6.815 2.66 6.815 2.86 6.585 2.86  ;
        POLYGON 3.03 2.705 6.105 2.705 6.105 3.09 7.09 3.09 7.09 2.89 8.6 2.89 8.6 3.12 9.785 3.12 9.785 2.69 10.015 2.69 10.015 3.35 8.37 3.35 8.37 3.12 7.32 3.12 7.32 3.32 5.875 3.32 5.875 2.935 3.03 2.935  ;
        POLYGON 3.27 0.845 4.655 0.845 4.655 1.305 6.03 1.305 6.03 0.53 7.55 0.53 7.55 1.305 8.375 1.305 8.375 0.53 10.07 0.53 10.07 1.14 9.84 1.14 9.84 0.76 8.605 0.76 8.605 1.535 7.32 1.535 7.32 0.76 6.26 0.76 6.26 1.535 4.425 1.535 4.425 1.075 3.27 1.075  ;
        POLYGON 10.855 1.47 10.96 1.47 10.96 0.8 11.19 0.8 11.19 1.47 13.965 1.47 13.965 1.7 11.085 1.7 11.085 2.87 10.855 2.87  ;
        POLYGON 12.2 2.07 14.285 2.07 14.285 0.8 14.515 0.8 14.515 2.07 14.555 2.07 14.555 2.87 14.325 2.87 14.325 2.3 12.2 2.3  ;
        POLYGON 9.295 1.82 10.555 1.82 10.555 3.15 12.26 3.15 12.26 2.53 13.9 2.53 13.9 3.16 14.785 3.16 14.785 1.26 15.015 1.26 15.015 3.16 15.905 3.16 15.905 2.07 16.245 2.07 16.245 3.39 13.67 3.39 13.67 2.765 12.49 2.765 12.49 3.39 10.325 3.39 10.325 2.05 9.13 2.05 9.13 2.86 8.9 2.86 8.9 1.82 9.065 1.82 9.065 0.99 9.405 0.99 9.405 1.275 9.295 1.275  ;
        POLYGON 15.425 0.8 15.675 0.8 15.675 1.54 16.885 1.54 16.885 2.315 18.29 2.315 18.29 1.46 18.63 1.46 18.63 2.55 16.655 2.55 16.655 1.775 15.675 1.775 15.675 2.87 15.425 2.87  ;
        POLYGON 17.195 0.995 18.965 0.995 18.965 0.575 19.195 0.575 19.195 1.565 20.245 1.565 20.245 1.275 20.515 1.275 20.515 2.085 20.245 2.085 20.245 1.795 19.195 1.795 19.195 3.345 18.965 3.345 18.965 1.23 17.455 1.23 17.455 2.08 17.195 2.08  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 24.08 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.095 1.765 4.39 1.765 4.39 2.19 3.095 2.19  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.155 1.21 20.04 1.21 20.04 0.645 20.67 0.645 20.67 1.02 20.41 1.02 20.41 1.635 19.155 1.635  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.765 6.63 1.765 6.63 2.155 5.13 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.891 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.59 0.555 23.95 0.555 23.95 3.38 23.59 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 10.125 3.62 10.62 3.62 13.12 3.62 13.12 3 13.46 3 13.46 3.62 14.645 3.62 15.135 3.62 15.135 2.665 15.365 2.665 15.365 3.62 16.385 3.62 19.48 3.62 19.48 2.845 19.82 2.845 19.82 3.62 21.345 3.62 21.675 3.62 21.675 2.675 21.905 2.675 21.905 3.62 22.535 3.62 22.535 2.36 22.765 2.36 22.765 3.62 23.24 3.62 24.08 3.62 24.08 4.22 23.24 4.22 21.345 4.22 16.385 4.22 14.645 4.22 10.62 4.22 10.125 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 24.08 -0.3 24.08 0.3 22.715 0.3 22.715 0.925 22.485 0.925 22.485 0.3 19.7 0.3 19.7 0.915 19.36 0.915 19.36 0.3 14.71 0.3 14.71 0.915 14.37 0.915 14.37 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.75 4.63 1.75 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.275 6.835 1.275 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.23 2.745 4.845 2.745 4.845 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.895 3.16 9.895 2.645 10.125 2.645 10.125 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 5.075 2.655 5.075 2.975 3.23 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.375 1.26 6.375 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.97 9.925 0.97 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.605 0.76 6.605 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.62 1.8 10.62 2.035 9.115 2.035 9.115 2.845 8.885 2.845  ;
        POLYGON 11.935 2.53 14.645 2.53 14.645 3.005 14.415 3.005 14.415 2.76 12.165 2.76 12.165 3.005 11.935 3.005  ;
        POLYGON 10.915 2.065 11.045 2.065 11.045 0.63 11.275 0.63 11.275 2.065 11.965 2.065 11.965 1.61 15.37 1.61 15.37 1.84 12.195 1.84 12.195 2.295 11.145 2.295 11.145 3.125 10.915 3.125  ;
        POLYGON 12.46 2.07 15.71 2.07 15.71 0.99 16.05 0.99 16.05 2.07 16.385 2.07 16.385 3.035 16.155 3.035 16.155 2.3 12.46 2.3  ;
        POLYGON 11.505 1.145 14.98 1.145 14.98 0.53 17.845 0.53 17.845 2.06 17.99 2.06 17.99 2.4 17.615 2.4 17.615 0.76 16.6 0.76 16.6 1.735 16.37 1.735 16.37 0.76 15.21 0.76 15.21 1.375 11.735 1.375 11.735 1.72 11.505 1.72  ;
        POLYGON 18.075 0.79 18.305 0.79 18.305 1.51 18.45 1.51 18.45 2.42 18.57 2.42 18.57 2.93 18.22 2.93 18.22 1.745 18.075 1.745  ;
        POLYGON 16.83 0.99 17.385 0.99 17.385 2.69 17.46 2.69 17.46 3.16 18.845 3.16 18.845 2.385 20.425 2.385 20.425 3.155 21.115 3.155 21.115 2.03 21.345 2.03 21.345 3.39 20.195 3.39 20.195 2.615 19.075 2.615 19.075 3.39 17.155 3.39 17.155 1.22 16.83 1.22  ;
        POLYGON 18.68 1.68 18.91 1.68 18.91 1.925 20.655 1.925 20.655 1.56 21.675 1.56 21.675 0.81 21.905 0.81 21.905 1.56 23.24 1.56 23.24 1.79 20.885 1.79 20.885 2.86 20.655 2.86 20.655 2.155 18.68 2.155  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 25.2 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.095 1.765 4.39 1.765 4.39 2.19 3.095 2.19  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.315 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.155 1.21 20.035 1.21 20.035 0.665 20.7 0.665 20.7 1.02 20.41 1.02 20.41 1.635 19.155 1.635  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.765 6.63 1.765 6.63 2.155 5.13 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.11375 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.46 0.6 23.98 0.6 23.98 3.36 23.46 3.36  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 10.125 3.62 10.62 3.62 13.12 3.62 13.12 3 13.46 3 13.46 3.62 14.645 3.62 15.135 3.62 15.135 2.665 15.365 2.665 15.365 3.62 16.385 3.62 19.48 3.62 19.48 2.845 19.82 2.845 19.82 3.62 21.345 3.62 21.675 3.62 21.675 2.57 21.905 2.57 21.905 3.62 22.445 3.62 22.445 2.56 22.675 2.56 22.675 3.62 23.145 3.62 24.535 3.62 24.535 2.56 24.765 2.56 24.765 3.62 25.2 3.62 25.2 4.22 23.145 4.22 21.345 4.22 16.385 4.22 14.645 4.22 10.62 4.22 10.125 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 25.2 -0.3 25.2 0.3 24.865 0.3 24.865 0.925 24.635 0.925 24.635 0.3 22.625 0.3 22.625 0.925 22.395 0.925 22.395 0.3 19.7 0.3 19.7 0.915 19.36 0.915 19.36 0.3 14.71 0.3 14.71 0.915 14.37 0.915 14.37 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.75 4.63 1.75 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.275 6.835 1.275 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.27 2.745 4.845 2.745 4.845 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.895 3.16 9.895 2.645 10.125 2.645 10.125 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 5.075 2.655 5.075 2.975 3.27 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.375 1.26 6.375 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.97 9.925 0.97 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.605 0.76 6.605 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.62 1.8 10.62 2.035 9.115 2.035 9.115 2.845 8.885 2.845  ;
        POLYGON 11.935 2.53 14.645 2.53 14.645 3.005 14.415 3.005 14.415 2.76 12.165 2.76 12.165 3.005 11.935 3.005  ;
        POLYGON 10.915 2.065 11.045 2.065 11.045 0.63 11.275 0.63 11.275 2.065 11.965 2.065 11.965 1.61 15.37 1.61 15.37 1.84 12.195 1.84 12.195 2.295 11.145 2.295 11.145 3.125 10.915 3.125  ;
        POLYGON 12.46 2.07 15.71 2.07 15.71 0.99 16.05 0.99 16.05 2.07 16.385 2.07 16.385 3.035 16.155 3.035 16.155 2.3 12.46 2.3  ;
        POLYGON 11.505 1.145 14.98 1.145 14.98 0.53 17.845 0.53 17.845 2.06 17.99 2.06 17.99 2.4 17.615 2.4 17.615 0.76 16.6 0.76 16.6 1.735 16.37 1.735 16.37 0.76 15.21 0.76 15.21 1.375 11.735 1.375 11.735 1.72 11.505 1.72  ;
        POLYGON 18.075 0.79 18.305 0.79 18.305 1.51 18.45 1.51 18.45 2.42 18.57 2.42 18.57 2.93 18.22 2.93 18.22 1.745 18.075 1.745  ;
        POLYGON 16.83 0.99 17.385 0.99 17.385 2.69 17.46 2.69 17.46 3.16 18.845 3.16 18.845 2.385 20.425 2.385 20.425 3.155 21.115 3.155 21.115 2.03 21.345 2.03 21.345 3.39 20.195 3.39 20.195 2.615 19.075 2.615 19.075 3.39 17.155 3.39 17.155 1.22 16.83 1.22  ;
        POLYGON 18.68 1.68 18.91 1.68 18.91 1.925 20.655 1.925 20.655 1.405 21.675 1.405 21.675 0.81 21.905 0.81 21.905 1.405 23.145 1.405 23.145 2.25 22.915 2.25 22.915 1.635 20.885 1.635 20.885 2.86 20.655 2.86 20.655 2.155 18.68 2.155  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 27.44 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.095 1.765 4.39 1.765 4.39 2.19 3.095 2.19  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.315 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.155 1.17 20.035 1.17 20.035 0.665 20.7 0.665 20.7 1.02 20.41 1.02 20.41 1.635 19.155 1.635  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.09 1.765 6.63 1.765 6.63 2.155 5.09 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2275 ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.46 0.6 23.98 0.6 23.98 1.66 25.7 1.66 25.7 0.6 26.22 0.6 26.22 3.36 25.7 3.36 25.7 2.18 23.98 2.18 23.98 3.36 23.46 3.36  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 10.125 3.62 10.62 3.62 13.12 3.62 13.12 3 13.46 3 13.46 3.62 14.645 3.62 15.135 3.62 15.135 2.665 15.365 2.665 15.365 3.62 16.385 3.62 19.48 3.62 19.48 2.845 19.82 2.845 19.82 3.62 21.345 3.62 21.675 3.62 21.675 2.535 21.905 2.535 21.905 3.62 22.445 3.62 22.445 2.56 22.675 2.56 22.675 3.62 23.145 3.62 24.61 3.62 24.61 2.56 24.84 2.56 24.84 3.62 26.775 3.62 26.775 2.56 27.005 2.56 27.005 3.62 27.44 3.62 27.44 4.22 23.145 4.22 21.345 4.22 16.385 4.22 14.645 4.22 10.62 4.22 10.125 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 27.44 -0.3 27.44 0.3 27.105 0.3 27.105 0.925 26.875 0.925 26.875 0.3 24.865 0.3 24.865 0.925 24.635 0.925 24.635 0.3 22.625 0.3 22.625 0.925 22.395 0.925 22.395 0.3 19.7 0.3 19.7 0.915 19.36 0.915 19.36 0.3 14.71 0.3 14.71 0.915 14.37 0.915 14.37 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.75 4.63 1.75 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.275 6.835 1.275 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.27 2.745 4.845 2.745 4.845 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.895 3.16 9.895 2.645 10.125 2.645 10.125 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 5.075 2.655 5.075 2.975 3.27 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.375 1.26 6.375 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.97 9.925 0.97 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.605 0.76 6.605 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.62 1.8 10.62 2.035 9.115 2.035 9.115 2.845 8.885 2.845  ;
        POLYGON 11.935 2.53 14.645 2.53 14.645 3.005 14.415 3.005 14.415 2.76 12.165 2.76 12.165 3.005 11.935 3.005  ;
        POLYGON 10.915 2.065 11.045 2.065 11.045 0.63 11.275 0.63 11.275 2.065 11.965 2.065 11.965 1.61 15.37 1.61 15.37 1.84 12.195 1.84 12.195 2.295 11.145 2.295 11.145 3.125 10.915 3.125  ;
        POLYGON 12.46 2.07 15.71 2.07 15.71 0.99 16.05 0.99 16.05 2.07 16.385 2.07 16.385 3.035 16.155 3.035 16.155 2.3 12.46 2.3  ;
        POLYGON 11.505 1.145 14.98 1.145 14.98 0.53 17.845 0.53 17.845 2.06 17.99 2.06 17.99 2.4 17.615 2.4 17.615 0.76 16.6 0.76 16.6 1.735 16.37 1.735 16.37 0.76 15.21 0.76 15.21 1.375 11.735 1.375 11.735 1.72 11.505 1.72  ;
        POLYGON 18.075 0.79 18.305 0.79 18.305 1.51 18.45 1.51 18.45 2.42 18.57 2.42 18.57 2.93 18.22 2.93 18.22 1.745 18.075 1.745  ;
        POLYGON 16.83 0.99 17.385 0.99 17.385 2.69 17.46 2.69 17.46 3.16 18.845 3.16 18.845 2.385 20.425 2.385 20.425 3.155 21.115 3.155 21.115 2.03 21.345 2.03 21.345 3.39 20.195 3.39 20.195 2.615 19.075 2.615 19.075 3.39 17.155 3.39 17.155 1.22 16.83 1.22  ;
        POLYGON 18.68 1.68 18.91 1.68 18.91 1.925 20.655 1.925 20.655 1.405 21.675 1.405 21.675 0.81 21.905 0.81 21.905 1.405 23.145 1.405 23.145 2.25 22.915 2.25 22.915 1.635 20.885 1.635 20.885 2.86 20.655 2.86 20.655 2.155 18.68 2.155  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 26.88 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.405 1.765 4.39 1.765 4.39 2.19 3.405 2.19  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.2045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 22.525 1.765 23.43 1.765 23.43 2.155 22.525 2.155  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.605 1.21 21.14 1.21 21.14 2.195 20.605 2.195  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.765 6.63 1.765 6.63 2.155 5.13 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 25.86 2.205 26.255 2.205 26.255 1.16 25.755 1.16 25.755 0.655 26.555 0.655 26.555 2.505 26.32 2.505 26.32 3.38 25.86 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 9.835 3.62 10.405 3.62 13.01 3.62 13.01 3.445 13.35 3.445 13.35 3.62 16.2 3.62 16.2 3.445 16.56 3.445 16.56 3.62 18.275 3.62 20.465 3.62 20.465 2.915 20.695 2.915 20.695 3.62 22.63 3.62 22.63 2.97 22.97 2.97 22.97 3.62 24.49 3.62 25.055 3.62 25.055 2.53 25.285 2.53 25.285 3.62 25.78 3.62 26.88 3.62 26.88 4.22 25.78 4.22 24.49 4.22 18.275 4.22 10.405 4.22 9.835 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 26.88 -0.3 26.88 0.3 25.285 0.3 25.285 1.16 25.055 1.16 25.055 0.3 22.2 0.3 22.2 1.075 21.86 1.075 21.86 0.3 14.14 0.3 14.14 0.915 13.78 0.915 13.78 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.75 4.63 1.75 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.275 6.835 1.275 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.27 2.745 4.845 2.745 4.845 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.605 3.16 9.605 2.485 9.835 2.485 9.835 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 5.075 2.655 5.075 2.975 3.27 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.01 1.26 6.01 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.98 9.925 0.98 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.24 0.76 6.24 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.405 1.8 10.405 2.035 9.115 2.035 9.115 2.845 8.885 2.845  ;
        POLYGON 11.68 2.525 14.6 2.525 14.6 2.78 14.16 2.78 14.16 2.755 12.2 2.755 12.2 2.775 11.68 2.775  ;
        POLYGON 10.8 2.065 11.045 2.065 11.045 0.62 11.275 0.62 11.275 2.065 15.905 2.065 15.905 2.295 11.03 2.295 11.03 2.87 10.8 2.87  ;
        POLYGON 14.96 2.525 16.325 2.525 16.325 1.835 12.295 1.835 12.295 1.605 16.325 1.605 16.325 0.99 16.665 0.99 16.665 2.525 17.79 2.525 17.79 2.78 17.36 2.78 17.36 2.755 15.4 2.755 15.4 2.78 14.96 2.78  ;
        POLYGON 11.265 3.16 12.55 3.16 12.55 2.985 13.81 2.985 13.81 3.16 15.74 3.16 15.74 2.985 17.02 2.985 17.02 3.16 18.045 3.16 18.045 2.035 18.275 2.035 18.275 3.39 16.79 3.39 16.79 3.215 15.97 3.215 15.97 3.39 13.58 3.39 13.58 3.215 12.78 3.215 12.78 3.39 11.265 3.39  ;
        POLYGON 11.625 1.145 14.37 1.145 14.37 0.53 19.675 0.53 19.675 1.765 19.445 1.765 19.445 0.76 17.17 0.76 17.17 1.745 16.94 1.745 16.94 0.76 14.6 0.76 14.6 1.375 11.855 1.375 11.855 1.7 11.625 1.7  ;
        POLYGON 18.57 0.99 19.215 0.99 19.215 1.995 19.955 1.995 19.955 0.715 21.63 0.715 21.63 1.925 21.77 1.925 21.77 2.93 21.43 2.93 21.43 2.155 21.4 2.155 21.4 0.96 20.185 0.96 20.185 2.225 19.775 2.225 19.775 2.835 19.545 2.835 19.545 2.225 18.985 2.225 18.985 1.22 18.57 1.22  ;
        POLYGON 17.445 0.99 17.785 0.99 17.785 1.575 18.755 1.575 18.755 3.16 20.005 3.16 20.005 2.455 21.155 2.455 21.155 3.16 22.08 3.16 22.08 2.51 23.43 2.51 23.43 3.16 24.26 3.16 24.26 2.06 24.49 2.06 24.49 3.39 23.2 3.39 23.2 2.74 22.31 2.74 22.31 3.39 20.925 3.39 20.925 2.685 20.235 2.685 20.235 3.39 18.525 3.39 18.525 1.805 17.445 1.805  ;
        POLYGON 22.065 1.305 24.335 1.305 24.335 0.78 24.565 0.78 24.565 1.6 25.78 1.6 25.78 1.83 24.335 1.83 24.335 1.535 24.03 1.535 24.03 2.93 23.69 2.93 23.69 1.535 22.295 1.535 22.295 2.2 22.065 2.2  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 28 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.765 4.39 1.765 4.39 2.155 3.41 2.155  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.3545 ;
    PORT
      LAYER Metal1 ;
        POLYGON 22.49 1.765 23.43 1.765 23.43 2.155 22.49 2.155  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.605 1.21 21.14 1.21 21.14 2.19 20.605 2.19  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.765 6.63 1.765 6.63 2.155 5.13 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 25.85 2.385 26.79 2.385 27.025 2.385 27.025 1.535 25.85 1.535 25.85 0.61 26.435 0.61 26.435 1.21 27.31 1.21 27.31 2.66 26.79 2.66 26.3 2.66 26.3 3.38 25.85 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 9.835 3.62 10.39 3.62 13.01 3.62 13.01 3.445 13.35 3.445 13.35 3.62 16.2 3.62 16.2 3.445 16.56 3.445 16.56 3.62 18.275 3.62 20.465 3.62 20.465 2.915 20.695 2.915 20.695 3.62 22.63 3.62 22.63 2.97 22.97 2.97 22.97 3.62 24.49 3.62 24.885 3.62 24.885 2.53 25.115 2.53 25.115 3.62 26.79 3.62 27.055 3.62 27.055 2.94 27.285 2.94 27.285 3.62 28 3.62 28 4.22 26.79 4.22 24.49 4.22 18.275 4.22 10.39 4.22 9.835 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 28 -0.3 28 0.3 27.525 0.3 27.525 0.85 27.295 0.85 27.295 0.3 25.285 0.3 25.285 0.85 25.055 0.85 25.055 0.3 22.2 0.3 22.2 1.075 21.86 1.075 21.86 0.3 14.14 0.3 14.14 0.915 13.78 0.915 13.78 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.75 4.63 1.75 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.275 6.835 1.275 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.27 2.745 3.89 2.745 3.89 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.605 3.16 9.605 2.485 9.835 2.485 9.835 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 4.12 2.655 4.12 2.975 3.27 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.01 1.26 6.01 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.98 9.925 0.98 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.24 0.76 6.24 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.39 1.8 10.39 2.035 9.115 2.035 9.115 2.89 8.885 2.89  ;
        POLYGON 11.68 2.525 14.6 2.525 14.6 2.78 14.16 2.78 14.16 2.755 12.2 2.755 12.2 2.775 11.68 2.775  ;
        POLYGON 10.8 2.065 11.045 2.065 11.045 0.62 11.275 0.62 11.275 2.065 15.905 2.065 15.905 2.295 11.03 2.295 11.03 2.87 10.8 2.87  ;
        POLYGON 14.96 2.525 16.325 2.525 16.325 1.835 12.295 1.835 12.295 1.605 16.325 1.605 16.325 0.99 16.665 0.99 16.665 2.525 17.79 2.525 17.79 2.78 17.36 2.78 17.36 2.755 15.4 2.755 15.4 2.78 14.96 2.78  ;
        POLYGON 11.265 3.16 12.55 3.16 12.55 2.985 13.81 2.985 13.81 3.16 15.74 3.16 15.74 2.985 17.02 2.985 17.02 3.16 18.045 3.16 18.045 2.035 18.275 2.035 18.275 3.39 16.79 3.39 16.79 3.215 15.97 3.215 15.97 3.39 13.58 3.39 13.58 3.215 12.78 3.215 12.78 3.39 11.265 3.39  ;
        POLYGON 11.625 1.145 14.37 1.145 14.37 0.53 19.675 0.53 19.675 1.765 19.445 1.765 19.445 0.76 17.17 0.76 17.17 1.745 16.94 1.745 16.94 0.76 14.6 0.76 14.6 1.375 11.855 1.375 11.855 1.7 11.625 1.7  ;
        POLYGON 18.57 0.99 19.215 0.99 19.215 1.995 19.955 1.995 19.955 0.715 21.63 0.715 21.63 1.925 21.77 1.925 21.77 2.93 21.43 2.93 21.43 2.155 21.4 2.155 21.4 0.96 20.185 0.96 20.185 2.225 19.775 2.225 19.775 2.835 19.545 2.835 19.545 2.225 18.985 2.225 18.985 1.22 18.57 1.22  ;
        POLYGON 17.445 0.99 17.785 0.99 17.785 1.575 18.755 1.575 18.755 3.16 20.005 3.16 20.005 2.455 21.155 2.455 21.155 3.16 22.08 3.16 22.08 2.51 23.43 2.51 23.43 3.16 24.26 3.16 24.26 1.91 24.49 1.91 24.49 3.39 23.2 3.39 23.2 2.74 22.315 2.74 22.315 3.39 20.925 3.39 20.925 2.685 20.235 2.685 20.235 3.39 18.525 3.39 18.525 1.805 17.445 1.805  ;
        POLYGON 22.01 1.305 24.335 1.305 24.335 0.64 24.565 0.64 24.565 1.305 25.175 1.305 25.175 1.825 26.79 1.825 26.79 2.095 24.945 2.095 24.945 1.535 24.03 1.535 24.03 2.93 23.69 2.93 23.69 1.535 22.24 1.535 22.24 2.2 22.01 2.2  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 30.24 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.765 4.39 1.765 4.39 2.155 3.41 2.155  ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.3545 ;
    PORT
      LAYER Metal1 ;
        POLYGON 22.49 1.765 23.43 1.765 23.43 2.155 22.49 2.155  ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.605 1.21 21.14 1.21 21.14 2.19 20.605 2.19  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.765 6.63 1.765 6.63 2.155 5.13 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.1216 ;
    PORT
      LAYER Metal1 ;
        POLYGON 25.785 2.385 28.725 2.385 29.255 2.385 29.255 1.535 25.85 1.535 25.85 0.61 26.435 0.61 26.435 1.205 28.135 1.205 28.135 0.61 28.695 0.61 28.695 1.205 29.54 1.205 29.54 2.655 28.725 2.655 28.085 2.655 28.085 3.38 27.585 3.38 27.585 2.655 26.18 2.655 26.18 3.38 25.785 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 9.835 3.62 10.395 3.62 13.01 3.62 13.01 3.445 13.35 3.445 13.35 3.62 16.2 3.62 16.2 3.445 16.56 3.445 16.56 3.62 18.275 3.62 20.465 3.62 20.465 2.915 20.695 2.915 20.695 3.62 22.63 3.62 22.63 2.97 22.97 2.97 22.97 3.62 24.49 3.62 24.765 3.62 24.765 2.53 24.995 2.53 24.995 3.62 26.805 3.62 26.805 3 27.035 3 27.035 3.62 28.725 3.62 28.845 3.62 28.845 3 29.075 3 29.075 3.62 30.24 3.62 30.24 4.22 28.725 4.22 24.49 4.22 18.275 4.22 10.395 4.22 9.835 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 30.24 -0.3 30.24 0.3 29.765 0.3 29.765 0.925 29.535 0.925 29.535 0.3 27.525 0.3 27.525 0.925 27.295 0.925 27.295 0.3 25.285 0.3 25.285 0.925 25.055 0.925 25.055 0.3 22.2 0.3 22.2 1.075 21.86 1.075 21.86 0.3 14.14 0.3 14.14 0.915 13.78 0.915 13.78 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.75 4.63 1.75 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.285 6.835 1.285 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.27 2.745 3.89 2.745 3.89 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.605 3.16 9.605 2.385 9.835 2.385 9.835 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 4.12 2.655 4.12 2.975 3.27 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.01 1.26 6.01 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.98 9.925 0.98 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.24 0.76 6.24 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.395 1.8 10.395 2.035 9.115 2.035 9.115 2.89 8.885 2.89  ;
        POLYGON 11.68 2.525 14.6 2.525 14.6 2.78 14.16 2.78 14.16 2.755 12.2 2.755 12.2 2.775 11.68 2.775  ;
        POLYGON 10.8 2.065 11.045 2.065 11.045 0.62 11.275 0.62 11.275 2.065 15.905 2.065 15.905 2.295 11.03 2.295 11.03 2.87 10.8 2.87  ;
        POLYGON 14.96 2.525 16.325 2.525 16.325 1.835 12.295 1.835 12.295 1.605 16.325 1.605 16.325 0.99 16.665 0.99 16.665 2.525 17.79 2.525 17.79 2.78 17.36 2.78 17.36 2.755 15.4 2.755 15.4 2.78 14.96 2.78  ;
        POLYGON 11.265 3.16 12.55 3.16 12.55 2.985 13.81 2.985 13.81 3.16 15.74 3.16 15.74 2.985 17.02 2.985 17.02 3.16 18.045 3.16 18.045 2.035 18.275 2.035 18.275 3.39 16.79 3.39 16.79 3.215 15.97 3.215 15.97 3.39 13.58 3.39 13.58 3.215 12.78 3.215 12.78 3.39 11.265 3.39  ;
        POLYGON 11.625 1.145 14.37 1.145 14.37 0.53 19.675 0.53 19.675 1.765 19.445 1.765 19.445 0.76 17.17 0.76 17.17 1.745 16.94 1.745 16.94 0.76 14.6 0.76 14.6 1.375 11.855 1.375 11.855 1.7 11.625 1.7  ;
        POLYGON 18.57 0.99 19.215 0.99 19.215 1.995 19.955 1.995 19.955 0.715 21.63 0.715 21.63 1.925 21.77 1.925 21.77 2.93 21.43 2.93 21.43 2.155 21.4 2.155 21.4 0.96 20.185 0.96 20.185 2.225 19.775 2.225 19.775 2.835 19.545 2.835 19.545 2.225 18.985 2.225 18.985 1.22 18.57 1.22  ;
        POLYGON 17.445 0.99 17.785 0.99 17.785 1.575 18.755 1.575 18.755 3.16 20.005 3.16 20.005 2.455 21.155 2.455 21.155 3.16 22.08 3.16 22.08 2.51 23.43 2.51 23.43 3.16 24.26 3.16 24.26 1.91 24.49 1.91 24.49 3.39 23.2 3.39 23.2 2.74 22.315 2.74 22.315 3.39 20.925 3.39 20.925 2.685 20.235 2.685 20.235 3.39 18.525 3.39 18.525 1.805 17.445 1.805  ;
        POLYGON 22.01 1.305 24.335 1.305 24.335 0.655 24.565 0.655 24.565 1.305 25.175 1.305 25.175 1.825 28.725 1.825 28.725 2.095 24.945 2.095 24.945 1.535 24.03 1.535 24.03 2.93 23.69 2.93 23.69 1.535 22.24 1.535 22.24 2.2 22.01 2.2  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffrsnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 25.2 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.765 4.39 1.765 4.39 2.155 3.41 2.155  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.62 1.17 20.11 1.17 20.11 2.19 19.62 2.19  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.765 6.63 1.765 6.63 2.155 5.13 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.8976 ;
    PORT
      LAYER Metal1 ;
        POLYGON 24.22 0.595 24.77 0.595 24.77 3.38 24.22 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 9.835 3.62 10.39 3.62 13.19 3.62 13.19 3.445 13.53 3.445 13.53 3.62 15.46 3.62 15.46 2.91 15.82 2.91 15.82 3.62 17.25 3.62 19.47 3.62 19.47 2.965 19.81 2.965 19.81 3.62 21.59 3.62 21.59 2.965 21.93 2.965 21.93 3.62 22.53 3.62 23.515 3.62 23.515 2.53 23.745 2.53 23.745 3.62 23.99 3.62 25.2 3.62 25.2 4.22 23.99 4.22 22.53 4.22 17.25 4.22 10.39 4.22 9.835 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 25.2 -0.3 25.2 0.3 23.545 0.3 23.545 0.905 23.315 0.905 23.315 0.3 21.705 0.3 21.705 0.89 21.475 0.89 21.475 0.3 13.48 0.3 13.48 0.915 13.12 0.915 13.12 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.74 4.63 1.74 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.275 6.835 1.275 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.27 2.745 3.89 2.745 3.89 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.605 3.16 9.605 2.485 9.835 2.485 9.835 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 4.12 2.655 4.12 2.975 3.27 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.01 1.26 6.01 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.98 9.925 0.98 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.24 0.76 6.24 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.39 1.8 10.39 2.035 9.115 2.035 9.115 2.89 8.885 2.89  ;
        POLYGON 10.8 2.065 11.045 2.065 11.045 0.62 11.275 0.62 11.275 2.065 14.255 2.065 14.255 2.295 11.03 2.295 11.03 2.87 10.8 2.87  ;
        POLYGON 12.475 1.605 14.715 1.605 14.715 1.99 15.47 1.99 15.47 0.99 15.81 0.99 15.81 1.99 16.74 1.99 16.74 2.885 16.51 2.885 16.51 2.22 14.715 2.22 14.715 2.93 14.485 2.93 14.485 1.835 12.475 1.835  ;
        POLYGON 11.265 3.16 12.55 3.16 12.55 2.985 13.99 2.985 13.99 3.16 15 3.16 15 2.45 16.28 2.45 16.28 3.115 17.02 3.115 17.02 2.065 17.25 2.065 17.25 3.345 16.05 3.345 16.05 2.68 15.23 2.68 15.23 3.39 13.76 3.39 13.76 3.215 12.78 3.215 12.78 3.39 11.265 3.39  ;
        POLYGON 11.625 1.145 14.1 1.145 14.1 0.53 18.82 0.53 18.82 1.815 18.45 1.815 18.45 0.76 16.32 0.76 16.32 1.74 16.09 1.74 16.09 0.76 14.33 0.76 14.33 1.375 11.955 1.375 11.955 1.7 11.625 1.7  ;
        POLYGON 17.71 0.99 18.22 0.99 18.22 2.045 19.05 2.045 19.05 0.53 20.84 0.53 20.84 2.93 20.5 2.93 20.5 0.76 19.28 0.76 19.28 2.275 18.78 2.275 18.78 2.885 18.55 2.885 18.55 2.315 17.99 2.315 17.99 1.265 17.71 1.265  ;
        POLYGON 16.59 0.99 16.93 0.99 16.93 1.525 17.76 1.525 17.76 3.115 19.01 3.115 19.01 2.505 20.27 2.505 20.27 3.16 21.11 3.16 21.11 2.505 22.19 2.505 22.19 1.96 22.53 1.96 22.53 2.735 21.34 2.735 21.34 3.39 20.04 3.39 20.04 2.735 19.24 2.735 19.24 3.345 17.53 3.345 17.53 1.76 16.59 1.76  ;
        POLYGON 21.115 1.495 22.54 1.495 22.54 0.655 22.89 0.655 22.89 1.44 23.99 1.44 23.99 1.78 23.005 1.78 23.005 3.15 22.775 3.15 22.775 1.725 21.345 1.725 21.345 2.17 21.115 2.17  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffsnq_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 26.32 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.765 4.39 1.765 4.39 2.155 3.41 2.155  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.062 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.057 ;
    PORT
      LAYER Metal1 ;
        POLYGON 19.62 1.17 20.11 1.17 20.11 2.19 19.62 2.19  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.531 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.7415 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.13 1.765 6.63 1.765 6.63 2.155 5.13 2.155  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0791 ;
    PORT
      LAYER Metal1 ;
        POLYGON 24.555 2.38 25.3 2.38 25.53 2.38 25.53 1.535 24.17 1.535 24.17 0.61 24.695 0.61 24.695 1.265 25.795 1.265 25.795 2.655 25.3 2.655 25.1 2.655 25.1 3.38 24.555 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.375 3.62 5.375 2.885 5.605 2.885 5.605 3.62 7.59 3.62 7.59 3.35 7.93 3.35 7.93 3.62 9.835 3.62 10.39 3.62 13.19 3.62 13.19 3.445 13.53 3.445 13.53 3.62 15.46 3.62 15.46 2.91 15.82 2.91 15.82 3.62 17.25 3.62 19.485 3.62 19.485 2.965 19.825 2.965 19.825 3.62 21.58 3.62 21.58 2.965 21.92 2.965 21.92 3.62 22.54 3.62 23.54 3.62 23.54 2.53 23.77 2.53 23.77 3.62 25.3 3.62 25.595 3.62 25.595 2.945 25.825 2.945 25.825 3.62 26.32 3.62 26.32 4.22 25.3 4.22 22.54 4.22 17.25 4.22 10.39 4.22 9.835 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 26.32 -0.3 26.32 0.3 25.825 0.3 25.825 0.905 25.595 0.905 25.595 0.3 23.545 0.3 23.545 0.905 23.315 0.905 23.315 0.3 21.705 0.3 21.705 0.89 21.475 0.89 21.475 0.3 13.48 0.3 13.48 0.915 13.12 0.915 13.12 0.3 8.095 0.3 8.095 1.045 7.865 1.045 7.865 0.3 5.78 0.3 5.78 1.025 5.55 1.025 5.55 0.3 1.595 0.3 1.595 1.14 1.365 1.14 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.625 2.385 2.625 1.305 4.86 1.305 4.86 1.74 4.63 1.74 4.63 1.535 2.855 1.535 2.855 2.615 0.475 2.615 0.475 3.04 0.245 3.04  ;
        POLYGON 6.61 2.385 6.945 2.385 6.945 1.275 6.835 1.275 6.835 0.99 7.175 0.99 7.175 2.385 8.305 2.385 8.305 1.91 8.535 1.91 8.535 2.62 6.84 2.62 6.84 2.89 6.61 2.89  ;
        POLYGON 3.27 2.745 3.89 2.745 3.89 2.42 6.315 2.42 6.315 3.16 7.13 3.16 7.13 2.89 8.435 2.89 8.435 3.16 9.605 3.16 9.605 2.485 9.835 2.485 9.835 3.39 8.205 3.39 8.205 3.12 7.36 3.12 7.36 3.39 6.085 3.39 6.085 2.655 4.12 2.655 4.12 2.975 3.27 2.975  ;
        POLYGON 3.25 0.845 5.32 0.845 5.32 1.26 6.01 1.26 6.01 0.53 7.635 0.53 7.635 1.295 8.45 1.295 8.45 0.53 10.155 0.53 10.155 0.98 9.925 0.98 9.925 0.76 8.68 0.76 8.68 1.53 7.405 1.53 7.405 0.76 6.24 0.76 6.24 1.49 5.09 1.49 5.09 1.075 3.25 1.075  ;
        POLYGON 8.885 1.8 9.15 1.8 9.15 0.99 9.49 0.99 9.49 1.8 10.39 1.8 10.39 2.035 9.115 2.035 9.115 2.89 8.885 2.89  ;
        POLYGON 10.8 2.065 11.045 2.065 11.045 0.62 11.275 0.62 11.275 2.065 14.255 2.065 14.255 2.295 11.03 2.295 11.03 2.87 10.8 2.87  ;
        POLYGON 12.475 1.605 14.715 1.605 14.715 1.99 15.47 1.99 15.47 0.99 15.81 0.99 15.81 1.99 16.74 1.99 16.74 2.885 16.51 2.885 16.51 2.22 14.715 2.22 14.715 2.93 14.485 2.93 14.485 1.835 12.475 1.835  ;
        POLYGON 11.265 3.16 12.55 3.16 12.55 2.985 13.99 2.985 13.99 3.16 15 3.16 15 2.45 16.28 2.45 16.28 3.115 17.02 3.115 17.02 2.065 17.25 2.065 17.25 3.345 16.05 3.345 16.05 2.68 15.23 2.68 15.23 3.39 13.76 3.39 13.76 3.215 12.78 3.215 12.78 3.39 11.265 3.39  ;
        POLYGON 11.625 1.145 14.1 1.145 14.1 0.53 18.82 0.53 18.82 1.815 18.45 1.815 18.45 0.76 16.32 0.76 16.32 1.74 16.09 1.74 16.09 0.76 14.33 0.76 14.33 1.375 11.855 1.375 11.855 1.7 11.625 1.7  ;
        POLYGON 17.71 0.99 18.22 0.99 18.22 2.045 19.05 2.045 19.05 0.53 20.865 0.53 20.865 2.93 20.525 2.93 20.525 0.76 19.28 0.76 19.28 2.275 18.78 2.275 18.78 2.885 18.55 2.885 18.55 2.315 17.99 2.315 17.99 1.265 17.71 1.265  ;
        POLYGON 16.59 0.99 16.93 0.99 16.93 1.525 17.76 1.525 17.76 3.115 19.01 3.115 19.01 2.505 20.285 2.505 20.285 3.16 21.1 3.16 21.1 2.505 22.2 2.505 22.2 1.96 22.54 1.96 22.54 2.735 21.33 2.735 21.33 3.39 20.055 3.39 20.055 2.735 19.24 2.735 19.24 3.345 17.53 3.345 17.53 1.76 16.59 1.76  ;
        POLYGON 21.115 1.495 22.595 1.495 22.595 0.655 23.03 0.655 23.03 1.825 25.3 1.825 25.3 2.095 23.03 2.095 23.03 3.38 22.8 3.38 22.8 1.725 21.345 1.725 21.345 2.17 21.115 2.17  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffsnq_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 29.68 BY 3.92 ;
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 1.77 4.43 1.77 4.43 2.15 3.41 2.15  ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.816 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.595 1.03 0.595 1.03 2.15 0.705 2.15  ;
    END
  END SE
  PIN SETN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.0805 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.075 1.21 21.23 1.21 21.23 1.59 20.075 1.59  ;
    END
  END SETN
  PIN SI
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.408 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 0.595 2.15 0.595 2.15 2.15 1.825 2.15  ;
    END
  END SI
  PIN CLK
    DIRECTION INPUT ;
    USE clock ;
    ANTENNAGATEAREA 0.6865 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.21 1.77 7.79 1.77 7.79 2.15 6.21 2.15  ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.3055 ;
    PORT
      LAYER Metal1 ;
        POLYGON 25.31 2.055 27.105 2.055 27.44 2.055 27.44 1.345 25.31 1.345 25.31 0.805 25.54 0.805 25.54 1.115 27.44 1.115 27.44 0.595 27.91 0.595 27.91 3.38 27.44 3.38 27.44 2.29 27.105 2.29 25.64 2.29 25.64 3.38 25.31 3.38  ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 1.26 3.62 1.26 2.845 1.6 2.845 1.6 3.62 5.25 3.62 5.25 3.305 5.59 3.305 5.59 3.62 8.1 3.62 8.1 3.35 8.44 3.35 8.44 3.62 10.85 3.62 11.29 3.62 13.51 3.62 13.51 3.36 13.85 3.36 13.85 3.62 15.985 3.62 15.985 2.93 16.215 2.93 16.215 3.62 17.99 3.62 19.93 3.62 19.93 2.66 20.27 2.66 20.27 3.62 21.235 3.62 22.285 3.62 22.285 2.53 22.515 2.53 22.515 3.62 24.325 3.62 24.325 2.53 24.555 2.53 24.555 3.62 26.38 3.62 26.38 2.53 26.61 2.53 26.61 3.62 27.105 3.62 28.57 3.62 28.57 2.53 28.8 2.53 28.8 3.62 29.68 3.62 29.68 4.22 27.105 4.22 21.235 4.22 17.99 4.22 11.29 4.22 10.85 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 29.68 -0.3 29.68 0.3 28.9 0.3 28.9 1.145 28.67 1.145 28.67 0.3 26.715 0.3 26.715 0.75 26.375 0.75 26.375 0.3 24.42 0.3 24.42 1.145 24.19 1.145 24.19 0.3 22.18 0.3 22.18 1.02 21.95 1.02 21.95 0.3 14.19 0.3 14.19 0.915 13.85 0.915 13.85 0.3 8.41 0.3 8.41 0.475 8.07 0.475 8.07 0.3 5.79 0.3 5.79 0.475 5.45 0.475 5.45 0.3 1.595 0.3 1.595 1.16 1.365 1.16 1.365 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.245 0.78 0.475 0.78 0.475 2.385 2.6 2.385 2.6 2.105 2.83 2.105 2.83 2.385 4.725 2.385 4.725 1.455 5.065 1.455 5.065 2.615 0.475 2.615 0.475 3.14 0.245 3.14  ;
        POLYGON 6.785 2.43 8.815 2.43 8.815 1.395 6.51 1.395 6.51 0.99 6.85 0.99 6.85 1.165 9.045 1.165 9.045 2.66 7.07 2.66 7.07 2.835 6.785 2.835  ;
        POLYGON 3.27 2.845 6.05 2.845 6.05 3.16 7.56 3.16 7.56 2.89 9.095 2.89 9.095 3.065 10.51 3.065 10.51 2.655 10.85 2.655 10.85 3.295 8.865 3.295 8.865 3.12 7.79 3.12 7.79 3.39 5.82 3.39 5.82 3.075 3.27 3.075  ;
        POLYGON 3.27 0.705 6.02 0.705 6.02 0.53 7.84 0.53 7.84 0.705 9.085 0.705 9.085 0.53 10.895 0.53 10.895 0.97 10.665 0.97 10.665 0.76 9.315 0.76 9.315 0.935 7.61 0.935 7.61 0.76 6.25 0.76 6.25 0.935 3.61 0.935 3.61 1.095 3.27 1.095  ;
        POLYGON 9.395 2.495 9.71 2.495 9.71 0.99 10.05 0.99 10.05 2.045 11.29 2.045 11.29 2.28 9.995 2.28 9.995 2.835 9.395 2.835  ;
        POLYGON 11.585 1.725 11.785 1.725 11.785 0.68 12.015 0.68 12.015 1.725 14.67 1.725 14.67 1.96 11.815 1.96 11.815 3.015 11.585 3.015  ;
        POLYGON 12.31 1.26 14.745 1.26 14.745 0.53 16.81 0.53 16.81 0.76 14.975 0.76 14.975 1.495 12.31 1.495  ;
        POLYGON 12.85 2.19 14.965 2.19 14.965 1.805 16.03 1.805 16.03 0.99 16.37 0.99 16.37 1.805 17.51 1.805 17.51 2.81 17.17 2.81 17.17 2.04 15.25 2.04 15.25 2.78 14.91 2.78 14.91 2.425 12.85 2.425  ;
        POLYGON 12.11 2.9 14.55 2.9 14.55 3.16 15.48 3.16 15.48 2.465 16.93 2.465 16.93 3.04 17.99 3.04 17.99 3.31 16.7 3.31 16.7 2.7 15.71 2.7 15.71 3.39 14.32 3.39 14.32 3.13 12.45 3.13 12.45 3.355 12.11 3.355  ;
        POLYGON 19.495 2.2 21.235 2.2 21.235 2.835 21.005 2.835 21.005 2.43 19.495 2.43 19.495 2.89 19.265 2.89 19.265 1.22 18.27 1.22 18.27 0.99 19.77 0.99 19.77 1.22 19.495 1.22  ;
        POLYGON 17.15 0.99 17.81 0.99 17.81 0.53 21.72 0.53 21.72 1.45 22.775 1.45 22.775 1.685 21.49 1.685 21.49 0.76 18.04 0.76 18.04 1.875 18.475 1.875 18.475 2.89 18.245 2.89 18.245 2.105 17.81 2.105 17.81 1.22 17.15 1.22  ;
        POLYGON 21.53 1.965 23.07 1.965 23.07 0.805 23.3 0.805 23.3 1.575 27.105 1.575 27.105 1.805 23.535 1.805 23.535 3.38 23.305 3.38 23.305 2.195 21.53 2.195  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__sdffsnq_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__tieh
  CLASS core TIEHIGH ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__tieh 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 2.24 BY 3.92 ;
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.5368 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.22 2.305 1.58 2.305 1.58 3.39 1.22 3.39  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.25 3.62 0.25 2.36 0.48 2.36 0.48 3.62 1.6 3.62 2.24 3.62 2.24 4.22 1.6 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 2.24 -0.3 2.24 0.3 0.48 0.3 0.48 1.16 0.25 1.16 0.25 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.875 1.335 1.37 1.335 1.37 0.53 1.6 0.53 1.6 1.57 0.875 1.57  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__tieh

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__tiel
  CLASS core TIELOW ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__tiel 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 2.24 BY 3.92 ;
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.3608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.22 0.53 1.595 0.53 1.595 1.65 1.22 1.65  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.345 3.62 0.345 2.345 0.575 2.345 0.575 3.62 1.595 3.62 2.24 3.62 2.24 4.22 1.595 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 2.24 -0.3 2.24 0.3 0.475 0.3 0.475 1.16 0.245 1.16 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.87 1.95 1.595 1.95 1.595 3.39 1.365 3.39 1.365 2.185 0.87 2.185  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__tiel

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xnor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 7.28 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.815 1.45 2.22 1.45 2.22 1.825 3.445 1.825 4.57 1.825 4.57 2.095 3.445 2.095 1.815 2.095  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.91 1.625 1.535 1.625 1.535 2.385 3.445 2.385 5.185 2.385 5.185 1.51 6.01 1.51 6.01 1.74 5.455 1.74 5.455 2.655 3.445 2.655 1.305 2.655 1.305 1.855 0.91 1.855  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.45635 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.305 2.945 3.445 2.945 5.745 2.945 5.745 1.98 6.29 1.98 6.29 1.22 4.98 1.22 4.98 0.99 6.58 0.99 6.58 2.215 6.02 2.215 6.02 3.215 3.445 3.215 3.305 3.215  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.385 3.62 0.385 2.72 0.615 2.72 0.615 3.62 2.65 3.62 2.65 2.93 2.99 2.93 2.99 3.62 3.445 3.62 6.305 3.62 6.305 2.69 6.535 2.69 6.535 3.62 6.69 3.62 7.28 3.62 7.28 4.22 6.69 4.22 3.445 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 7.28 -0.3 7.28 0.3 2.71 0.3 2.71 0.76 2.37 0.76 2.37 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.33 0.53 0.67 0.53 0.67 0.99 3.445 0.99 3.445 1.565 3.105 1.565 3.105 1.22 0.615 1.22 0.615 2.18 1.075 2.18 1.075 2.945 1.78 2.945 1.78 3.215 0.845 3.215 0.845 2.415 0.33 2.415  ;
        POLYGON 3.63 0.53 6.69 0.53 6.69 0.76 3.63 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor2_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xnor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 9.52 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.6005 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.825 1.57 2.29 1.57 2.29 1.825 3.535 1.825 3.855 1.825 3.855 1.255 4.48 1.255 4.48 1.745 4.105 1.745 4.105 2.095 3.535 2.095 1.825 2.095  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.6005 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.835 1.655 1.535 1.655 1.535 2.325 3.535 2.325 4.29 2.325 4.29 2.235 5.215 2.235 5.215 1.785 5.475 1.785 5.475 2.47 4.52 2.47 4.52 2.66 3.535 2.66 1.26 2.66 1.26 1.885 0.835 1.885  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.1828 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.585 0.6 8.265 0.6 8.265 3.38 7.585 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.435 3.62 2.435 2.915 2.665 2.915 2.665 3.62 3.535 3.62 6.11 3.62 6.545 3.62 6.545 2.53 6.775 2.53 6.775 3.62 7.29 3.62 8.685 3.62 8.685 2.53 8.915 2.53 8.915 3.62 9.52 3.62 9.52 4.22 7.29 4.22 6.11 4.22 3.535 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 9.52 -0.3 9.52 0.3 9.015 0.3 9.015 1.115 8.785 1.115 8.785 0.3 6.775 0.3 6.775 0.915 6.545 0.915 6.545 0.3 6.055 0.3 6.055 0.915 5.825 0.915 5.825 0.3 2.715 0.3 2.715 0.825 2.485 0.825 2.485 0.3 0.475 0.3 0.475 0.825 0.245 0.825 0.245 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 1.055 1.31 1.055 1.31 0.53 1.65 0.53 1.65 1.055 3.27 1.055 3.27 1.365 3.535 1.365 3.535 1.595 3.04 1.595 3.04 1.29 0.575 1.29 0.575 3.36 0.345 3.36  ;
        POLYGON 3.64 3.16 6.11 3.16 6.11 3.39 3.64 3.39  ;
        POLYGON 4.75 2.7 5.705 2.7 5.705 1.555 4.81 1.555 4.81 0.82 3.64 0.82 3.64 0.59 5.04 0.59 5.04 1.155 7.29 1.155 7.29 2.11 6.92 2.11 6.92 1.555 5.935 1.555 5.935 2.93 4.75 2.93  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor2_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xnor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 11.76 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.498 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.58 2.225 1.58 2.225 1.795 3.4 1.795 3.785 1.795 3.785 1.66 4.55 1.66 4.55 2.01 4.06 2.01 4.06 2.12 3.4 2.12 1.83 2.12  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.498 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.755 1.81 1.535 1.81 1.535 2.36 3.4 2.36 4.29 2.36 4.29 2.24 4.84 2.24 4.84 1.81 5.63 1.81 5.63 2.1 5.07 2.1 5.07 2.47 4.52 2.47 4.52 2.68 3.4 2.68 1.26 2.68 1.26 2.095 0.755 2.095  ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2436 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.61 2.36 10.5 2.36 10.775 2.36 10.775 1.43 7.665 1.43 7.665 0.53 7.895 0.53 7.895 1.195 9.905 1.195 9.905 0.53 10.135 0.53 10.135 1.195 11.06 1.195 11.06 2.7 10.5 2.7 10.14 2.7 10.14 3.38 9.8 3.38 9.8 2.7 7.95 2.7 7.95 3.38 7.61 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.665 3.62 2.665 2.94 2.895 2.94 2.895 3.62 3.4 3.62 6.11 3.62 6.645 3.62 6.645 2.53 6.875 2.53 6.875 3.62 8.735 3.62 8.735 3.015 8.965 3.015 8.965 3.62 10.5 3.62 10.925 3.62 10.925 3.015 11.155 3.015 11.155 3.62 11.76 3.62 11.76 4.22 10.5 4.22 6.11 4.22 3.4 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 11.76 -0.3 11.76 0.3 11.255 0.3 11.255 0.915 11.025 0.915 11.025 0.3 9.015 0.3 9.015 0.915 8.785 0.915 8.785 0.3 6.775 0.3 6.775 0.915 6.545 0.915 6.545 0.3 6.055 0.3 6.055 0.915 5.825 0.915 5.825 0.3 2.77 0.3 2.77 0.76 2.43 0.76 2.43 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.23 0.99 1.31 0.99 1.31 0.53 1.65 0.53 1.65 0.99 3.4 0.99 3.4 1.555 3 1.555 3 1.225 0.525 1.225 0.525 2.72 0.23 2.72  ;
        POLYGON 3.575 3.16 6.11 3.16 6.11 3.39 3.575 3.39  ;
        POLYGON 4.75 2.7 6.01 2.7 6.01 1.43 3.785 1.43 3.785 0.53 4.015 0.53 4.015 1.195 6.24 1.195 6.24 1.665 10.5 1.665 10.5 1.895 6.24 1.895 6.24 2.93 4.75 2.93  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor2_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xnor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 13.44 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.77 1.455 2.225 1.455 2.225 1.825 3.495 1.825 3.67 1.825 3.67 1.455 4.77 1.455 4.77 1.69 3.9 1.69 3.9 2.095 3.495 2.095 1.77 2.095  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.87 2.385 3.495 2.385 4.13 2.385 4.13 1.92 5.175 1.92 5.175 1.595 5.62 1.595 5.62 2.15 4.36 2.15 4.36 2.655 3.495 2.655 0.87 2.655  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.085 1.825 9.54 1.825 10.765 1.825 10.765 2.095 9.54 2.095 8.085 2.095  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.5111 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.57 2.92 11.88 2.92 11.88 2.36 12.17 2.36 12.44 2.36 12.44 1.58 11.17 1.58 11.17 0.99 12.76 0.99 12.76 2.68 12.215 2.68 12.215 3.24 12.17 3.24 9.57 3.24  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.37 3.62 2.37 2.9 2.73 2.9 2.73 3.62 3.495 3.62 6.12 3.62 6.545 3.62 6.545 2.84 6.775 2.84 6.775 3.62 8.76 3.62 8.76 2.815 9.1 2.815 9.1 3.62 12.17 3.62 12.465 3.62 12.465 3.015 12.695 3.015 12.695 3.62 12.86 3.62 13.44 3.62 13.44 4.22 12.86 4.22 12.17 4.22 6.12 4.22 3.495 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 13.44 -0.3 13.44 0.3 8.87 0.3 8.87 0.76 8.53 0.76 8.53 0.3 6.11 0.3 6.11 0.76 5.77 0.76 5.77 0.3 2.77 0.3 2.77 0.76 2.43 0.76 2.43 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 0.99 1.305 0.99 1.305 0.53 1.65 0.53 1.65 0.99 3.495 0.99 3.495 1.22 0.575 1.22 0.575 3.195 0.345 3.195  ;
        POLYGON 3.72 2.9 4.08 2.9 4.08 3.16 5.76 3.16 5.76 2.9 6.12 2.9 6.12 3.39 3.72 3.39  ;
        POLYGON 6.49 0.53 6.83 0.53 6.83 0.99 9.54 0.99 9.54 1.565 9.2 1.565 9.2 1.225 7.85 1.225 7.85 2.93 7.51 2.93 7.51 1.225 6.49 1.225  ;
        POLYGON 4.74 2.38 5.88 2.38 5.88 1.225 3.73 1.225 3.73 0.53 4.07 0.53 4.07 0.99 6.11 0.99 6.11 2.38 7.03 2.38 7.03 1.535 7.26 1.535 7.26 3.16 8.27 3.16 8.27 2.33 11.22 2.33 11.22 1.86 12.17 1.86 12.17 2.095 11.45 2.095 11.45 2.565 8.5 2.565 8.5 3.39 7.03 3.39 7.03 2.61 5.1 2.61 5.1 2.93 4.74 2.93  ;
        POLYGON 9.74 0.53 12.86 0.53 12.86 0.76 9.74 0.76  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor3_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xnor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 15.68 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.935 1.265 4.905 1.265 4.905 1.535 1.935 1.535  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.9045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 2.385 3.57 2.385 3.935 2.385 3.935 1.815 5.715 1.815 5.715 2.1 4.24 2.1 4.24 2.655 3.57 2.655 0.825 2.655  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.598 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.3 1.815 9.905 1.815 10.17 1.815 10.17 1.21 11.075 1.21 11.075 1.61 10.425 1.61 10.425 2.095 9.905 2.095 8.3 2.095  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7952 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.015 2.36 14.915 2.36 15.155 2.36 15.155 1.56 12.965 1.56 12.965 0.6 13.31 0.6 13.31 1.24 15.155 1.24 15.155 0.6 15.535 0.6 15.535 3.39 15.155 3.39 15.155 2.68 14.915 2.68 13.295 2.68 13.295 3.39 13.015 3.39  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.42 3.62 2.42 2.895 2.78 2.895 2.78 3.62 3.57 3.62 6.055 3.62 9.09 3.62 9.09 2.785 9.43 2.785 9.43 3.62 12.575 3.62 14.035 3.62 14.035 2.95 14.265 2.95 14.265 3.62 14.915 3.62 15.68 3.62 15.68 4.22 14.915 4.22 12.575 4.22 6.055 4.22 3.57 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 15.68 -0.3 15.68 0.3 14.315 0.3 14.315 0.975 14.085 0.975 14.085 0.3 12.49 0.3 12.49 0.635 12.15 0.635 12.15 0.3 9.275 0.3 9.275 0.89 9.045 0.89 9.045 0.3 6.91 0.3 6.91 0.76 6.57 0.76 6.57 0.3 6.11 0.3 6.11 0.76 5.77 0.76 5.77 0.3 2.855 0.3 2.855 0.76 2.515 0.76 2.515 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 0.99 1.31 0.99 1.31 0.53 1.65 0.53 1.65 1.765 3.57 1.765 3.57 1.995 1.365 1.995 1.365 1.225 0.575 1.225 0.575 3.19 0.345 3.19  ;
        POLYGON 3.72 2.895 4.08 2.895 4.08 3.155 5.76 3.155 5.76 2.84 6.055 2.84 6.055 3.39 3.72 3.39  ;
        POLYGON 6.745 1.86 7.69 1.86 7.69 0.53 8.03 0.53 8.03 1.15 9.905 1.15 9.905 1.555 9.515 1.555 9.515 1.38 8.03 1.38 8.03 2.095 7.085 2.095 7.085 2.925 6.745 2.925  ;
        POLYGON 6.515 3.155 7.835 3.155 7.835 2.325 10.655 2.325 10.655 2.24 11.765 2.24 11.765 1.715 11.995 1.715 11.995 2.47 10.885 2.47 10.885 2.555 8.065 2.555 8.065 3.39 6.285 3.39 6.285 2.565 5.09 2.565 5.09 2.925 4.75 2.925 4.75 2.335 6.285 2.335 6.285 1.22 5.23 1.22 5.23 0.76 3.73 0.76 3.73 0.53 5.46 0.53 5.46 0.99 7.435 0.99 7.435 1.225 6.515 1.225  ;
        POLYGON 10.045 3.16 12.575 3.16 12.575 3.39 10.045 3.39  ;
        POLYGON 11.115 2.7 12.345 2.7 12.345 1.095 11.405 1.095 11.405 0.765 10.035 0.765 10.035 0.53 11.71 0.53 11.71 0.865 12.575 0.865 12.575 1.815 14.915 1.815 14.915 2.045 12.575 2.045 12.575 2.93 11.115 2.93  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor3_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xnor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xnor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 17.92 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.88 1.24 4.42 1.24 4.42 1.535 1.88 1.535  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.875 1.565 1.105 1.565 1.105 2.265 3.22 2.265 3.45 2.265 3.45 1.82 5.26 1.82 5.26 2.095 3.89 2.095 3.89 2.495 3.22 2.495 0.875 2.495  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5105 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.175 1.8 9.745 1.8 10.02 1.8 10.02 1.255 11.15 1.255 11.15 1.565 10.275 1.565 10.275 2.095 9.745 2.095 8.175 2.095  ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.978 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.94 2.36 17.06 2.36 17.32 2.36 17.32 1.535 12.84 1.535 12.84 0.655 13.07 0.655 13.07 1.26 15.08 1.26 15.08 0.655 15.31 0.655 15.31 1.26 17.32 1.26 17.32 0.6 17.775 0.6 17.775 3.38 17.22 3.38 17.22 2.68 17.06 2.68 15.26 2.68 15.26 3.38 15.03 3.38 15.03 2.68 13.17 2.68 13.17 3.38 12.94 3.38  ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.33 3.62 2.33 2.725 2.67 2.725 2.67 3.62 3.22 3.62 6.165 3.62 8.965 3.62 8.965 2.785 9.305 2.785 9.305 3.62 12.375 3.62 13.96 3.62 13.96 3.015 14.19 3.015 14.19 3.62 16.15 3.62 16.15 3.015 16.38 3.015 16.38 3.62 17.06 3.62 17.92 3.62 17.92 4.22 17.06 4.22 12.375 4.22 6.165 4.22 3.22 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 17.92 -0.3 17.92 0.3 16.43 0.3 16.43 0.905 16.2 0.905 16.2 0.3 14.19 0.3 14.19 0.905 13.96 0.905 13.96 0.3 12.365 0.3 12.365 0.64 12.025 0.64 12.025 0.3 9.145 0.3 9.145 0.84 8.915 0.84 8.915 0.3 6.74 0.3 6.74 0.76 5.59 0.76 5.59 0.3 2.77 0.3 2.77 0.76 2.43 0.76 2.43 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 0.99 1.31 0.99 1.31 0.53 1.65 0.53 1.65 1.765 3.22 1.765 3.22 2.035 1.42 2.035 1.42 1.225 0.575 1.225 0.575 3.015 0.345 3.015  ;
        POLYGON 3.55 2.725 3.89 2.725 3.89 3.16 5.825 3.16 5.825 2.725 6.165 2.725 6.165 3.39 3.55 3.39  ;
        POLYGON 6.905 1.8 7.52 1.8 7.52 0.53 7.86 0.53 7.86 1.075 9.745 1.075 9.745 1.56 9.405 1.56 9.405 1.305 7.86 1.305 7.86 2.095 7.245 2.095 7.245 2.93 6.905 2.93  ;
        POLYGON 6.625 3.16 8.115 3.16 8.115 2.325 10.505 2.325 10.505 1.82 11.76 1.82 11.76 2.18 10.735 2.18 10.735 2.555 8.39 2.555 8.39 3.39 6.395 3.39 6.395 2.495 5.67 2.495 5.67 2.555 4.91 2.555 4.91 2.93 4.57 2.93 4.57 2.325 5.44 2.325 5.44 2.265 6.395 2.265 6.395 1.535 5.115 1.535 5.115 0.76 3.55 0.76 3.55 0.53 5.345 0.53 5.345 1.3 7.275 1.3 7.275 1.535 6.625 1.535  ;
        POLYGON 9.895 3.16 12.375 3.16 12.375 3.39 9.895 3.39  ;
        POLYGON 10.915 2.7 12.145 2.7 12.145 1.485 11.565 1.485 11.565 0.76 9.895 0.76 9.895 0.53 11.795 0.53 11.795 1.255 12.375 1.255 12.375 1.765 17.06 1.765 17.06 1.995 12.375 1.995 12.375 2.93 10.915 2.93  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xnor3_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor2_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor2_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 6.72 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.598 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.875 1.82 3.51 1.82 3.785 1.82 3.785 1.34 4.525 1.34 4.525 1.57 4.015 1.57 4.015 2.1 3.51 2.1 1.875 2.1  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.598 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.88 1.69 1.56 1.69 1.56 2.33 3.51 2.33 4.255 2.33 4.255 1.8 5.49 1.8 5.49 2.155 4.495 2.155 4.495 2.56 3.51 2.56 2.325 2.56 2.325 2.73 0.88 2.73  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.75 2.695 5.72 2.695 5.72 1.11 3.785 1.11 3.785 0.53 4.015 0.53 4.015 0.875 6.04 0.875 6.04 2.925 4.75 2.925  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.71 3.62 2.71 2.79 3.05 2.79 3.05 3.62 3.51 3.62 6.12 3.62 6.72 3.62 6.72 4.22 6.12 4.22 3.51 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 6.72 -0.3 6.72 0.3 6.11 0.3 6.11 0.635 5.77 0.635 5.77 0.3 2.95 0.3 2.95 0.76 2.61 0.76 2.61 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.29 0.99 1.31 0.99 1.31 0.53 1.65 0.53 1.65 0.99 3.51 0.99 3.51 1.555 3.17 1.555 3.17 1.29 0.63 1.29 0.63 3.35 0.29 3.35  ;
        POLYGON 3.59 3.155 6.12 3.155 6.12 3.39 3.59 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor2_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor2_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor2_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 10.08 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.85 1.45 2.87 1.45 2.87 1.795 3.52 1.795 4.27 1.795 4.27 1.265 4.565 1.265 4.565 2.095 3.52 2.095 2.595 2.095 2.595 1.68 1.85 1.68  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.915 1.8 1.61 1.8 1.61 1.91 2.315 1.91 2.315 2.325 3.52 2.325 4.83 2.325 4.83 1.8 6.225 1.8 6.225 2.12 5.105 2.12 5.105 2.68 3.52 2.68 3.375 2.68 3.375 2.555 2.035 2.555 2.035 2.14 0.915 2.14  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.195 2.36 9.08 2.36 9.315 2.36 9.315 1.56 8.195 1.56 8.195 0.61 8.545 0.61 8.545 1.24 9.6 1.24 9.6 2.68 9.08 2.68 8.56 2.68 8.56 3.38 8.195 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.455 3.62 0.455 2.83 0.685 2.83 0.685 3.62 2.72 3.62 2.72 2.79 3.06 2.79 3.06 3.62 3.52 3.62 6.32 3.62 6.32 2.815 6.66 2.815 6.66 3.62 7.295 3.62 7.295 2.53 7.525 2.53 7.525 3.62 9.08 3.62 9.335 3.62 9.335 2.94 9.565 2.94 9.565 3.62 10.08 3.62 10.08 4.22 9.08 4.22 3.52 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 10.08 -0.3 10.08 0.3 9.665 0.3 9.665 0.99 9.435 0.99 9.435 0.3 7.425 0.3 7.425 0.99 7.195 0.99 7.195 0.3 2.96 0.3 2.96 0.76 2.62 0.76 2.62 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.4 0.53 0.74 0.53 0.74 0.99 3.52 0.99 3.52 1.555 3.18 1.555 3.18 1.22 0.68 1.22 0.68 2.37 1.705 2.37 1.705 3.35 1.475 3.35 1.475 2.6 0.4 2.6  ;
        POLYGON 3.65 0.53 6.77 0.53 6.77 0.76 3.65 0.76  ;
        POLYGON 3.6 2.99 5.4 2.99 5.4 2.35 6.54 2.35 6.54 1.22 5.07 1.22 5.07 0.99 6.77 0.99 6.77 1.82 9.08 1.82 9.08 2.095 6.77 2.095 6.77 2.58 5.63 2.58 5.63 3.22 3.6 3.22  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor2_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor2_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor2_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.32 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.448 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.935 1.825 3.51 1.825 4.225 1.825 4.225 1.23 4.525 1.23 4.525 2.095 3.51 2.095 1.935 2.095  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.448 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.86 1.81 1.7 1.81 1.7 2.325 3.51 2.325 4.795 2.325 4.795 1.8 6.18 1.8 6.18 2.12 5.025 2.12 5.025 2.68 3.51 2.68 3 2.68 3 2.555 1.425 2.555 1.425 2.1 0.86 2.1  ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.2436 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.27 2.36 11.275 2.36 11.51 2.36 11.51 1.56 8.27 1.56 8.27 0.655 8.5 0.655 8.5 1.24 10.51 1.24 10.51 0.655 10.74 0.655 10.74 1.24 11.78 1.24 11.78 2.68 11.275 2.68 10.69 2.68 10.69 3.38 10.46 3.38 10.46 2.68 8.5 2.68 8.5 3.38 8.27 3.38  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 0.355 3.62 0.355 2.795 0.695 2.795 0.695 3.62 2.395 3.62 2.395 2.785 2.735 2.785 2.735 3.62 3.51 3.62 6.275 3.62 6.275 2.815 6.615 2.815 6.615 3.62 7.25 3.62 7.25 2.53 7.48 2.53 7.48 3.62 9.34 3.62 9.34 3 9.57 3 9.57 3.62 11.275 3.62 11.53 3.62 11.53 3 11.76 3 11.76 3.62 12.32 3.62 12.32 4.22 11.275 4.22 3.51 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.32 -0.3 12.32 0.3 11.86 0.3 11.86 0.985 11.63 0.985 11.63 0.3 9.62 0.3 9.62 0.985 9.39 0.985 9.39 0.3 7.38 0.3 7.38 0.905 7.15 0.905 7.15 0.3 2.915 0.3 2.915 0.76 2.575 0.76 2.575 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.355 0.53 0.695 0.53 0.695 0.99 3.51 0.99 3.51 1.555 3.17 1.555 3.17 1.22 0.585 1.22 0.585 2.33 1.19 2.33 1.19 2.785 1.805 2.785 1.805 3.015 0.93 3.015 0.93 2.565 0.355 2.565  ;
        POLYGON 3.605 0.53 6.725 0.53 6.725 0.76 3.605 0.76  ;
        POLYGON 3.66 2.965 5.45 2.965 5.45 2.35 6.495 2.35 6.495 1.22 4.92 1.22 4.92 0.99 6.725 0.99 6.725 1.815 11.275 1.815 11.275 2.105 6.725 2.105 6.725 2.585 5.68 2.585 5.68 3.195 3.66 3.195  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor2_4

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor3_1
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor3_1 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 12.88 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8945 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.89 1.265 4.6 1.265 4.6 1.535 1.89 1.535  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8945 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.865 1.57 1.095 1.57 1.095 2.225 3.51 2.225 3.915 2.225 3.915 1.82 5.6 1.82 5.6 2.095 4.195 2.095 4.195 2.455 3.51 2.455 2.1 2.455 2.1 2.71 0.865 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.6005 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.205 1.455 8.545 1.455 8.545 1.825 9.745 1.825 9.975 1.825 9.975 1.265 11.11 1.265 11.11 1.56 10.205 1.56 10.205 2.1 9.745 2.1 8.205 2.1  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.0608 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.77 2.7 11.585 2.7 11.88 2.7 11.88 1.295 11.56 1.295 11.56 1 10.045 1 10.045 0.67 11.83 0.67 11.83 1.015 12.2 1.015 12.2 2.93 11.585 2.93 10.77 2.93  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.33 3.62 2.33 2.685 2.67 2.685 2.67 3.62 3.51 3.62 6.055 3.62 8.75 3.62 8.75 2.79 9.09 2.79 9.09 3.62 12.16 3.62 12.88 3.62 12.88 4.22 12.16 4.22 6.055 4.22 3.51 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 12.88 -0.3 12.88 0.3 12.425 0.3 12.425 0.635 12.085 0.635 12.085 0.3 9.275 0.3 9.275 0.76 8.915 0.76 8.915 0.3 6.85 0.3 6.85 0.76 5.77 0.76 5.77 0.3 2.77 0.3 2.77 0.76 2.43 0.76 2.43 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.345 1.07 1.31 1.07 1.31 0.53 1.65 0.53 1.65 1.765 3.51 1.765 3.51 1.995 1.385 1.995 1.385 1.305 0.575 1.305 0.575 2.98 0.345 2.98  ;
        POLYGON 3.73 2.755 4.07 2.755 4.07 3.16 5.825 3.16 5.825 2.815 6.055 2.815 6.055 3.39 3.73 3.39  ;
        POLYGON 6.745 1.535 7.625 1.535 7.625 0.53 7.965 0.53 7.965 0.99 9.745 0.99 9.745 1.555 9.395 1.555 9.395 1.22 7.93 1.22 7.93 1.765 6.975 1.765 6.975 2.925 6.745 2.925  ;
        POLYGON 6.11 2.325 6.515 2.325 6.515 3.16 7.695 3.16 7.695 2.33 10.395 2.33 10.395 2.24 11.35 2.24 11.35 1.76 11.585 1.76 11.585 2.47 10.585 2.47 10.585 2.56 7.925 2.56 7.925 3.39 6.285 3.39 6.285 2.555 5.09 2.555 5.09 2.915 4.75 2.915 4.75 2.325 5.88 2.325 5.88 1.305 5.195 1.305 5.195 0.76 3.7 0.76 3.7 0.53 5.425 0.53 5.425 1.07 7.39 1.07 7.39 1.305 6.11 1.305  ;
        POLYGON 9.64 3.16 12.16 3.16 12.16 3.39 9.64 3.39  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor3_1

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor3_2
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor3_2 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 16.24 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.05 1.265 4.535 1.265 4.535 1.535 2.05 1.535  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.892 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.075 1.49 1.305 1.49 1.305 2.225 3.56 2.225 3.835 2.225 3.835 1.765 4.8 1.765 4.8 1.485 5.695 1.485 5.695 1.72 5.095 1.72 5.095 2.095 4.065 2.095 4.065 2.455 3.56 2.455 2.275 2.455 2.275 2.66 1.075 2.66  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.5355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.115 1.825 9.61 1.825 10.71 1.825 10.71 2.095 9.61 2.095 8.115 2.095  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 1.7952 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.29 2.36 15.21 2.36 15.46 2.36 15.46 1.56 13.29 1.56 13.29 0.655 13.52 0.655 13.52 1.24 15.53 1.24 15.53 0.655 15.76 0.655 15.76 3.36 15.24 3.36 15.24 2.68 15.21 2.68 13.52 2.68 13.52 3.36 13.29 3.36  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.725 3.62 2.725 2.735 3.065 2.735 3.065 3.62 3.56 3.62 6.07 3.62 6.525 3.62 6.525 2.68 6.81 2.68 6.81 3.62 8.775 3.62 8.775 2.795 9.135 2.795 9.135 3.62 11.99 3.62 11.99 3.28 12.355 3.28 12.355 3.62 14.31 3.62 14.31 3.015 14.54 3.015 14.54 3.62 15.21 3.62 16.24 3.62 16.24 4.22 15.21 4.22 6.07 4.22 3.56 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 16.24 -0.3 16.24 0.3 14.64 0.3 14.64 0.905 14.41 0.905 14.41 0.3 8.88 0.3 8.88 0.76 8.535 0.76 8.535 0.3 6.095 0.3 6.095 0.76 5.755 0.76 5.755 0.3 2.935 0.3 2.935 0.775 2.595 0.775 2.595 0.3 0.695 0.3 0.695 0.76 0.355 0.76 0.355 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 0.51 0.99 1.475 0.99 1.475 0.53 1.815 0.53 1.815 1.765 3.56 1.765 3.56 1.995 1.535 1.995 1.535 1.22 0.74 1.22 0.74 3.03 0.51 3.03  ;
        POLYGON 3.735 2.735 4.095 2.735 4.095 3.16 5.785 3.16 5.785 2.68 6.07 2.68 6.07 3.39 3.735 3.39  ;
        POLYGON 6.485 0.53 7.885 0.53 7.885 0.99 9.61 0.99 9.61 1.555 9.27 1.555 9.27 1.22 7.885 1.22 7.885 2.78 7.545 2.78 7.545 0.76 6.485 0.76  ;
        POLYGON 4.72 2.605 5.325 2.605 5.325 1.99 7.01 1.99 7.01 1.22 5.24 1.22 5.24 0.76 3.625 0.76 3.625 0.53 5.47 0.53 5.47 0.99 7.27 0.99 7.27 3.01 8.16 3.01 8.16 2.33 11.105 2.33 11.105 1.67 11.76 1.67 11.76 1.9 11.335 1.9 11.335 2.565 8.445 2.565 8.445 3.24 7.04 3.24 7.04 2.22 5.555 2.22 5.555 2.835 4.72 2.835  ;
        POLYGON 9.795 0.53 12.865 0.53 12.865 0.76 9.795 0.76  ;
        POLYGON 9.75 2.815 12.125 2.815 12.125 1.22 11.17 1.22 11.17 0.99 12.355 0.99 12.355 1.825 15.21 1.825 15.21 2.095 12.355 2.095 12.355 3.05 9.75 3.05  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor3_2

# Copyright 2022 GlobalFoundries PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.

MACRO gf180mcu_fd_sc_mcu7t5v0__xor3_4
  CLASS core ;
  FOREIGN gf180mcu_fd_sc_mcu7t5v0__xor3_4 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  SIZE 18.48 BY 3.92 ;
  PIN A1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.88 1.265 4.36 1.265 4.36 1.535 1.88 1.535  ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.8045 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.865 1.6 1.105 1.6 1.105 2.225 3.41 2.225 3.645 2.225 3.645 1.82 4.615 1.82 4.615 1.56 5.36 1.56 5.36 1.79 4.895 1.79 4.895 2.095 3.875 2.095 3.875 2.455 3.41 2.455 2.1 2.455 2.1 2.71 0.865 2.71  ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    ANTENNAGATEAREA 1.4355 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.91 1.82 9.555 1.82 10.6 1.82 10.6 2.115 9.555 2.115 7.91 2.115  ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 2.978 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.025 2.36 17.225 2.36 17.48 2.36 17.48 1.56 13.025 1.56 13.025 0.6 13.335 0.6 13.335 1.24 15.265 1.24 15.265 0.6 15.575 0.6 15.575 1.24 17.505 1.24 17.505 0.6 17.815 0.6 17.815 3.325 17.37 3.325 17.37 2.68 17.225 2.68 15.69 2.68 15.69 3.315 15.265 3.315 15.265 2.68 13.505 2.68 13.505 3.315 13.025 3.315  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 3.62 2.33 3.62 2.33 2.685 2.67 2.685 2.67 3.62 3.41 3.62 5.875 3.62 6.365 3.62 6.365 2.485 6.595 2.485 6.595 3.62 8.57 3.62 8.57 2.805 8.91 2.805 8.91 3.62 12.23 3.62 12.23 3.285 12.57 3.285 12.57 3.62 14.225 3.62 14.225 2.94 14.455 2.94 14.455 3.62 16.415 3.62 16.415 2.94 16.645 2.94 16.645 3.62 17.225 3.62 18.48 3.62 18.48 4.22 17.225 4.22 5.875 4.22 3.41 4.22 0 4.22  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        POLYGON 0 -0.3 18.48 -0.3 18.48 0.3 16.695 0.3 16.695 0.84 16.465 0.84 16.465 0.3 14.455 0.3 14.455 0.85 14.225 0.85 14.225 0.3 8.69 0.3 8.69 0.775 8.35 0.775 8.35 0.3 5.93 0.3 5.93 0.76 5.59 0.76 5.59 0.3 2.77 0.3 2.77 0.76 2.43 0.76 2.43 0.3 0.53 0.3 0.53 0.76 0.19 0.76 0.19 0.3 0 0.3  ;
    END
  END VSS
  OBS
      LAYER Metal1 ;
        POLYGON 1.085 1.12 1.58 1.12 1.58 1.765 3.41 1.765 3.41 1.995 1.35 1.995 1.35 1.355 0.575 1.355 0.575 2.98 0.345 2.98 0.345 1.12 0.835 1.12 0.835 0.53 1.65 0.53 1.65 0.76 1.085 0.76  ;
        POLYGON 3.55 2.685 3.89 2.685 3.89 3.16 5.645 3.16 5.645 2.61 5.875 2.61 5.875 3.39 3.55 3.39  ;
        POLYGON 6.31 0.53 7.615 0.53 7.615 1.35 9.555 1.35 9.555 1.585 7.615 1.585 7.615 2.845 7.385 2.845 7.385 0.765 6.31 0.765  ;
        POLYGON 4.57 2.685 5.14 2.685 5.14 2.025 5.705 2.025 5.705 1.305 5.035 1.305 5.035 0.76 3.55 0.76 3.55 0.53 5.265 0.53 5.265 1.075 7.115 1.075 7.115 3.14 7.97 3.14 7.97 2.345 11.765 2.345 11.765 1.695 11.995 1.695 11.995 2.575 8.205 2.575 8.205 3.39 6.885 3.39 6.885 1.305 5.935 1.305 5.935 2.26 5.37 2.26 5.37 2.915 4.57 2.915  ;
        POLYGON 9.56 0.53 12.68 0.53 12.68 0.76 9.56 0.76  ;
        POLYGON 9.635 2.815 12.345 2.815 12.345 1.22 10.98 1.22 10.98 0.99 12.575 0.99 12.575 1.825 17.225 1.825 17.225 2.095 12.575 2.095 12.575 3.05 9.635 3.05  ;
  END
END gf180mcu_fd_sc_mcu7t5v0__xor3_4


END LIBRARY
