VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_256x64
  FOREIGN fakeram_256x64 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 8.360 BY 67.200 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.048 0.024 0.072 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.528 0.024 0.552 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.008 0.024 1.032 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.488 0.024 1.512 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.968 0.024 1.992 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.448 0.024 2.472 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.928 0.024 2.952 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.408 0.024 3.432 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.888 0.024 3.912 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.368 0.024 4.392 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.848 0.024 4.872 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.328 0.024 5.352 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.808 0.024 5.832 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.288 0.024 6.312 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.768 0.024 6.792 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.248 0.024 7.272 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.728 0.024 7.752 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.208 0.024 8.232 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.688 0.024 8.712 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.168 0.024 9.192 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.648 0.024 9.672 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.128 0.024 10.152 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.608 0.024 10.632 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.088 0.024 11.112 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.568 0.024 11.592 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.048 0.024 12.072 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.528 0.024 12.552 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.008 0.024 13.032 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.488 0.024 13.512 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.968 0.024 13.992 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.448 0.024 14.472 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.928 0.024 14.952 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.408 0.024 15.432 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.888 0.024 15.912 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.368 0.024 16.392 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.848 0.024 16.872 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.328 0.024 17.352 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.808 0.024 17.832 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.288 0.024 18.312 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.768 0.024 18.792 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.248 0.024 19.272 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.728 0.024 19.752 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.208 0.024 20.232 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.688 0.024 20.712 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.168 0.024 21.192 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.648 0.024 21.672 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.128 0.024 22.152 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.608 0.024 22.632 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.088 0.024 23.112 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.568 0.024 23.592 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.048 0.024 24.072 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.528 0.024 24.552 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.008 0.024 25.032 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.488 0.024 25.512 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.968 0.024 25.992 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.448 0.024 26.472 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.928 0.024 26.952 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.408 0.024 27.432 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.888 0.024 27.912 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.368 0.024 28.392 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.848 0.024 28.872 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.328 0.024 29.352 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.808 0.024 29.832 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.288 0.024 30.312 ;
    END
  END rd_out[63]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.384 0.024 30.408 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.864 0.024 30.888 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.344 0.024 31.368 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.824 0.024 31.848 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.304 0.024 32.328 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.784 0.024 32.808 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 33.264 0.024 33.288 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 33.744 0.024 33.768 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 34.224 0.024 34.248 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 34.704 0.024 34.728 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 35.184 0.024 35.208 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 35.664 0.024 35.688 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.144 0.024 36.168 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.624 0.024 36.648 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.104 0.024 37.128 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.584 0.024 37.608 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 38.064 0.024 38.088 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 38.544 0.024 38.568 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 39.024 0.024 39.048 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 39.504 0.024 39.528 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 39.984 0.024 40.008 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 40.464 0.024 40.488 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 40.944 0.024 40.968 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 41.424 0.024 41.448 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 41.904 0.024 41.928 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 42.384 0.024 42.408 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 42.864 0.024 42.888 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 43.344 0.024 43.368 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 43.824 0.024 43.848 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 44.304 0.024 44.328 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 44.784 0.024 44.808 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 45.264 0.024 45.288 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 45.744 0.024 45.768 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 46.224 0.024 46.248 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 46.704 0.024 46.728 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 47.184 0.024 47.208 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 47.664 0.024 47.688 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 48.144 0.024 48.168 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 48.624 0.024 48.648 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.104 0.024 49.128 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.584 0.024 49.608 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 50.064 0.024 50.088 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 50.544 0.024 50.568 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.024 0.024 51.048 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.504 0.024 51.528 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.984 0.024 52.008 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 52.464 0.024 52.488 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 52.944 0.024 52.968 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 53.424 0.024 53.448 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 53.904 0.024 53.928 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.384 0.024 54.408 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.864 0.024 54.888 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 55.344 0.024 55.368 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 55.824 0.024 55.848 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 56.304 0.024 56.328 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 56.784 0.024 56.808 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 57.264 0.024 57.288 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 57.744 0.024 57.768 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 58.224 0.024 58.248 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 58.704 0.024 58.728 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.184 0.024 59.208 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.664 0.024 59.688 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 60.144 0.024 60.168 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 60.624 0.024 60.648 ;
    END
  END wd_in[63]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 60.720 0.024 60.744 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 61.200 0.024 61.224 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 61.680 0.024 61.704 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 62.160 0.024 62.184 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 62.640 0.024 62.664 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 63.120 0.024 63.144 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 63.600 0.024 63.624 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 64.080 0.024 64.104 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 64.176 0.024 64.200 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 64.656 0.024 64.680 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 65.136 0.024 65.160 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.000 8.312 0.096 ;
      RECT 0.048 0.768 8.312 0.864 ;
      RECT 0.048 1.536 8.312 1.632 ;
      RECT 0.048 2.304 8.312 2.400 ;
      RECT 0.048 3.072 8.312 3.168 ;
      RECT 0.048 3.840 8.312 3.936 ;
      RECT 0.048 4.608 8.312 4.704 ;
      RECT 0.048 5.376 8.312 5.472 ;
      RECT 0.048 6.144 8.312 6.240 ;
      RECT 0.048 6.912 8.312 7.008 ;
      RECT 0.048 7.680 8.312 7.776 ;
      RECT 0.048 8.448 8.312 8.544 ;
      RECT 0.048 9.216 8.312 9.312 ;
      RECT 0.048 9.984 8.312 10.080 ;
      RECT 0.048 10.752 8.312 10.848 ;
      RECT 0.048 11.520 8.312 11.616 ;
      RECT 0.048 12.288 8.312 12.384 ;
      RECT 0.048 13.056 8.312 13.152 ;
      RECT 0.048 13.824 8.312 13.920 ;
      RECT 0.048 14.592 8.312 14.688 ;
      RECT 0.048 15.360 8.312 15.456 ;
      RECT 0.048 16.128 8.312 16.224 ;
      RECT 0.048 16.896 8.312 16.992 ;
      RECT 0.048 17.664 8.312 17.760 ;
      RECT 0.048 18.432 8.312 18.528 ;
      RECT 0.048 19.200 8.312 19.296 ;
      RECT 0.048 19.968 8.312 20.064 ;
      RECT 0.048 20.736 8.312 20.832 ;
      RECT 0.048 21.504 8.312 21.600 ;
      RECT 0.048 22.272 8.312 22.368 ;
      RECT 0.048 23.040 8.312 23.136 ;
      RECT 0.048 23.808 8.312 23.904 ;
      RECT 0.048 24.576 8.312 24.672 ;
      RECT 0.048 25.344 8.312 25.440 ;
      RECT 0.048 26.112 8.312 26.208 ;
      RECT 0.048 26.880 8.312 26.976 ;
      RECT 0.048 27.648 8.312 27.744 ;
      RECT 0.048 28.416 8.312 28.512 ;
      RECT 0.048 29.184 8.312 29.280 ;
      RECT 0.048 29.952 8.312 30.048 ;
      RECT 0.048 30.720 8.312 30.816 ;
      RECT 0.048 31.488 8.312 31.584 ;
      RECT 0.048 32.256 8.312 32.352 ;
      RECT 0.048 33.024 8.312 33.120 ;
      RECT 0.048 33.792 8.312 33.888 ;
      RECT 0.048 34.560 8.312 34.656 ;
      RECT 0.048 35.328 8.312 35.424 ;
      RECT 0.048 36.096 8.312 36.192 ;
      RECT 0.048 36.864 8.312 36.960 ;
      RECT 0.048 37.632 8.312 37.728 ;
      RECT 0.048 38.400 8.312 38.496 ;
      RECT 0.048 39.168 8.312 39.264 ;
      RECT 0.048 39.936 8.312 40.032 ;
      RECT 0.048 40.704 8.312 40.800 ;
      RECT 0.048 41.472 8.312 41.568 ;
      RECT 0.048 42.240 8.312 42.336 ;
      RECT 0.048 43.008 8.312 43.104 ;
      RECT 0.048 43.776 8.312 43.872 ;
      RECT 0.048 44.544 8.312 44.640 ;
      RECT 0.048 45.312 8.312 45.408 ;
      RECT 0.048 46.080 8.312 46.176 ;
      RECT 0.048 46.848 8.312 46.944 ;
      RECT 0.048 47.616 8.312 47.712 ;
      RECT 0.048 48.384 8.312 48.480 ;
      RECT 0.048 49.152 8.312 49.248 ;
      RECT 0.048 49.920 8.312 50.016 ;
      RECT 0.048 50.688 8.312 50.784 ;
      RECT 0.048 51.456 8.312 51.552 ;
      RECT 0.048 52.224 8.312 52.320 ;
      RECT 0.048 52.992 8.312 53.088 ;
      RECT 0.048 53.760 8.312 53.856 ;
      RECT 0.048 54.528 8.312 54.624 ;
      RECT 0.048 55.296 8.312 55.392 ;
      RECT 0.048 56.064 8.312 56.160 ;
      RECT 0.048 56.832 8.312 56.928 ;
      RECT 0.048 57.600 8.312 57.696 ;
      RECT 0.048 58.368 8.312 58.464 ;
      RECT 0.048 59.136 8.312 59.232 ;
      RECT 0.048 59.904 8.312 60.000 ;
      RECT 0.048 60.672 8.312 60.768 ;
      RECT 0.048 61.440 8.312 61.536 ;
      RECT 0.048 62.208 8.312 62.304 ;
      RECT 0.048 62.976 8.312 63.072 ;
      RECT 0.048 63.744 8.312 63.840 ;
      RECT 0.048 64.512 8.312 64.608 ;
      RECT 0.048 65.280 8.312 65.376 ;
      RECT 0.048 66.048 8.312 66.144 ;
      RECT 0.048 66.816 8.312 66.912 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.384 8.312 0.480 ;
      RECT 0.048 1.152 8.312 1.248 ;
      RECT 0.048 1.920 8.312 2.016 ;
      RECT 0.048 2.688 8.312 2.784 ;
      RECT 0.048 3.456 8.312 3.552 ;
      RECT 0.048 4.224 8.312 4.320 ;
      RECT 0.048 4.992 8.312 5.088 ;
      RECT 0.048 5.760 8.312 5.856 ;
      RECT 0.048 6.528 8.312 6.624 ;
      RECT 0.048 7.296 8.312 7.392 ;
      RECT 0.048 8.064 8.312 8.160 ;
      RECT 0.048 8.832 8.312 8.928 ;
      RECT 0.048 9.600 8.312 9.696 ;
      RECT 0.048 10.368 8.312 10.464 ;
      RECT 0.048 11.136 8.312 11.232 ;
      RECT 0.048 11.904 8.312 12.000 ;
      RECT 0.048 12.672 8.312 12.768 ;
      RECT 0.048 13.440 8.312 13.536 ;
      RECT 0.048 14.208 8.312 14.304 ;
      RECT 0.048 14.976 8.312 15.072 ;
      RECT 0.048 15.744 8.312 15.840 ;
      RECT 0.048 16.512 8.312 16.608 ;
      RECT 0.048 17.280 8.312 17.376 ;
      RECT 0.048 18.048 8.312 18.144 ;
      RECT 0.048 18.816 8.312 18.912 ;
      RECT 0.048 19.584 8.312 19.680 ;
      RECT 0.048 20.352 8.312 20.448 ;
      RECT 0.048 21.120 8.312 21.216 ;
      RECT 0.048 21.888 8.312 21.984 ;
      RECT 0.048 22.656 8.312 22.752 ;
      RECT 0.048 23.424 8.312 23.520 ;
      RECT 0.048 24.192 8.312 24.288 ;
      RECT 0.048 24.960 8.312 25.056 ;
      RECT 0.048 25.728 8.312 25.824 ;
      RECT 0.048 26.496 8.312 26.592 ;
      RECT 0.048 27.264 8.312 27.360 ;
      RECT 0.048 28.032 8.312 28.128 ;
      RECT 0.048 28.800 8.312 28.896 ;
      RECT 0.048 29.568 8.312 29.664 ;
      RECT 0.048 30.336 8.312 30.432 ;
      RECT 0.048 31.104 8.312 31.200 ;
      RECT 0.048 31.872 8.312 31.968 ;
      RECT 0.048 32.640 8.312 32.736 ;
      RECT 0.048 33.408 8.312 33.504 ;
      RECT 0.048 34.176 8.312 34.272 ;
      RECT 0.048 34.944 8.312 35.040 ;
      RECT 0.048 35.712 8.312 35.808 ;
      RECT 0.048 36.480 8.312 36.576 ;
      RECT 0.048 37.248 8.312 37.344 ;
      RECT 0.048 38.016 8.312 38.112 ;
      RECT 0.048 38.784 8.312 38.880 ;
      RECT 0.048 39.552 8.312 39.648 ;
      RECT 0.048 40.320 8.312 40.416 ;
      RECT 0.048 41.088 8.312 41.184 ;
      RECT 0.048 41.856 8.312 41.952 ;
      RECT 0.048 42.624 8.312 42.720 ;
      RECT 0.048 43.392 8.312 43.488 ;
      RECT 0.048 44.160 8.312 44.256 ;
      RECT 0.048 44.928 8.312 45.024 ;
      RECT 0.048 45.696 8.312 45.792 ;
      RECT 0.048 46.464 8.312 46.560 ;
      RECT 0.048 47.232 8.312 47.328 ;
      RECT 0.048 48.000 8.312 48.096 ;
      RECT 0.048 48.768 8.312 48.864 ;
      RECT 0.048 49.536 8.312 49.632 ;
      RECT 0.048 50.304 8.312 50.400 ;
      RECT 0.048 51.072 8.312 51.168 ;
      RECT 0.048 51.840 8.312 51.936 ;
      RECT 0.048 52.608 8.312 52.704 ;
      RECT 0.048 53.376 8.312 53.472 ;
      RECT 0.048 54.144 8.312 54.240 ;
      RECT 0.048 54.912 8.312 55.008 ;
      RECT 0.048 55.680 8.312 55.776 ;
      RECT 0.048 56.448 8.312 56.544 ;
      RECT 0.048 57.216 8.312 57.312 ;
      RECT 0.048 57.984 8.312 58.080 ;
      RECT 0.048 58.752 8.312 58.848 ;
      RECT 0.048 59.520 8.312 59.616 ;
      RECT 0.048 60.288 8.312 60.384 ;
      RECT 0.048 61.056 8.312 61.152 ;
      RECT 0.048 61.824 8.312 61.920 ;
      RECT 0.048 62.592 8.312 62.688 ;
      RECT 0.048 63.360 8.312 63.456 ;
      RECT 0.048 64.128 8.312 64.224 ;
      RECT 0.048 64.896 8.312 64.992 ;
      RECT 0.048 65.664 8.312 65.760 ;
      RECT 0.048 66.432 8.312 66.528 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 8.360 67.200 ;
    LAYER M2 ;
    RECT 0 0 8.360 67.200 ;
    LAYER M3 ;
    RECT 0 0 8.360 67.200 ;
    LAYER M4 ;
    RECT 0.024 0 0.048 67.200 ;
    RECT 8.312 0 8.360 67.200 ;
    RECT 0.048 0.000 8.312 0.000 ;
    RECT 0.048 0.096 8.312 0.384 ;
    RECT 0.048 0.480 8.312 0.768 ;
    RECT 0.048 0.864 8.312 1.152 ;
    RECT 0.048 1.248 8.312 1.536 ;
    RECT 0.048 1.632 8.312 1.920 ;
    RECT 0.048 2.016 8.312 2.304 ;
    RECT 0.048 2.400 8.312 2.688 ;
    RECT 0.048 2.784 8.312 3.072 ;
    RECT 0.048 3.168 8.312 3.456 ;
    RECT 0.048 3.552 8.312 3.840 ;
    RECT 0.048 3.936 8.312 4.224 ;
    RECT 0.048 4.320 8.312 4.608 ;
    RECT 0.048 4.704 8.312 4.992 ;
    RECT 0.048 5.088 8.312 5.376 ;
    RECT 0.048 5.472 8.312 5.760 ;
    RECT 0.048 5.856 8.312 6.144 ;
    RECT 0.048 6.240 8.312 6.528 ;
    RECT 0.048 6.624 8.312 6.912 ;
    RECT 0.048 7.008 8.312 7.296 ;
    RECT 0.048 7.392 8.312 7.680 ;
    RECT 0.048 7.776 8.312 8.064 ;
    RECT 0.048 8.160 8.312 8.448 ;
    RECT 0.048 8.544 8.312 8.832 ;
    RECT 0.048 8.928 8.312 9.216 ;
    RECT 0.048 9.312 8.312 9.600 ;
    RECT 0.048 9.696 8.312 9.984 ;
    RECT 0.048 10.080 8.312 10.368 ;
    RECT 0.048 10.464 8.312 10.752 ;
    RECT 0.048 10.848 8.312 11.136 ;
    RECT 0.048 11.232 8.312 11.520 ;
    RECT 0.048 11.616 8.312 11.904 ;
    RECT 0.048 12.000 8.312 12.288 ;
    RECT 0.048 12.384 8.312 12.672 ;
    RECT 0.048 12.768 8.312 13.056 ;
    RECT 0.048 13.152 8.312 13.440 ;
    RECT 0.048 13.536 8.312 13.824 ;
    RECT 0.048 13.920 8.312 14.208 ;
    RECT 0.048 14.304 8.312 14.592 ;
    RECT 0.048 14.688 8.312 14.976 ;
    RECT 0.048 15.072 8.312 15.360 ;
    RECT 0.048 15.456 8.312 15.744 ;
    RECT 0.048 15.840 8.312 16.128 ;
    RECT 0.048 16.224 8.312 16.512 ;
    RECT 0.048 16.608 8.312 16.896 ;
    RECT 0.048 16.992 8.312 17.280 ;
    RECT 0.048 17.376 8.312 17.664 ;
    RECT 0.048 17.760 8.312 18.048 ;
    RECT 0.048 18.144 8.312 18.432 ;
    RECT 0.048 18.528 8.312 18.816 ;
    RECT 0.048 18.912 8.312 19.200 ;
    RECT 0.048 19.296 8.312 19.584 ;
    RECT 0.048 19.680 8.312 19.968 ;
    RECT 0.048 20.064 8.312 20.352 ;
    RECT 0.048 20.448 8.312 20.736 ;
    RECT 0.048 20.832 8.312 21.120 ;
    RECT 0.048 21.216 8.312 21.504 ;
    RECT 0.048 21.600 8.312 21.888 ;
    RECT 0.048 21.984 8.312 22.272 ;
    RECT 0.048 22.368 8.312 22.656 ;
    RECT 0.048 22.752 8.312 23.040 ;
    RECT 0.048 23.136 8.312 23.424 ;
    RECT 0.048 23.520 8.312 23.808 ;
    RECT 0.048 23.904 8.312 24.192 ;
    RECT 0.048 24.288 8.312 24.576 ;
    RECT 0.048 24.672 8.312 24.960 ;
    RECT 0.048 25.056 8.312 25.344 ;
    RECT 0.048 25.440 8.312 25.728 ;
    RECT 0.048 25.824 8.312 26.112 ;
    RECT 0.048 26.208 8.312 26.496 ;
    RECT 0.048 26.592 8.312 26.880 ;
    RECT 0.048 26.976 8.312 27.264 ;
    RECT 0.048 27.360 8.312 27.648 ;
    RECT 0.048 27.744 8.312 28.032 ;
    RECT 0.048 28.128 8.312 28.416 ;
    RECT 0.048 28.512 8.312 28.800 ;
    RECT 0.048 28.896 8.312 29.184 ;
    RECT 0.048 29.280 8.312 29.568 ;
    RECT 0.048 29.664 8.312 29.952 ;
    RECT 0.048 30.048 8.312 30.336 ;
    RECT 0.048 30.432 8.312 30.720 ;
    RECT 0.048 30.816 8.312 31.104 ;
    RECT 0.048 31.200 8.312 31.488 ;
    RECT 0.048 31.584 8.312 31.872 ;
    RECT 0.048 31.968 8.312 32.256 ;
    RECT 0.048 32.352 8.312 32.640 ;
    RECT 0.048 32.736 8.312 33.024 ;
    RECT 0.048 33.120 8.312 33.408 ;
    RECT 0.048 33.504 8.312 33.792 ;
    RECT 0.048 33.888 8.312 34.176 ;
    RECT 0.048 34.272 8.312 34.560 ;
    RECT 0.048 34.656 8.312 34.944 ;
    RECT 0.048 35.040 8.312 35.328 ;
    RECT 0.048 35.424 8.312 35.712 ;
    RECT 0.048 35.808 8.312 36.096 ;
    RECT 0.048 36.192 8.312 36.480 ;
    RECT 0.048 36.576 8.312 36.864 ;
    RECT 0.048 36.960 8.312 37.248 ;
    RECT 0.048 37.344 8.312 37.632 ;
    RECT 0.048 37.728 8.312 38.016 ;
    RECT 0.048 38.112 8.312 38.400 ;
    RECT 0.048 38.496 8.312 38.784 ;
    RECT 0.048 38.880 8.312 39.168 ;
    RECT 0.048 39.264 8.312 39.552 ;
    RECT 0.048 39.648 8.312 39.936 ;
    RECT 0.048 40.032 8.312 40.320 ;
    RECT 0.048 40.416 8.312 40.704 ;
    RECT 0.048 40.800 8.312 41.088 ;
    RECT 0.048 41.184 8.312 41.472 ;
    RECT 0.048 41.568 8.312 41.856 ;
    RECT 0.048 41.952 8.312 42.240 ;
    RECT 0.048 42.336 8.312 42.624 ;
    RECT 0.048 42.720 8.312 43.008 ;
    RECT 0.048 43.104 8.312 43.392 ;
    RECT 0.048 43.488 8.312 43.776 ;
    RECT 0.048 43.872 8.312 44.160 ;
    RECT 0.048 44.256 8.312 44.544 ;
    RECT 0.048 44.640 8.312 44.928 ;
    RECT 0.048 45.024 8.312 45.312 ;
    RECT 0.048 45.408 8.312 45.696 ;
    RECT 0.048 45.792 8.312 46.080 ;
    RECT 0.048 46.176 8.312 46.464 ;
    RECT 0.048 46.560 8.312 46.848 ;
    RECT 0.048 46.944 8.312 47.232 ;
    RECT 0.048 47.328 8.312 47.616 ;
    RECT 0.048 47.712 8.312 48.000 ;
    RECT 0.048 48.096 8.312 48.384 ;
    RECT 0.048 48.480 8.312 48.768 ;
    RECT 0.048 48.864 8.312 49.152 ;
    RECT 0.048 49.248 8.312 49.536 ;
    RECT 0.048 49.632 8.312 49.920 ;
    RECT 0.048 50.016 8.312 50.304 ;
    RECT 0.048 50.400 8.312 50.688 ;
    RECT 0.048 50.784 8.312 51.072 ;
    RECT 0.048 51.168 8.312 51.456 ;
    RECT 0.048 51.552 8.312 51.840 ;
    RECT 0.048 51.936 8.312 52.224 ;
    RECT 0.048 52.320 8.312 52.608 ;
    RECT 0.048 52.704 8.312 52.992 ;
    RECT 0.048 53.088 8.312 53.376 ;
    RECT 0.048 53.472 8.312 53.760 ;
    RECT 0.048 53.856 8.312 54.144 ;
    RECT 0.048 54.240 8.312 54.528 ;
    RECT 0.048 54.624 8.312 54.912 ;
    RECT 0.048 55.008 8.312 55.296 ;
    RECT 0.048 55.392 8.312 55.680 ;
    RECT 0.048 55.776 8.312 56.064 ;
    RECT 0.048 56.160 8.312 56.448 ;
    RECT 0.048 56.544 8.312 56.832 ;
    RECT 0.048 56.928 8.312 57.216 ;
    RECT 0.048 57.312 8.312 57.600 ;
    RECT 0.048 57.696 8.312 57.984 ;
    RECT 0.048 58.080 8.312 58.368 ;
    RECT 0.048 58.464 8.312 58.752 ;
    RECT 0.048 58.848 8.312 59.136 ;
    RECT 0.048 59.232 8.312 59.520 ;
    RECT 0.048 59.616 8.312 59.904 ;
    RECT 0.048 60.000 8.312 60.288 ;
    RECT 0.048 60.384 8.312 60.672 ;
    RECT 0.048 60.768 8.312 61.056 ;
    RECT 0.048 61.152 8.312 61.440 ;
    RECT 0.048 61.536 8.312 61.824 ;
    RECT 0.048 61.920 8.312 62.208 ;
    RECT 0.048 62.304 8.312 62.592 ;
    RECT 0.048 62.688 8.312 62.976 ;
    RECT 0.048 63.072 8.312 63.360 ;
    RECT 0.048 63.456 8.312 63.744 ;
    RECT 0.048 63.840 8.312 64.128 ;
    RECT 0.048 64.224 8.312 64.512 ;
    RECT 0.048 64.608 8.312 64.896 ;
    RECT 0.048 64.992 8.312 65.280 ;
    RECT 0.048 65.376 8.312 65.664 ;
    RECT 0.048 65.760 8.312 66.048 ;
    RECT 0.048 66.144 8.312 66.432 ;
    RECT 0.048 66.528 8.312 66.816 ;
    RECT 0.048 66.912 8.312 67.200 ;
    RECT 0 0.000 0.024 0.048 ;
    RECT 0 0.072 0.024 0.528 ;
    RECT 0 0.552 0.024 1.008 ;
    RECT 0 1.032 0.024 1.488 ;
    RECT 0 1.512 0.024 1.968 ;
    RECT 0 1.992 0.024 2.448 ;
    RECT 0 2.472 0.024 2.928 ;
    RECT 0 2.952 0.024 3.408 ;
    RECT 0 3.432 0.024 3.888 ;
    RECT 0 3.912 0.024 4.368 ;
    RECT 0 4.392 0.024 4.848 ;
    RECT 0 4.872 0.024 5.328 ;
    RECT 0 5.352 0.024 5.808 ;
    RECT 0 5.832 0.024 6.288 ;
    RECT 0 6.312 0.024 6.768 ;
    RECT 0 6.792 0.024 7.248 ;
    RECT 0 7.272 0.024 7.728 ;
    RECT 0 7.752 0.024 8.208 ;
    RECT 0 8.232 0.024 8.688 ;
    RECT 0 8.712 0.024 9.168 ;
    RECT 0 9.192 0.024 9.648 ;
    RECT 0 9.672 0.024 10.128 ;
    RECT 0 10.152 0.024 10.608 ;
    RECT 0 10.632 0.024 11.088 ;
    RECT 0 11.112 0.024 11.568 ;
    RECT 0 11.592 0.024 12.048 ;
    RECT 0 12.072 0.024 12.528 ;
    RECT 0 12.552 0.024 13.008 ;
    RECT 0 13.032 0.024 13.488 ;
    RECT 0 13.512 0.024 13.968 ;
    RECT 0 13.992 0.024 14.448 ;
    RECT 0 14.472 0.024 14.928 ;
    RECT 0 14.952 0.024 15.408 ;
    RECT 0 15.432 0.024 15.888 ;
    RECT 0 15.912 0.024 16.368 ;
    RECT 0 16.392 0.024 16.848 ;
    RECT 0 16.872 0.024 17.328 ;
    RECT 0 17.352 0.024 17.808 ;
    RECT 0 17.832 0.024 18.288 ;
    RECT 0 18.312 0.024 18.768 ;
    RECT 0 18.792 0.024 19.248 ;
    RECT 0 19.272 0.024 19.728 ;
    RECT 0 19.752 0.024 20.208 ;
    RECT 0 20.232 0.024 20.688 ;
    RECT 0 20.712 0.024 21.168 ;
    RECT 0 21.192 0.024 21.648 ;
    RECT 0 21.672 0.024 22.128 ;
    RECT 0 22.152 0.024 22.608 ;
    RECT 0 22.632 0.024 23.088 ;
    RECT 0 23.112 0.024 23.568 ;
    RECT 0 23.592 0.024 24.048 ;
    RECT 0 24.072 0.024 24.528 ;
    RECT 0 24.552 0.024 25.008 ;
    RECT 0 25.032 0.024 25.488 ;
    RECT 0 25.512 0.024 25.968 ;
    RECT 0 25.992 0.024 26.448 ;
    RECT 0 26.472 0.024 26.928 ;
    RECT 0 26.952 0.024 27.408 ;
    RECT 0 27.432 0.024 27.888 ;
    RECT 0 27.912 0.024 28.368 ;
    RECT 0 28.392 0.024 28.848 ;
    RECT 0 28.872 0.024 29.328 ;
    RECT 0 29.352 0.024 29.808 ;
    RECT 0 29.832 0.024 30.288 ;
    RECT 0 30.312 0.024 30.384 ;
    RECT 0 30.408 0.024 30.864 ;
    RECT 0 30.888 0.024 31.344 ;
    RECT 0 31.368 0.024 31.824 ;
    RECT 0 31.848 0.024 32.304 ;
    RECT 0 32.328 0.024 32.784 ;
    RECT 0 32.808 0.024 33.264 ;
    RECT 0 33.288 0.024 33.744 ;
    RECT 0 33.768 0.024 34.224 ;
    RECT 0 34.248 0.024 34.704 ;
    RECT 0 34.728 0.024 35.184 ;
    RECT 0 35.208 0.024 35.664 ;
    RECT 0 35.688 0.024 36.144 ;
    RECT 0 36.168 0.024 36.624 ;
    RECT 0 36.648 0.024 37.104 ;
    RECT 0 37.128 0.024 37.584 ;
    RECT 0 37.608 0.024 38.064 ;
    RECT 0 38.088 0.024 38.544 ;
    RECT 0 38.568 0.024 39.024 ;
    RECT 0 39.048 0.024 39.504 ;
    RECT 0 39.528 0.024 39.984 ;
    RECT 0 40.008 0.024 40.464 ;
    RECT 0 40.488 0.024 40.944 ;
    RECT 0 40.968 0.024 41.424 ;
    RECT 0 41.448 0.024 41.904 ;
    RECT 0 41.928 0.024 42.384 ;
    RECT 0 42.408 0.024 42.864 ;
    RECT 0 42.888 0.024 43.344 ;
    RECT 0 43.368 0.024 43.824 ;
    RECT 0 43.848 0.024 44.304 ;
    RECT 0 44.328 0.024 44.784 ;
    RECT 0 44.808 0.024 45.264 ;
    RECT 0 45.288 0.024 45.744 ;
    RECT 0 45.768 0.024 46.224 ;
    RECT 0 46.248 0.024 46.704 ;
    RECT 0 46.728 0.024 47.184 ;
    RECT 0 47.208 0.024 47.664 ;
    RECT 0 47.688 0.024 48.144 ;
    RECT 0 48.168 0.024 48.624 ;
    RECT 0 48.648 0.024 49.104 ;
    RECT 0 49.128 0.024 49.584 ;
    RECT 0 49.608 0.024 50.064 ;
    RECT 0 50.088 0.024 50.544 ;
    RECT 0 50.568 0.024 51.024 ;
    RECT 0 51.048 0.024 51.504 ;
    RECT 0 51.528 0.024 51.984 ;
    RECT 0 52.008 0.024 52.464 ;
    RECT 0 52.488 0.024 52.944 ;
    RECT 0 52.968 0.024 53.424 ;
    RECT 0 53.448 0.024 53.904 ;
    RECT 0 53.928 0.024 54.384 ;
    RECT 0 54.408 0.024 54.864 ;
    RECT 0 54.888 0.024 55.344 ;
    RECT 0 55.368 0.024 55.824 ;
    RECT 0 55.848 0.024 56.304 ;
    RECT 0 56.328 0.024 56.784 ;
    RECT 0 56.808 0.024 57.264 ;
    RECT 0 57.288 0.024 57.744 ;
    RECT 0 57.768 0.024 58.224 ;
    RECT 0 58.248 0.024 58.704 ;
    RECT 0 58.728 0.024 59.184 ;
    RECT 0 59.208 0.024 59.664 ;
    RECT 0 59.688 0.024 60.144 ;
    RECT 0 60.168 0.024 60.624 ;
    RECT 0 60.648 0.024 60.720 ;
    RECT 0 60.744 0.024 61.200 ;
    RECT 0 61.224 0.024 61.680 ;
    RECT 0 61.704 0.024 62.160 ;
    RECT 0 62.184 0.024 62.640 ;
    RECT 0 62.664 0.024 63.120 ;
    RECT 0 63.144 0.024 63.600 ;
    RECT 0 63.624 0.024 64.080 ;
    RECT 0 64.104 0.024 64.560 ;
    RECT 0 64.584 0.024 65.040 ;
    RECT 0 65.064 0.024 65.520 ;
    RECT 0 65.544 0.024 66.000 ;
    RECT 0 66.024 0.024 66.480 ;
    RECT 0 66.504 0.024 66.960 ;
    RECT 0 66.984 0.024 67.440 ;
    RECT 0 67.464 0.024 67.920 ;
    RECT 0 67.944 0.024 68.400 ;
    RECT 0 68.424 0.024 68.880 ;
    RECT 0 68.904 0.024 69.360 ;
    RECT 0 69.384 0.024 69.840 ;
    RECT 0 69.864 0.024 70.320 ;
    RECT 0 70.344 0.024 70.800 ;
    RECT 0 70.824 0.024 71.280 ;
    RECT 0 71.304 0.024 71.760 ;
    RECT 0 71.784 0.024 72.240 ;
    RECT 0 72.264 0.024 72.720 ;
    RECT 0 72.744 0.024 73.200 ;
    RECT 0 73.224 0.024 73.680 ;
    RECT 0 73.704 0.024 74.160 ;
    RECT 0 74.184 0.024 74.640 ;
    RECT 0 74.664 0.024 75.120 ;
    RECT 0 75.144 0.024 75.600 ;
    RECT 0 75.624 0.024 76.080 ;
    RECT 0 76.104 0.024 76.560 ;
    RECT 0 76.584 0.024 77.040 ;
    RECT 0 77.064 0.024 77.520 ;
    RECT 0 77.544 0.024 78.000 ;
    RECT 0 78.024 0.024 78.480 ;
    RECT 0 78.504 0.024 78.960 ;
    RECT 0 78.984 0.024 79.440 ;
    RECT 0 79.464 0.024 79.920 ;
    RECT 0 79.944 0.024 80.400 ;
    RECT 0 80.424 0.024 80.880 ;
    RECT 0 80.904 0.024 81.360 ;
    RECT 0 81.384 0.024 81.840 ;
    RECT 0 81.864 0.024 82.320 ;
    RECT 0 82.344 0.024 82.800 ;
    RECT 0 82.824 0.024 83.280 ;
    RECT 0 83.304 0.024 83.760 ;
    RECT 0 83.784 0.024 84.240 ;
    RECT 0 84.264 0.024 84.720 ;
    RECT 0 84.744 0.024 85.200 ;
    RECT 0 85.224 0.024 85.680 ;
    RECT 0 85.704 0.024 86.160 ;
    RECT 0 86.184 0.024 86.640 ;
    RECT 0 86.664 0.024 87.120 ;
    RECT 0 87.144 0.024 87.600 ;
    RECT 0 87.624 0.024 88.080 ;
    RECT 0 88.104 0.024 88.560 ;
    RECT 0 88.584 0.024 89.040 ;
    RECT 0 89.064 0.024 89.520 ;
    RECT 0 89.544 0.024 90.000 ;
    RECT 0 90.024 0.024 90.480 ;
    RECT 0 90.504 0.024 90.960 ;
    RECT 0 90.984 0.024 91.056 ;
    RECT 0 91.080 0.024 91.536 ;
    RECT 0 91.560 0.024 92.016 ;
    RECT 0 92.040 0.024 92.496 ;
    RECT 0 92.520 0.024 92.976 ;
    RECT 0 93.000 0.024 93.456 ;
    RECT 0 93.480 0.024 93.936 ;
    RECT 0 93.960 0.024 94.416 ;
    RECT 0 94.440 0.024 94.512 ;
    RECT 0 94.536 0.024 94.992 ;
    RECT 0 95.016 0.024 95.472 ;
    RECT 0 95.496 0.024 67.200 ;
#    LAYER OVERLAP ;
#    RECT 0 0 8.360 67.200 ;
  END
END fakeram_256x64

END LIBRARY
