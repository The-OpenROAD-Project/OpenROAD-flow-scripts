VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO or1200_spram3
  FOREIGN or1200_spram3 0 0 ;
  CLASS BLOCK ;
  SIZE 116.625 BY 139.55 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.94 122.7 115.34 124.1 ;
        RECT  2.94 82.7 115.34 84.1 ;
        RECT  2.94 42.7 115.34 44.1 ;
        RECT  2.94 2.7 115.34 4.1 ;
      LAYER metal4 ;
        RECT  115.04 1.33 115.24 135.87 ;
        RECT  59.04 1.33 59.24 135.87 ;
        RECT  3.04 1.33 3.24 135.87 ;
      LAYER metal1 ;
        RECT  1.14 135.75 115.52 135.85 ;
        RECT  1.14 132.95 115.52 133.05 ;
        RECT  1.14 130.15 115.52 130.25 ;
        RECT  1.14 127.35 115.52 127.45 ;
        RECT  1.14 124.55 115.52 124.65 ;
        RECT  1.14 121.75 115.52 121.85 ;
        RECT  1.14 118.95 115.52 119.05 ;
        RECT  1.14 116.15 115.52 116.25 ;
        RECT  1.14 113.35 115.52 113.45 ;
        RECT  1.14 110.55 115.52 110.65 ;
        RECT  1.14 107.75 115.52 107.85 ;
        RECT  1.14 104.95 115.52 105.05 ;
        RECT  1.14 102.15 115.52 102.25 ;
        RECT  1.14 99.35 115.52 99.45 ;
        RECT  1.14 96.55 115.52 96.65 ;
        RECT  1.14 93.75 115.52 93.85 ;
        RECT  1.14 90.95 115.52 91.05 ;
        RECT  1.14 88.15 115.52 88.25 ;
        RECT  1.14 85.35 115.52 85.45 ;
        RECT  1.14 82.55 115.52 82.65 ;
        RECT  1.14 79.75 115.52 79.85 ;
        RECT  1.14 76.95 115.52 77.05 ;
        RECT  1.14 74.15 115.52 74.25 ;
        RECT  1.14 71.35 115.52 71.45 ;
        RECT  1.14 68.55 115.52 68.65 ;
        RECT  1.14 65.75 115.52 65.85 ;
        RECT  1.14 62.95 115.52 63.05 ;
        RECT  1.14 60.15 115.52 60.25 ;
        RECT  1.14 57.35 115.52 57.45 ;
        RECT  1.14 54.55 115.52 54.65 ;
        RECT  1.14 51.75 115.52 51.85 ;
        RECT  1.14 48.95 115.52 49.05 ;
        RECT  1.14 46.15 115.52 46.25 ;
        RECT  1.14 43.35 115.52 43.45 ;
        RECT  1.14 40.55 115.52 40.65 ;
        RECT  1.14 37.75 115.52 37.85 ;
        RECT  1.14 34.95 115.52 35.05 ;
        RECT  1.14 32.15 115.52 32.25 ;
        RECT  1.14 29.35 115.52 29.45 ;
        RECT  1.14 26.55 115.52 26.65 ;
        RECT  1.14 23.75 115.52 23.85 ;
        RECT  1.14 20.95 115.52 21.05 ;
        RECT  1.14 18.15 115.52 18.25 ;
        RECT  1.14 15.35 115.52 15.45 ;
        RECT  1.14 12.55 115.52 12.65 ;
        RECT  1.14 9.75 115.52 9.85 ;
        RECT  1.14 6.95 115.52 7.05 ;
        RECT  1.14 4.15 115.52 4.25 ;
        RECT  1.14 1.35 115.52 1.45 ;
      VIA 115.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 1.4 via1_2_400_200_1_1_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.94 102.7 87.34 104.1 ;
        RECT  30.94 62.7 87.34 64.1 ;
        RECT  30.94 22.7 87.34 24.1 ;
      LAYER metal4 ;
        RECT  87.04 2.73 87.24 137.27 ;
        RECT  31.04 2.73 31.24 137.27 ;
      LAYER metal1 ;
        RECT  1.14 137.15 115.52 137.25 ;
        RECT  1.14 134.35 115.52 134.45 ;
        RECT  1.14 131.55 115.52 131.65 ;
        RECT  1.14 128.75 115.52 128.85 ;
        RECT  1.14 125.95 115.52 126.05 ;
        RECT  1.14 123.15 115.52 123.25 ;
        RECT  1.14 120.35 115.52 120.45 ;
        RECT  1.14 117.55 115.52 117.65 ;
        RECT  1.14 114.75 115.52 114.85 ;
        RECT  1.14 111.95 115.52 112.05 ;
        RECT  1.14 109.15 115.52 109.25 ;
        RECT  1.14 106.35 115.52 106.45 ;
        RECT  1.14 103.55 115.52 103.65 ;
        RECT  1.14 100.75 115.52 100.85 ;
        RECT  1.14 97.95 115.52 98.05 ;
        RECT  1.14 95.15 115.52 95.25 ;
        RECT  1.14 92.35 115.52 92.45 ;
        RECT  1.14 89.55 115.52 89.65 ;
        RECT  1.14 86.75 115.52 86.85 ;
        RECT  1.14 83.95 115.52 84.05 ;
        RECT  1.14 81.15 115.52 81.25 ;
        RECT  1.14 78.35 115.52 78.45 ;
        RECT  1.14 75.55 115.52 75.65 ;
        RECT  1.14 72.75 115.52 72.85 ;
        RECT  1.14 69.95 115.52 70.05 ;
        RECT  1.14 67.15 115.52 67.25 ;
        RECT  1.14 64.35 115.52 64.45 ;
        RECT  1.14 61.55 115.52 61.65 ;
        RECT  1.14 58.75 115.52 58.85 ;
        RECT  1.14 55.95 115.52 56.05 ;
        RECT  1.14 53.15 115.52 53.25 ;
        RECT  1.14 50.35 115.52 50.45 ;
        RECT  1.14 47.55 115.52 47.65 ;
        RECT  1.14 44.75 115.52 44.85 ;
        RECT  1.14 41.95 115.52 42.05 ;
        RECT  1.14 39.15 115.52 39.25 ;
        RECT  1.14 36.35 115.52 36.45 ;
        RECT  1.14 33.55 115.52 33.65 ;
        RECT  1.14 30.75 115.52 30.85 ;
        RECT  1.14 27.95 115.52 28.05 ;
        RECT  1.14 25.15 115.52 25.25 ;
        RECT  1.14 22.35 115.52 22.45 ;
        RECT  1.14 19.55 115.52 19.65 ;
        RECT  1.14 16.75 115.52 16.85 ;
        RECT  1.14 13.95 115.52 14.05 ;
        RECT  1.14 11.15 115.52 11.25 ;
        RECT  1.14 8.35 115.52 8.45 ;
        RECT  1.14 5.55 115.52 5.65 ;
        RECT  1.14 2.75 115.52 2.85 ;
      VIA 87.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 2.8 via1_2_400_200_1_1_300_300 ;
    END
  END VDD
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  29.145 0 29.285 0.14 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 76.72 0.14 76.86 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  105.865 0 106.005 0.14 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 134.4 0.14 134.54 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 76.16 116.625 76.3 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  95.785 0 95.925 0.14 ;
    END
  END addr[5]
  PIN ce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  76.745 0 76.885 0.14 ;
    END
  END ce
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 95.76 0.14 95.9 ;
    END
  END clk
  PIN di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 124.88 0.14 125.02 ;
    END
  END di[0]
  PIN di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 28.56 116.625 28.7 ;
    END
  END di[10]
  PIN di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  72.825 139.41 72.965 139.55 ;
    END
  END di[11]
  PIN di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 19.04 116.625 19.18 ;
    END
  END di[12]
  PIN di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  91.865 139.41 92.005 139.55 ;
    END
  END di[13]
  PIN di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 38.08 116.625 38.22 ;
    END
  END di[14]
  PIN di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  5.625 139.41 5.765 139.55 ;
    END
  END di[15]
  PIN di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 47.6 116.625 47.74 ;
    END
  END di[16]
  PIN di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 86.24 0.14 86.38 ;
    END
  END di[17]
  PIN di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 124.32 116.625 124.46 ;
    END
  END di[18]
  PIN di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 38.64 0.14 38.78 ;
    END
  END di[19]
  PIN di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 57.68 0.14 57.82 ;
    END
  END di[1]
  PIN di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 105.84 0.14 105.98 ;
    END
  END di[20]
  PIN di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 9.52 116.625 9.66 ;
    END
  END di[21]
  PIN di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 67.2 0.14 67.34 ;
    END
  END di[2]
  PIN di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 105.28 116.625 105.42 ;
    END
  END di[3]
  PIN di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 19.6 0.14 19.74 ;
    END
  END di[4]
  PIN di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  62.745 139.41 62.885 139.55 ;
    END
  END di[5]
  PIN di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 29.12 0.14 29.26 ;
    END
  END di[6]
  PIN di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 133.84 116.625 133.98 ;
    END
  END di[7]
  PIN di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  43.705 139.41 43.845 139.55 ;
    END
  END di[8]
  PIN di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 85.68 116.625 85.82 ;
    END
  END di[9]
  PIN doq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  82.345 139.41 82.485 139.55 ;
    END
  END doq[0]
  PIN doq[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  10.105 0 10.245 0.14 ;
    END
  END doq[10]
  PIN doq[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END doq[11]
  PIN doq[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  24.665 139.41 24.805 139.55 ;
    END
  END doq[12]
  PIN doq[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 114.8 116.625 114.94 ;
    END
  END doq[13]
  PIN doq[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  48.185 0 48.325 0.14 ;
    END
  END doq[14]
  PIN doq[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 95.76 116.625 95.9 ;
    END
  END doq[15]
  PIN doq[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  115.385 0 115.525 0.14 ;
    END
  END doq[16]
  PIN doq[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  53.225 139.41 53.365 139.55 ;
    END
  END doq[17]
  PIN doq[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 57.12 116.625 57.26 ;
    END
  END doq[18]
  PIN doq[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  19.625 0 19.765 0.14 ;
    END
  END doq[19]
  PIN doq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  38.665 0 38.805 0.14 ;
    END
  END doq[1]
  PIN doq[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  57.705 0 57.845 0.14 ;
    END
  END doq[20]
  PIN doq[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 10.08 0.14 10.22 ;
    END
  END doq[21]
  PIN doq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  67.225 0 67.365 0.14 ;
    END
  END doq[2]
  PIN doq[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  110.905 139.41 111.045 139.55 ;
    END
  END doq[3]
  PIN doq[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  101.385 139.41 101.525 139.55 ;
    END
  END doq[4]
  PIN doq[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  15.145 139.41 15.285 139.55 ;
    END
  END doq[5]
  PIN doq[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  34.185 139.41 34.325 139.55 ;
    END
  END doq[6]
  PIN doq[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  86.265 0 86.405 0.14 ;
    END
  END doq[7]
  PIN doq[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 48.16 0.14 48.3 ;
    END
  END doq[8]
  PIN doq[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 115.36 0.14 115.5 ;
    END
  END doq[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  116.485 66.64 116.625 66.78 ;
    END
  END we
  OBS
    LAYER metal1 ;
     RECT  0 0 116.625 139.55 ;
    LAYER metal2 ;
     RECT  0 0 116.625 139.55 ;
    LAYER metal3 ;
     RECT  0 0 116.625 139.55 ;
    LAYER metal4 ;
     RECT  0 0 116.625 139.55 ;
    LAYER metal5 ;
     RECT  0 0 116.625 139.55 ;
    LAYER metal6 ;
     RECT  0 0 116.625 139.55 ;
    LAYER metal7 ;
     RECT  0 0 116.625 139.55 ;
  END
END or1200_spram3
END LIBRARY
