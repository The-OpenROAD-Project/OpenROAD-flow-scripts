VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_256x34
  FOREIGN fakeram45_256x34 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 98.420 BY 65.800 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.400 0.070 1.470 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.820 0.070 1.890 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.240 0.070 2.310 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.660 0.070 2.730 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.080 0.070 3.150 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.500 0.070 3.570 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.920 0.070 3.990 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.340 0.070 4.410 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.760 0.070 4.830 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.180 0.070 5.250 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.600 0.070 5.670 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.020 0.070 6.090 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.440 0.070 6.510 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.860 0.070 6.930 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.280 0.070 7.350 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.700 0.070 7.770 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.120 0.070 8.190 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.540 0.070 8.610 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.960 0.070 9.030 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.380 0.070 9.450 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.800 0.070 9.870 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.220 0.070 10.290 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.640 0.070 10.710 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.060 0.070 11.130 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.480 0.070 11.550 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.900 0.070 11.970 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.320 0.070 12.390 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.740 0.070 12.810 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.160 0.070 13.230 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.580 0.070 13.650 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.000 0.070 14.070 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.420 0.070 14.490 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.840 0.070 14.910 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.260 0.070 15.330 ;
    END
  END w_mask_in[33]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.040 0.070 19.110 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.460 0.070 19.530 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.880 0.070 19.950 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.300 0.070 20.370 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.720 0.070 20.790 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.140 0.070 21.210 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.560 0.070 21.630 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.980 0.070 22.050 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.400 0.070 22.470 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.820 0.070 22.890 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.240 0.070 23.310 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.660 0.070 23.730 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.080 0.070 24.150 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.500 0.070 24.570 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.920 0.070 24.990 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.340 0.070 25.410 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.760 0.070 25.830 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.180 0.070 26.250 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.600 0.070 26.670 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.020 0.070 27.090 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.440 0.070 27.510 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.860 0.070 27.930 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.280 0.070 28.350 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.700 0.070 28.770 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.120 0.070 29.190 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.540 0.070 29.610 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.960 0.070 30.030 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.380 0.070 30.450 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.800 0.070 30.870 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.220 0.070 31.290 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.640 0.070 31.710 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.060 0.070 32.130 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.480 0.070 32.550 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.900 0.070 32.970 ;
    END
  END rd_out[33]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.680 0.070 36.750 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.100 0.070 37.170 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.520 0.070 37.590 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.940 0.070 38.010 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.360 0.070 38.430 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.780 0.070 38.850 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.200 0.070 39.270 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.620 0.070 39.690 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.040 0.070 40.110 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.460 0.070 40.530 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.880 0.070 40.950 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.300 0.070 41.370 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.720 0.070 41.790 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.140 0.070 42.210 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.560 0.070 42.630 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.980 0.070 43.050 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.400 0.070 43.470 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.820 0.070 43.890 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.240 0.070 44.310 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.660 0.070 44.730 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.080 0.070 45.150 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.500 0.070 45.570 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.920 0.070 45.990 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.340 0.070 46.410 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.760 0.070 46.830 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.180 0.070 47.250 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.600 0.070 47.670 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.020 0.070 48.090 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.440 0.070 48.510 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.860 0.070 48.930 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.280 0.070 49.350 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.700 0.070 49.770 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.120 0.070 50.190 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.540 0.070 50.610 ;
    END
  END wd_in[33]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.320 0.070 54.390 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.740 0.070 54.810 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.160 0.070 55.230 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.580 0.070 55.650 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.000 0.070 56.070 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.420 0.070 56.490 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.840 0.070 56.910 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.260 0.070 57.330 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.040 0.070 61.110 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.460 0.070 61.530 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.880 0.070 61.950 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 64.400 ;
      RECT 3.500 1.400 3.780 64.400 ;
      RECT 5.740 1.400 6.020 64.400 ;
      RECT 7.980 1.400 8.260 64.400 ;
      RECT 10.220 1.400 10.500 64.400 ;
      RECT 12.460 1.400 12.740 64.400 ;
      RECT 14.700 1.400 14.980 64.400 ;
      RECT 16.940 1.400 17.220 64.400 ;
      RECT 19.180 1.400 19.460 64.400 ;
      RECT 21.420 1.400 21.700 64.400 ;
      RECT 23.660 1.400 23.940 64.400 ;
      RECT 25.900 1.400 26.180 64.400 ;
      RECT 28.140 1.400 28.420 64.400 ;
      RECT 30.380 1.400 30.660 64.400 ;
      RECT 32.620 1.400 32.900 64.400 ;
      RECT 34.860 1.400 35.140 64.400 ;
      RECT 37.100 1.400 37.380 64.400 ;
      RECT 39.340 1.400 39.620 64.400 ;
      RECT 41.580 1.400 41.860 64.400 ;
      RECT 43.820 1.400 44.100 64.400 ;
      RECT 46.060 1.400 46.340 64.400 ;
      RECT 48.300 1.400 48.580 64.400 ;
      RECT 50.540 1.400 50.820 64.400 ;
      RECT 52.780 1.400 53.060 64.400 ;
      RECT 55.020 1.400 55.300 64.400 ;
      RECT 57.260 1.400 57.540 64.400 ;
      RECT 59.500 1.400 59.780 64.400 ;
      RECT 61.740 1.400 62.020 64.400 ;
      RECT 63.980 1.400 64.260 64.400 ;
      RECT 66.220 1.400 66.500 64.400 ;
      RECT 68.460 1.400 68.740 64.400 ;
      RECT 70.700 1.400 70.980 64.400 ;
      RECT 72.940 1.400 73.220 64.400 ;
      RECT 75.180 1.400 75.460 64.400 ;
      RECT 77.420 1.400 77.700 64.400 ;
      RECT 79.660 1.400 79.940 64.400 ;
      RECT 81.900 1.400 82.180 64.400 ;
      RECT 84.140 1.400 84.420 64.400 ;
      RECT 86.380 1.400 86.660 64.400 ;
      RECT 88.620 1.400 88.900 64.400 ;
      RECT 90.860 1.400 91.140 64.400 ;
      RECT 93.100 1.400 93.380 64.400 ;
      RECT 95.340 1.400 95.620 64.400 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 64.400 ;
      RECT 4.620 1.400 4.900 64.400 ;
      RECT 6.860 1.400 7.140 64.400 ;
      RECT 9.100 1.400 9.380 64.400 ;
      RECT 11.340 1.400 11.620 64.400 ;
      RECT 13.580 1.400 13.860 64.400 ;
      RECT 15.820 1.400 16.100 64.400 ;
      RECT 18.060 1.400 18.340 64.400 ;
      RECT 20.300 1.400 20.580 64.400 ;
      RECT 22.540 1.400 22.820 64.400 ;
      RECT 24.780 1.400 25.060 64.400 ;
      RECT 27.020 1.400 27.300 64.400 ;
      RECT 29.260 1.400 29.540 64.400 ;
      RECT 31.500 1.400 31.780 64.400 ;
      RECT 33.740 1.400 34.020 64.400 ;
      RECT 35.980 1.400 36.260 64.400 ;
      RECT 38.220 1.400 38.500 64.400 ;
      RECT 40.460 1.400 40.740 64.400 ;
      RECT 42.700 1.400 42.980 64.400 ;
      RECT 44.940 1.400 45.220 64.400 ;
      RECT 47.180 1.400 47.460 64.400 ;
      RECT 49.420 1.400 49.700 64.400 ;
      RECT 51.660 1.400 51.940 64.400 ;
      RECT 53.900 1.400 54.180 64.400 ;
      RECT 56.140 1.400 56.420 64.400 ;
      RECT 58.380 1.400 58.660 64.400 ;
      RECT 60.620 1.400 60.900 64.400 ;
      RECT 62.860 1.400 63.140 64.400 ;
      RECT 65.100 1.400 65.380 64.400 ;
      RECT 67.340 1.400 67.620 64.400 ;
      RECT 69.580 1.400 69.860 64.400 ;
      RECT 71.820 1.400 72.100 64.400 ;
      RECT 74.060 1.400 74.340 64.400 ;
      RECT 76.300 1.400 76.580 64.400 ;
      RECT 78.540 1.400 78.820 64.400 ;
      RECT 80.780 1.400 81.060 64.400 ;
      RECT 83.020 1.400 83.300 64.400 ;
      RECT 85.260 1.400 85.540 64.400 ;
      RECT 87.500 1.400 87.780 64.400 ;
      RECT 89.740 1.400 90.020 64.400 ;
      RECT 91.980 1.400 92.260 64.400 ;
      RECT 94.220 1.400 94.500 64.400 ;
      RECT 96.460 1.400 96.740 64.400 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 98.420 65.800 ;
    LAYER metal2 ;
    RECT 0 0 98.420 65.800 ;
    LAYER metal3 ;
    RECT 0.070 0 98.420 65.800 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.785 ;
    RECT 0 1.855 0.070 2.205 ;
    RECT 0 2.275 0.070 2.625 ;
    RECT 0 2.695 0.070 3.045 ;
    RECT 0 3.115 0.070 3.465 ;
    RECT 0 3.535 0.070 3.885 ;
    RECT 0 3.955 0.070 4.305 ;
    RECT 0 4.375 0.070 4.725 ;
    RECT 0 4.795 0.070 5.145 ;
    RECT 0 5.215 0.070 5.565 ;
    RECT 0 5.635 0.070 5.985 ;
    RECT 0 6.055 0.070 6.405 ;
    RECT 0 6.475 0.070 6.825 ;
    RECT 0 6.895 0.070 7.245 ;
    RECT 0 7.315 0.070 7.665 ;
    RECT 0 7.735 0.070 8.085 ;
    RECT 0 8.155 0.070 8.505 ;
    RECT 0 8.575 0.070 8.925 ;
    RECT 0 8.995 0.070 9.345 ;
    RECT 0 9.415 0.070 9.765 ;
    RECT 0 9.835 0.070 10.185 ;
    RECT 0 10.255 0.070 10.605 ;
    RECT 0 10.675 0.070 11.025 ;
    RECT 0 11.095 0.070 11.445 ;
    RECT 0 11.515 0.070 11.865 ;
    RECT 0 11.935 0.070 12.285 ;
    RECT 0 12.355 0.070 12.705 ;
    RECT 0 12.775 0.070 13.125 ;
    RECT 0 13.195 0.070 13.545 ;
    RECT 0 13.615 0.070 13.965 ;
    RECT 0 14.035 0.070 14.385 ;
    RECT 0 14.455 0.070 14.805 ;
    RECT 0 14.875 0.070 15.225 ;
    RECT 0 15.295 0.070 19.005 ;
    RECT 0 19.075 0.070 19.425 ;
    RECT 0 19.495 0.070 19.845 ;
    RECT 0 19.915 0.070 20.265 ;
    RECT 0 20.335 0.070 20.685 ;
    RECT 0 20.755 0.070 21.105 ;
    RECT 0 21.175 0.070 21.525 ;
    RECT 0 21.595 0.070 21.945 ;
    RECT 0 22.015 0.070 22.365 ;
    RECT 0 22.435 0.070 22.785 ;
    RECT 0 22.855 0.070 23.205 ;
    RECT 0 23.275 0.070 23.625 ;
    RECT 0 23.695 0.070 24.045 ;
    RECT 0 24.115 0.070 24.465 ;
    RECT 0 24.535 0.070 24.885 ;
    RECT 0 24.955 0.070 25.305 ;
    RECT 0 25.375 0.070 25.725 ;
    RECT 0 25.795 0.070 26.145 ;
    RECT 0 26.215 0.070 26.565 ;
    RECT 0 26.635 0.070 26.985 ;
    RECT 0 27.055 0.070 27.405 ;
    RECT 0 27.475 0.070 27.825 ;
    RECT 0 27.895 0.070 28.245 ;
    RECT 0 28.315 0.070 28.665 ;
    RECT 0 28.735 0.070 29.085 ;
    RECT 0 29.155 0.070 29.505 ;
    RECT 0 29.575 0.070 29.925 ;
    RECT 0 29.995 0.070 30.345 ;
    RECT 0 30.415 0.070 30.765 ;
    RECT 0 30.835 0.070 31.185 ;
    RECT 0 31.255 0.070 31.605 ;
    RECT 0 31.675 0.070 32.025 ;
    RECT 0 32.095 0.070 32.445 ;
    RECT 0 32.515 0.070 32.865 ;
    RECT 0 32.935 0.070 36.645 ;
    RECT 0 36.715 0.070 37.065 ;
    RECT 0 37.135 0.070 37.485 ;
    RECT 0 37.555 0.070 37.905 ;
    RECT 0 37.975 0.070 38.325 ;
    RECT 0 38.395 0.070 38.745 ;
    RECT 0 38.815 0.070 39.165 ;
    RECT 0 39.235 0.070 39.585 ;
    RECT 0 39.655 0.070 40.005 ;
    RECT 0 40.075 0.070 40.425 ;
    RECT 0 40.495 0.070 40.845 ;
    RECT 0 40.915 0.070 41.265 ;
    RECT 0 41.335 0.070 41.685 ;
    RECT 0 41.755 0.070 42.105 ;
    RECT 0 42.175 0.070 42.525 ;
    RECT 0 42.595 0.070 42.945 ;
    RECT 0 43.015 0.070 43.365 ;
    RECT 0 43.435 0.070 43.785 ;
    RECT 0 43.855 0.070 44.205 ;
    RECT 0 44.275 0.070 44.625 ;
    RECT 0 44.695 0.070 45.045 ;
    RECT 0 45.115 0.070 45.465 ;
    RECT 0 45.535 0.070 45.885 ;
    RECT 0 45.955 0.070 46.305 ;
    RECT 0 46.375 0.070 46.725 ;
    RECT 0 46.795 0.070 47.145 ;
    RECT 0 47.215 0.070 47.565 ;
    RECT 0 47.635 0.070 47.985 ;
    RECT 0 48.055 0.070 48.405 ;
    RECT 0 48.475 0.070 48.825 ;
    RECT 0 48.895 0.070 49.245 ;
    RECT 0 49.315 0.070 49.665 ;
    RECT 0 49.735 0.070 50.085 ;
    RECT 0 50.155 0.070 50.505 ;
    RECT 0 50.575 0.070 54.285 ;
    RECT 0 54.355 0.070 54.705 ;
    RECT 0 54.775 0.070 55.125 ;
    RECT 0 55.195 0.070 55.545 ;
    RECT 0 55.615 0.070 55.965 ;
    RECT 0 56.035 0.070 56.385 ;
    RECT 0 56.455 0.070 56.805 ;
    RECT 0 56.875 0.070 57.225 ;
    RECT 0 57.295 0.070 61.005 ;
    RECT 0 61.075 0.070 61.425 ;
    RECT 0 61.495 0.070 61.845 ;
    RECT 0 61.915 0.070 65.800 ;
    LAYER metal4 ;
    RECT 0 0 98.420 1.400 ;
    RECT 0 64.400 98.420 65.800 ;
    RECT 0.000 1.400 1.260 64.400 ;
    RECT 1.540 1.400 2.380 64.400 ;
    RECT 2.660 1.400 3.500 64.400 ;
    RECT 3.780 1.400 4.620 64.400 ;
    RECT 4.900 1.400 5.740 64.400 ;
    RECT 6.020 1.400 6.860 64.400 ;
    RECT 7.140 1.400 7.980 64.400 ;
    RECT 8.260 1.400 9.100 64.400 ;
    RECT 9.380 1.400 10.220 64.400 ;
    RECT 10.500 1.400 11.340 64.400 ;
    RECT 11.620 1.400 12.460 64.400 ;
    RECT 12.740 1.400 13.580 64.400 ;
    RECT 13.860 1.400 14.700 64.400 ;
    RECT 14.980 1.400 15.820 64.400 ;
    RECT 16.100 1.400 16.940 64.400 ;
    RECT 17.220 1.400 18.060 64.400 ;
    RECT 18.340 1.400 19.180 64.400 ;
    RECT 19.460 1.400 20.300 64.400 ;
    RECT 20.580 1.400 21.420 64.400 ;
    RECT 21.700 1.400 22.540 64.400 ;
    RECT 22.820 1.400 23.660 64.400 ;
    RECT 23.940 1.400 24.780 64.400 ;
    RECT 25.060 1.400 25.900 64.400 ;
    RECT 26.180 1.400 27.020 64.400 ;
    RECT 27.300 1.400 28.140 64.400 ;
    RECT 28.420 1.400 29.260 64.400 ;
    RECT 29.540 1.400 30.380 64.400 ;
    RECT 30.660 1.400 31.500 64.400 ;
    RECT 31.780 1.400 32.620 64.400 ;
    RECT 32.900 1.400 33.740 64.400 ;
    RECT 34.020 1.400 34.860 64.400 ;
    RECT 35.140 1.400 35.980 64.400 ;
    RECT 36.260 1.400 37.100 64.400 ;
    RECT 37.380 1.400 38.220 64.400 ;
    RECT 38.500 1.400 39.340 64.400 ;
    RECT 39.620 1.400 40.460 64.400 ;
    RECT 40.740 1.400 41.580 64.400 ;
    RECT 41.860 1.400 42.700 64.400 ;
    RECT 42.980 1.400 43.820 64.400 ;
    RECT 44.100 1.400 44.940 64.400 ;
    RECT 45.220 1.400 46.060 64.400 ;
    RECT 46.340 1.400 47.180 64.400 ;
    RECT 47.460 1.400 48.300 64.400 ;
    RECT 48.580 1.400 49.420 64.400 ;
    RECT 49.700 1.400 50.540 64.400 ;
    RECT 50.820 1.400 51.660 64.400 ;
    RECT 51.940 1.400 52.780 64.400 ;
    RECT 53.060 1.400 53.900 64.400 ;
    RECT 54.180 1.400 55.020 64.400 ;
    RECT 55.300 1.400 56.140 64.400 ;
    RECT 56.420 1.400 57.260 64.400 ;
    RECT 57.540 1.400 58.380 64.400 ;
    RECT 58.660 1.400 59.500 64.400 ;
    RECT 59.780 1.400 60.620 64.400 ;
    RECT 60.900 1.400 61.740 64.400 ;
    RECT 62.020 1.400 62.860 64.400 ;
    RECT 63.140 1.400 63.980 64.400 ;
    RECT 64.260 1.400 65.100 64.400 ;
    RECT 65.380 1.400 66.220 64.400 ;
    RECT 66.500 1.400 67.340 64.400 ;
    RECT 67.620 1.400 68.460 64.400 ;
    RECT 68.740 1.400 69.580 64.400 ;
    RECT 69.860 1.400 70.700 64.400 ;
    RECT 70.980 1.400 71.820 64.400 ;
    RECT 72.100 1.400 72.940 64.400 ;
    RECT 73.220 1.400 74.060 64.400 ;
    RECT 74.340 1.400 75.180 64.400 ;
    RECT 75.460 1.400 76.300 64.400 ;
    RECT 76.580 1.400 77.420 64.400 ;
    RECT 77.700 1.400 78.540 64.400 ;
    RECT 78.820 1.400 79.660 64.400 ;
    RECT 79.940 1.400 80.780 64.400 ;
    RECT 81.060 1.400 81.900 64.400 ;
    RECT 82.180 1.400 83.020 64.400 ;
    RECT 83.300 1.400 84.140 64.400 ;
    RECT 84.420 1.400 85.260 64.400 ;
    RECT 85.540 1.400 86.380 64.400 ;
    RECT 86.660 1.400 87.500 64.400 ;
    RECT 87.780 1.400 88.620 64.400 ;
    RECT 88.900 1.400 89.740 64.400 ;
    RECT 90.020 1.400 90.860 64.400 ;
    RECT 91.140 1.400 91.980 64.400 ;
    RECT 92.260 1.400 93.100 64.400 ;
    RECT 93.380 1.400 94.220 64.400 ;
    RECT 94.500 1.400 95.340 64.400 ;
    RECT 95.620 1.400 96.460 64.400 ;
    RECT 96.740 1.400 98.420 64.400 ;
    LAYER OVERLAP ;
    RECT 0 0 98.420 65.800 ;
  END
END fakeram45_256x34

END LIBRARY
