VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_256x32
  FOREIGN fakeram45_256x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 60.610 BY 169.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.535 0.070 3.605 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.475 0.070 6.545 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.945 0.070 8.015 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.355 0.070 12.425 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.825 0.070 13.895 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.295 0.070 15.365 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.235 0.070 18.305 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.705 0.070 19.775 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.175 0.070 21.245 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.585 0.070 25.655 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.055 0.070 27.125 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.525 0.070 28.595 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.995 0.070 30.065 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.465 0.070 31.535 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.935 0.070 33.005 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.405 0.070 34.475 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.875 0.070 35.945 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.815 0.070 38.885 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.285 0.070 40.355 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.755 0.070 41.825 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.695 0.070 44.765 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.165 0.070 46.235 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.635 0.070 47.705 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.525 0.070 49.595 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.995 0.070 51.065 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.935 0.070 54.005 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.405 0.070 55.475 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.875 0.070 56.945 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.815 0.070 59.885 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.285 0.070 61.355 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.755 0.070 62.825 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 64.225 0.070 64.295 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 65.695 0.070 65.765 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 67.165 0.070 67.235 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 68.635 0.070 68.705 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.105 0.070 70.175 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.575 0.070 71.645 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.515 0.070 74.585 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.985 0.070 76.055 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.455 0.070 77.525 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.395 0.070 80.465 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.865 0.070 81.935 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.335 0.070 83.405 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.275 0.070 86.345 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.745 0.070 87.815 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.215 0.070 89.285 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.155 0.070 92.225 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.625 0.070 93.695 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.095 0.070 95.165 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.985 0.070 97.055 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 98.455 0.070 98.525 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 99.925 0.070 99.995 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 101.395 0.070 101.465 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 102.865 0.070 102.935 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 104.335 0.070 104.405 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.805 0.070 105.875 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.275 0.070 107.345 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 108.745 0.070 108.815 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 110.215 0.070 110.285 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 111.685 0.070 111.755 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 113.155 0.070 113.225 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 114.625 0.070 114.695 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 116.095 0.070 116.165 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 117.565 0.070 117.635 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 119.035 0.070 119.105 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 120.505 0.070 120.575 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 121.975 0.070 122.045 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 123.445 0.070 123.515 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 124.915 0.070 124.985 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 126.385 0.070 126.455 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 127.855 0.070 127.925 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 129.325 0.070 129.395 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 130.795 0.070 130.865 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 132.265 0.070 132.335 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 133.735 0.070 133.805 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 135.205 0.070 135.275 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 136.675 0.070 136.745 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 138.145 0.070 138.215 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 139.615 0.070 139.685 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 141.085 0.070 141.155 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 142.555 0.070 142.625 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 144.445 0.070 144.515 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 145.915 0.070 145.985 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 147.385 0.070 147.455 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 148.855 0.070 148.925 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 150.325 0.070 150.395 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 151.795 0.070 151.865 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 153.265 0.070 153.335 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 154.735 0.070 154.805 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 156.625 0.070 156.695 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 158.095 0.070 158.165 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 159.565 0.070 159.635 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 167.300 ;
      RECT 5.320 2.100 5.600 167.300 ;
      RECT 8.680 2.100 8.960 167.300 ;
      RECT 12.040 2.100 12.320 167.300 ;
      RECT 15.400 2.100 15.680 167.300 ;
      RECT 18.760 2.100 19.040 167.300 ;
      RECT 22.120 2.100 22.400 167.300 ;
      RECT 25.480 2.100 25.760 167.300 ;
      RECT 28.840 2.100 29.120 167.300 ;
      RECT 32.200 2.100 32.480 167.300 ;
      RECT 35.560 2.100 35.840 167.300 ;
      RECT 38.920 2.100 39.200 167.300 ;
      RECT 42.280 2.100 42.560 167.300 ;
      RECT 45.640 2.100 45.920 167.300 ;
      RECT 49.000 2.100 49.280 167.300 ;
      RECT 52.360 2.100 52.640 167.300 ;
      RECT 55.720 2.100 56.000 167.300 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 167.300 ;
      RECT 7.000 2.100 7.280 167.300 ;
      RECT 10.360 2.100 10.640 167.300 ;
      RECT 13.720 2.100 14.000 167.300 ;
      RECT 17.080 2.100 17.360 167.300 ;
      RECT 20.440 2.100 20.720 167.300 ;
      RECT 23.800 2.100 24.080 167.300 ;
      RECT 27.160 2.100 27.440 167.300 ;
      RECT 30.520 2.100 30.800 167.300 ;
      RECT 33.880 2.100 34.160 167.300 ;
      RECT 37.240 2.100 37.520 167.300 ;
      RECT 40.600 2.100 40.880 167.300 ;
      RECT 43.960 2.100 44.240 167.300 ;
      RECT 47.320 2.100 47.600 167.300 ;
      RECT 50.680 2.100 50.960 167.300 ;
      RECT 54.040 2.100 54.320 167.300 ;
      RECT 57.400 2.100 57.680 167.300 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 60.610 169.400 ;
    LAYER metal2 ;
    RECT 0 0 60.610 169.400 ;
    LAYER metal3 ;
    RECT 0.070 0 60.610 169.400 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 3.535 ;
    RECT 0 3.605 0.070 5.005 ;
    RECT 0 5.075 0.070 6.475 ;
    RECT 0 6.545 0.070 7.945 ;
    RECT 0 8.015 0.070 9.415 ;
    RECT 0 9.485 0.070 10.885 ;
    RECT 0 10.955 0.070 12.355 ;
    RECT 0 12.425 0.070 13.825 ;
    RECT 0 13.895 0.070 15.295 ;
    RECT 0 15.365 0.070 16.765 ;
    RECT 0 16.835 0.070 18.235 ;
    RECT 0 18.305 0.070 19.705 ;
    RECT 0 19.775 0.070 21.175 ;
    RECT 0 21.245 0.070 22.645 ;
    RECT 0 22.715 0.070 24.115 ;
    RECT 0 24.185 0.070 25.585 ;
    RECT 0 25.655 0.070 27.055 ;
    RECT 0 27.125 0.070 28.525 ;
    RECT 0 28.595 0.070 29.995 ;
    RECT 0 30.065 0.070 31.465 ;
    RECT 0 31.535 0.070 32.935 ;
    RECT 0 33.005 0.070 34.405 ;
    RECT 0 34.475 0.070 35.875 ;
    RECT 0 35.945 0.070 37.345 ;
    RECT 0 37.415 0.070 38.815 ;
    RECT 0 38.885 0.070 40.285 ;
    RECT 0 40.355 0.070 41.755 ;
    RECT 0 41.825 0.070 43.225 ;
    RECT 0 43.295 0.070 44.695 ;
    RECT 0 44.765 0.070 46.165 ;
    RECT 0 46.235 0.070 47.635 ;
    RECT 0 47.705 0.070 49.525 ;
    RECT 0 49.595 0.070 50.995 ;
    RECT 0 51.065 0.070 52.465 ;
    RECT 0 52.535 0.070 53.935 ;
    RECT 0 54.005 0.070 55.405 ;
    RECT 0 55.475 0.070 56.875 ;
    RECT 0 56.945 0.070 58.345 ;
    RECT 0 58.415 0.070 59.815 ;
    RECT 0 59.885 0.070 61.285 ;
    RECT 0 61.355 0.070 62.755 ;
    RECT 0 62.825 0.070 64.225 ;
    RECT 0 64.295 0.070 65.695 ;
    RECT 0 65.765 0.070 67.165 ;
    RECT 0 67.235 0.070 68.635 ;
    RECT 0 68.705 0.070 70.105 ;
    RECT 0 70.175 0.070 71.575 ;
    RECT 0 71.645 0.070 73.045 ;
    RECT 0 73.115 0.070 74.515 ;
    RECT 0 74.585 0.070 75.985 ;
    RECT 0 76.055 0.070 77.455 ;
    RECT 0 77.525 0.070 78.925 ;
    RECT 0 78.995 0.070 80.395 ;
    RECT 0 80.465 0.070 81.865 ;
    RECT 0 81.935 0.070 83.335 ;
    RECT 0 83.405 0.070 84.805 ;
    RECT 0 84.875 0.070 86.275 ;
    RECT 0 86.345 0.070 87.745 ;
    RECT 0 87.815 0.070 89.215 ;
    RECT 0 89.285 0.070 90.685 ;
    RECT 0 90.755 0.070 92.155 ;
    RECT 0 92.225 0.070 93.625 ;
    RECT 0 93.695 0.070 95.095 ;
    RECT 0 95.165 0.070 96.985 ;
    RECT 0 97.055 0.070 98.455 ;
    RECT 0 98.525 0.070 99.925 ;
    RECT 0 99.995 0.070 101.395 ;
    RECT 0 101.465 0.070 102.865 ;
    RECT 0 102.935 0.070 104.335 ;
    RECT 0 104.405 0.070 105.805 ;
    RECT 0 105.875 0.070 107.275 ;
    RECT 0 107.345 0.070 108.745 ;
    RECT 0 108.815 0.070 110.215 ;
    RECT 0 110.285 0.070 111.685 ;
    RECT 0 111.755 0.070 113.155 ;
    RECT 0 113.225 0.070 114.625 ;
    RECT 0 114.695 0.070 116.095 ;
    RECT 0 116.165 0.070 117.565 ;
    RECT 0 117.635 0.070 119.035 ;
    RECT 0 119.105 0.070 120.505 ;
    RECT 0 120.575 0.070 121.975 ;
    RECT 0 122.045 0.070 123.445 ;
    RECT 0 123.515 0.070 124.915 ;
    RECT 0 124.985 0.070 126.385 ;
    RECT 0 126.455 0.070 127.855 ;
    RECT 0 127.925 0.070 129.325 ;
    RECT 0 129.395 0.070 130.795 ;
    RECT 0 130.865 0.070 132.265 ;
    RECT 0 132.335 0.070 133.735 ;
    RECT 0 133.805 0.070 135.205 ;
    RECT 0 135.275 0.070 136.675 ;
    RECT 0 136.745 0.070 138.145 ;
    RECT 0 138.215 0.070 139.615 ;
    RECT 0 139.685 0.070 141.085 ;
    RECT 0 141.155 0.070 142.555 ;
    RECT 0 142.625 0.070 144.445 ;
    RECT 0 144.515 0.070 145.915 ;
    RECT 0 145.985 0.070 147.385 ;
    RECT 0 147.455 0.070 148.855 ;
    RECT 0 148.925 0.070 150.325 ;
    RECT 0 150.395 0.070 151.795 ;
    RECT 0 151.865 0.070 153.265 ;
    RECT 0 153.335 0.070 154.735 ;
    RECT 0 154.805 0.070 156.625 ;
    RECT 0 156.695 0.070 158.095 ;
    RECT 0 158.165 0.070 159.565 ;
    RECT 0 159.635 0.070 169.400 ;
    LAYER metal4 ;
    RECT 0 0 60.610 2.100 ;
    RECT 0 167.300 60.610 169.400 ;
    RECT 0.000 2.100 1.960 167.300 ;
    RECT 2.240 2.100 3.640 167.300 ;
    RECT 3.920 2.100 5.320 167.300 ;
    RECT 5.600 2.100 7.000 167.300 ;
    RECT 7.280 2.100 8.680 167.300 ;
    RECT 8.960 2.100 10.360 167.300 ;
    RECT 10.640 2.100 12.040 167.300 ;
    RECT 12.320 2.100 13.720 167.300 ;
    RECT 14.000 2.100 15.400 167.300 ;
    RECT 15.680 2.100 17.080 167.300 ;
    RECT 17.360 2.100 18.760 167.300 ;
    RECT 19.040 2.100 20.440 167.300 ;
    RECT 20.720 2.100 22.120 167.300 ;
    RECT 22.400 2.100 23.800 167.300 ;
    RECT 24.080 2.100 25.480 167.300 ;
    RECT 25.760 2.100 27.160 167.300 ;
    RECT 27.440 2.100 28.840 167.300 ;
    RECT 29.120 2.100 30.520 167.300 ;
    RECT 30.800 2.100 32.200 167.300 ;
    RECT 32.480 2.100 33.880 167.300 ;
    RECT 34.160 2.100 35.560 167.300 ;
    RECT 35.840 2.100 37.240 167.300 ;
    RECT 37.520 2.100 38.920 167.300 ;
    RECT 39.200 2.100 40.600 167.300 ;
    RECT 40.880 2.100 42.280 167.300 ;
    RECT 42.560 2.100 43.960 167.300 ;
    RECT 44.240 2.100 45.640 167.300 ;
    RECT 45.920 2.100 47.320 167.300 ;
    RECT 47.600 2.100 49.000 167.300 ;
    RECT 49.280 2.100 50.680 167.300 ;
    RECT 50.960 2.100 52.360 167.300 ;
    RECT 52.640 2.100 54.040 167.300 ;
    RECT 54.320 2.100 55.720 167.300 ;
    RECT 56.000 2.100 57.400 167.300 ;
    RECT 57.680 2.100 60.610 167.300 ;
    LAYER OVERLAP ;
    RECT 0 0 60.610 169.400 ;
  END
END fakeram45_256x32

END LIBRARY
