module MockArray(
  input        clock,
  input        reset,
  input  [7:0] io_insHorizontal_0_0,
  input  [7:0] io_insHorizontal_0_1,
  input  [7:0] io_insHorizontal_0_2,
  input  [7:0] io_insHorizontal_0_3,
  input  [7:0] io_insHorizontal_0_4,
  input  [7:0] io_insHorizontal_0_5,
  input  [7:0] io_insHorizontal_0_6,
  input  [7:0] io_insHorizontal_0_7,
  input  [7:0] io_insHorizontal_0_8,
  input  [7:0] io_insHorizontal_0_9,
  input  [7:0] io_insHorizontal_0_10,
  input  [7:0] io_insHorizontal_0_11,
  input  [7:0] io_insHorizontal_0_12,
  input  [7:0] io_insHorizontal_0_13,
  input  [7:0] io_insHorizontal_0_14,
  input  [7:0] io_insHorizontal_0_15,
  input  [7:0] io_insHorizontal_1_0,
  input  [7:0] io_insHorizontal_1_1,
  input  [7:0] io_insHorizontal_1_2,
  input  [7:0] io_insHorizontal_1_3,
  input  [7:0] io_insHorizontal_1_4,
  input  [7:0] io_insHorizontal_1_5,
  input  [7:0] io_insHorizontal_1_6,
  input  [7:0] io_insHorizontal_1_7,
  input  [7:0] io_insHorizontal_1_8,
  input  [7:0] io_insHorizontal_1_9,
  input  [7:0] io_insHorizontal_1_10,
  input  [7:0] io_insHorizontal_1_11,
  input  [7:0] io_insHorizontal_1_12,
  input  [7:0] io_insHorizontal_1_13,
  input  [7:0] io_insHorizontal_1_14,
  input  [7:0] io_insHorizontal_1_15,
  output [7:0] io_outsHorizontal_0_0,
  output [7:0] io_outsHorizontal_0_1,
  output [7:0] io_outsHorizontal_0_2,
  output [7:0] io_outsHorizontal_0_3,
  output [7:0] io_outsHorizontal_0_4,
  output [7:0] io_outsHorizontal_0_5,
  output [7:0] io_outsHorizontal_0_6,
  output [7:0] io_outsHorizontal_0_7,
  output [7:0] io_outsHorizontal_0_8,
  output [7:0] io_outsHorizontal_0_9,
  output [7:0] io_outsHorizontal_0_10,
  output [7:0] io_outsHorizontal_0_11,
  output [7:0] io_outsHorizontal_0_12,
  output [7:0] io_outsHorizontal_0_13,
  output [7:0] io_outsHorizontal_0_14,
  output [7:0] io_outsHorizontal_0_15,
  output [7:0] io_outsHorizontal_1_0,
  output [7:0] io_outsHorizontal_1_1,
  output [7:0] io_outsHorizontal_1_2,
  output [7:0] io_outsHorizontal_1_3,
  output [7:0] io_outsHorizontal_1_4,
  output [7:0] io_outsHorizontal_1_5,
  output [7:0] io_outsHorizontal_1_6,
  output [7:0] io_outsHorizontal_1_7,
  output [7:0] io_outsHorizontal_1_8,
  output [7:0] io_outsHorizontal_1_9,
  output [7:0] io_outsHorizontal_1_10,
  output [7:0] io_outsHorizontal_1_11,
  output [7:0] io_outsHorizontal_1_12,
  output [7:0] io_outsHorizontal_1_13,
  output [7:0] io_outsHorizontal_1_14,
  output [7:0] io_outsHorizontal_1_15,
  input  [7:0] io_insVertical_0_0,
  input  [7:0] io_insVertical_0_1,
  input  [7:0] io_insVertical_0_2,
  input  [7:0] io_insVertical_0_3,
  input  [7:0] io_insVertical_0_4,
  input  [7:0] io_insVertical_0_5,
  input  [7:0] io_insVertical_0_6,
  input  [7:0] io_insVertical_0_7,
  input  [7:0] io_insVertical_0_8,
  input  [7:0] io_insVertical_0_9,
  input  [7:0] io_insVertical_0_10,
  input  [7:0] io_insVertical_0_11,
  input  [7:0] io_insVertical_0_12,
  input  [7:0] io_insVertical_0_13,
  input  [7:0] io_insVertical_0_14,
  input  [7:0] io_insVertical_0_15,
  input  [7:0] io_insVertical_1_0,
  input  [7:0] io_insVertical_1_1,
  input  [7:0] io_insVertical_1_2,
  input  [7:0] io_insVertical_1_3,
  input  [7:0] io_insVertical_1_4,
  input  [7:0] io_insVertical_1_5,
  input  [7:0] io_insVertical_1_6,
  input  [7:0] io_insVertical_1_7,
  input  [7:0] io_insVertical_1_8,
  input  [7:0] io_insVertical_1_9,
  input  [7:0] io_insVertical_1_10,
  input  [7:0] io_insVertical_1_11,
  input  [7:0] io_insVertical_1_12,
  input  [7:0] io_insVertical_1_13,
  input  [7:0] io_insVertical_1_14,
  input  [7:0] io_insVertical_1_15,
  output [7:0] io_outsVertical_0_0,
  output [7:0] io_outsVertical_0_1,
  output [7:0] io_outsVertical_0_2,
  output [7:0] io_outsVertical_0_3,
  output [7:0] io_outsVertical_0_4,
  output [7:0] io_outsVertical_0_5,
  output [7:0] io_outsVertical_0_6,
  output [7:0] io_outsVertical_0_7,
  output [7:0] io_outsVertical_0_8,
  output [7:0] io_outsVertical_0_9,
  output [7:0] io_outsVertical_0_10,
  output [7:0] io_outsVertical_0_11,
  output [7:0] io_outsVertical_0_12,
  output [7:0] io_outsVertical_0_13,
  output [7:0] io_outsVertical_0_14,
  output [7:0] io_outsVertical_0_15,
  output [7:0] io_outsVertical_1_0,
  output [7:0] io_outsVertical_1_1,
  output [7:0] io_outsVertical_1_2,
  output [7:0] io_outsVertical_1_3,
  output [7:0] io_outsVertical_1_4,
  output [7:0] io_outsVertical_1_5,
  output [7:0] io_outsVertical_1_6,
  output [7:0] io_outsVertical_1_7,
  output [7:0] io_outsVertical_1_8,
  output [7:0] io_outsVertical_1_9,
  output [7:0] io_outsVertical_1_10,
  output [7:0] io_outsVertical_1_11,
  output [7:0] io_outsVertical_1_12,
  output [7:0] io_outsVertical_1_13,
  output [7:0] io_outsVertical_1_14,
  output [7:0] io_outsVertical_1_15
);
  wire  ces_0_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_0_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_0_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_1_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_1_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_2_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_2_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_3_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_3_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_4_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_4_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_5_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_5_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_6_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_6_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_7_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_7_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_8_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_8_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_9_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_9_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_10_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_10_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_11_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_11_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_12_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_12_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_13_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_13_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_14_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_14_15_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_0_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_0_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_0_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_0_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_0_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_0_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_0_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_0_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_0_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_1_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_1_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_1_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_1_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_1_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_1_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_1_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_1_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_1_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_2_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_2_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_2_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_2_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_2_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_2_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_2_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_2_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_2_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_3_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_3_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_3_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_3_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_3_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_3_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_3_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_3_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_3_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_4_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_4_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_4_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_4_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_4_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_4_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_4_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_4_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_4_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_5_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_5_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_5_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_5_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_5_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_5_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_5_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_5_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_5_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_6_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_6_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_6_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_6_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_6_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_6_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_6_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_6_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_6_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_7_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_7_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_7_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_7_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_7_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_7_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_7_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_7_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_7_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_8_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_8_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_8_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_8_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_8_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_8_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_8_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_8_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_8_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_9_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_9_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_9_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_9_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_9_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_9_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_9_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_9_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_9_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_10_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_10_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_10_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_10_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_10_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_10_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_10_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_10_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_10_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_11_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_11_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_11_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_11_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_11_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_11_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_11_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_11_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_11_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_12_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_12_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_12_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_12_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_12_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_12_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_12_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_12_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_12_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_13_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_13_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_13_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_13_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_13_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_13_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_13_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_13_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_13_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_14_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_14_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_14_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_14_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_14_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_14_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_14_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_14_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_14_io_outs_3; // @[MockArray.scala 37:53]
  wire  ces_15_15_clock; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_15_io_ins_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_15_io_ins_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_15_io_ins_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_15_io_ins_3; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_15_io_outs_0; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_15_io_outs_1; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_15_io_outs_2; // @[MockArray.scala 37:53]
  wire [7:0] ces_15_15_io_outs_3; // @[MockArray.scala 37:53]
  Element ces_0_0 ( // @[MockArray.scala 37:53]
    .clock(ces_0_0_clock),
    .io_ins_0(ces_0_0_io_ins_0),
    .io_ins_1(ces_0_0_io_ins_1),
    .io_ins_2(ces_0_0_io_ins_2),
    .io_ins_3(ces_0_0_io_ins_3),
    .io_outs_0(ces_0_0_io_outs_0),
    .io_outs_1(ces_0_0_io_outs_1),
    .io_outs_2(ces_0_0_io_outs_2),
    .io_outs_3(ces_0_0_io_outs_3)
  );
  Element ces_0_1 ( // @[MockArray.scala 37:53]
    .clock(ces_0_1_clock),
    .io_ins_0(ces_0_1_io_ins_0),
    .io_ins_1(ces_0_1_io_ins_1),
    .io_ins_2(ces_0_1_io_ins_2),
    .io_ins_3(ces_0_1_io_ins_3),
    .io_outs_0(ces_0_1_io_outs_0),
    .io_outs_1(ces_0_1_io_outs_1),
    .io_outs_2(ces_0_1_io_outs_2),
    .io_outs_3(ces_0_1_io_outs_3)
  );
  Element ces_0_2 ( // @[MockArray.scala 37:53]
    .clock(ces_0_2_clock),
    .io_ins_0(ces_0_2_io_ins_0),
    .io_ins_1(ces_0_2_io_ins_1),
    .io_ins_2(ces_0_2_io_ins_2),
    .io_ins_3(ces_0_2_io_ins_3),
    .io_outs_0(ces_0_2_io_outs_0),
    .io_outs_1(ces_0_2_io_outs_1),
    .io_outs_2(ces_0_2_io_outs_2),
    .io_outs_3(ces_0_2_io_outs_3)
  );
  Element ces_0_3 ( // @[MockArray.scala 37:53]
    .clock(ces_0_3_clock),
    .io_ins_0(ces_0_3_io_ins_0),
    .io_ins_1(ces_0_3_io_ins_1),
    .io_ins_2(ces_0_3_io_ins_2),
    .io_ins_3(ces_0_3_io_ins_3),
    .io_outs_0(ces_0_3_io_outs_0),
    .io_outs_1(ces_0_3_io_outs_1),
    .io_outs_2(ces_0_3_io_outs_2),
    .io_outs_3(ces_0_3_io_outs_3)
  );
  Element ces_0_4 ( // @[MockArray.scala 37:53]
    .clock(ces_0_4_clock),
    .io_ins_0(ces_0_4_io_ins_0),
    .io_ins_1(ces_0_4_io_ins_1),
    .io_ins_2(ces_0_4_io_ins_2),
    .io_ins_3(ces_0_4_io_ins_3),
    .io_outs_0(ces_0_4_io_outs_0),
    .io_outs_1(ces_0_4_io_outs_1),
    .io_outs_2(ces_0_4_io_outs_2),
    .io_outs_3(ces_0_4_io_outs_3)
  );
  Element ces_0_5 ( // @[MockArray.scala 37:53]
    .clock(ces_0_5_clock),
    .io_ins_0(ces_0_5_io_ins_0),
    .io_ins_1(ces_0_5_io_ins_1),
    .io_ins_2(ces_0_5_io_ins_2),
    .io_ins_3(ces_0_5_io_ins_3),
    .io_outs_0(ces_0_5_io_outs_0),
    .io_outs_1(ces_0_5_io_outs_1),
    .io_outs_2(ces_0_5_io_outs_2),
    .io_outs_3(ces_0_5_io_outs_3)
  );
  Element ces_0_6 ( // @[MockArray.scala 37:53]
    .clock(ces_0_6_clock),
    .io_ins_0(ces_0_6_io_ins_0),
    .io_ins_1(ces_0_6_io_ins_1),
    .io_ins_2(ces_0_6_io_ins_2),
    .io_ins_3(ces_0_6_io_ins_3),
    .io_outs_0(ces_0_6_io_outs_0),
    .io_outs_1(ces_0_6_io_outs_1),
    .io_outs_2(ces_0_6_io_outs_2),
    .io_outs_3(ces_0_6_io_outs_3)
  );
  Element ces_0_7 ( // @[MockArray.scala 37:53]
    .clock(ces_0_7_clock),
    .io_ins_0(ces_0_7_io_ins_0),
    .io_ins_1(ces_0_7_io_ins_1),
    .io_ins_2(ces_0_7_io_ins_2),
    .io_ins_3(ces_0_7_io_ins_3),
    .io_outs_0(ces_0_7_io_outs_0),
    .io_outs_1(ces_0_7_io_outs_1),
    .io_outs_2(ces_0_7_io_outs_2),
    .io_outs_3(ces_0_7_io_outs_3)
  );
  Element ces_0_8 ( // @[MockArray.scala 37:53]
    .clock(ces_0_8_clock),
    .io_ins_0(ces_0_8_io_ins_0),
    .io_ins_1(ces_0_8_io_ins_1),
    .io_ins_2(ces_0_8_io_ins_2),
    .io_ins_3(ces_0_8_io_ins_3),
    .io_outs_0(ces_0_8_io_outs_0),
    .io_outs_1(ces_0_8_io_outs_1),
    .io_outs_2(ces_0_8_io_outs_2),
    .io_outs_3(ces_0_8_io_outs_3)
  );
  Element ces_0_9 ( // @[MockArray.scala 37:53]
    .clock(ces_0_9_clock),
    .io_ins_0(ces_0_9_io_ins_0),
    .io_ins_1(ces_0_9_io_ins_1),
    .io_ins_2(ces_0_9_io_ins_2),
    .io_ins_3(ces_0_9_io_ins_3),
    .io_outs_0(ces_0_9_io_outs_0),
    .io_outs_1(ces_0_9_io_outs_1),
    .io_outs_2(ces_0_9_io_outs_2),
    .io_outs_3(ces_0_9_io_outs_3)
  );
  Element ces_0_10 ( // @[MockArray.scala 37:53]
    .clock(ces_0_10_clock),
    .io_ins_0(ces_0_10_io_ins_0),
    .io_ins_1(ces_0_10_io_ins_1),
    .io_ins_2(ces_0_10_io_ins_2),
    .io_ins_3(ces_0_10_io_ins_3),
    .io_outs_0(ces_0_10_io_outs_0),
    .io_outs_1(ces_0_10_io_outs_1),
    .io_outs_2(ces_0_10_io_outs_2),
    .io_outs_3(ces_0_10_io_outs_3)
  );
  Element ces_0_11 ( // @[MockArray.scala 37:53]
    .clock(ces_0_11_clock),
    .io_ins_0(ces_0_11_io_ins_0),
    .io_ins_1(ces_0_11_io_ins_1),
    .io_ins_2(ces_0_11_io_ins_2),
    .io_ins_3(ces_0_11_io_ins_3),
    .io_outs_0(ces_0_11_io_outs_0),
    .io_outs_1(ces_0_11_io_outs_1),
    .io_outs_2(ces_0_11_io_outs_2),
    .io_outs_3(ces_0_11_io_outs_3)
  );
  Element ces_0_12 ( // @[MockArray.scala 37:53]
    .clock(ces_0_12_clock),
    .io_ins_0(ces_0_12_io_ins_0),
    .io_ins_1(ces_0_12_io_ins_1),
    .io_ins_2(ces_0_12_io_ins_2),
    .io_ins_3(ces_0_12_io_ins_3),
    .io_outs_0(ces_0_12_io_outs_0),
    .io_outs_1(ces_0_12_io_outs_1),
    .io_outs_2(ces_0_12_io_outs_2),
    .io_outs_3(ces_0_12_io_outs_3)
  );
  Element ces_0_13 ( // @[MockArray.scala 37:53]
    .clock(ces_0_13_clock),
    .io_ins_0(ces_0_13_io_ins_0),
    .io_ins_1(ces_0_13_io_ins_1),
    .io_ins_2(ces_0_13_io_ins_2),
    .io_ins_3(ces_0_13_io_ins_3),
    .io_outs_0(ces_0_13_io_outs_0),
    .io_outs_1(ces_0_13_io_outs_1),
    .io_outs_2(ces_0_13_io_outs_2),
    .io_outs_3(ces_0_13_io_outs_3)
  );
  Element ces_0_14 ( // @[MockArray.scala 37:53]
    .clock(ces_0_14_clock),
    .io_ins_0(ces_0_14_io_ins_0),
    .io_ins_1(ces_0_14_io_ins_1),
    .io_ins_2(ces_0_14_io_ins_2),
    .io_ins_3(ces_0_14_io_ins_3),
    .io_outs_0(ces_0_14_io_outs_0),
    .io_outs_1(ces_0_14_io_outs_1),
    .io_outs_2(ces_0_14_io_outs_2),
    .io_outs_3(ces_0_14_io_outs_3)
  );
  Element ces_0_15 ( // @[MockArray.scala 37:53]
    .clock(ces_0_15_clock),
    .io_ins_0(ces_0_15_io_ins_0),
    .io_ins_1(ces_0_15_io_ins_1),
    .io_ins_2(ces_0_15_io_ins_2),
    .io_ins_3(ces_0_15_io_ins_3),
    .io_outs_0(ces_0_15_io_outs_0),
    .io_outs_1(ces_0_15_io_outs_1),
    .io_outs_2(ces_0_15_io_outs_2),
    .io_outs_3(ces_0_15_io_outs_3)
  );
  Element ces_1_0 ( // @[MockArray.scala 37:53]
    .clock(ces_1_0_clock),
    .io_ins_0(ces_1_0_io_ins_0),
    .io_ins_1(ces_1_0_io_ins_1),
    .io_ins_2(ces_1_0_io_ins_2),
    .io_ins_3(ces_1_0_io_ins_3),
    .io_outs_0(ces_1_0_io_outs_0),
    .io_outs_1(ces_1_0_io_outs_1),
    .io_outs_2(ces_1_0_io_outs_2),
    .io_outs_3(ces_1_0_io_outs_3)
  );
  Element ces_1_1 ( // @[MockArray.scala 37:53]
    .clock(ces_1_1_clock),
    .io_ins_0(ces_1_1_io_ins_0),
    .io_ins_1(ces_1_1_io_ins_1),
    .io_ins_2(ces_1_1_io_ins_2),
    .io_ins_3(ces_1_1_io_ins_3),
    .io_outs_0(ces_1_1_io_outs_0),
    .io_outs_1(ces_1_1_io_outs_1),
    .io_outs_2(ces_1_1_io_outs_2),
    .io_outs_3(ces_1_1_io_outs_3)
  );
  Element ces_1_2 ( // @[MockArray.scala 37:53]
    .clock(ces_1_2_clock),
    .io_ins_0(ces_1_2_io_ins_0),
    .io_ins_1(ces_1_2_io_ins_1),
    .io_ins_2(ces_1_2_io_ins_2),
    .io_ins_3(ces_1_2_io_ins_3),
    .io_outs_0(ces_1_2_io_outs_0),
    .io_outs_1(ces_1_2_io_outs_1),
    .io_outs_2(ces_1_2_io_outs_2),
    .io_outs_3(ces_1_2_io_outs_3)
  );
  Element ces_1_3 ( // @[MockArray.scala 37:53]
    .clock(ces_1_3_clock),
    .io_ins_0(ces_1_3_io_ins_0),
    .io_ins_1(ces_1_3_io_ins_1),
    .io_ins_2(ces_1_3_io_ins_2),
    .io_ins_3(ces_1_3_io_ins_3),
    .io_outs_0(ces_1_3_io_outs_0),
    .io_outs_1(ces_1_3_io_outs_1),
    .io_outs_2(ces_1_3_io_outs_2),
    .io_outs_3(ces_1_3_io_outs_3)
  );
  Element ces_1_4 ( // @[MockArray.scala 37:53]
    .clock(ces_1_4_clock),
    .io_ins_0(ces_1_4_io_ins_0),
    .io_ins_1(ces_1_4_io_ins_1),
    .io_ins_2(ces_1_4_io_ins_2),
    .io_ins_3(ces_1_4_io_ins_3),
    .io_outs_0(ces_1_4_io_outs_0),
    .io_outs_1(ces_1_4_io_outs_1),
    .io_outs_2(ces_1_4_io_outs_2),
    .io_outs_3(ces_1_4_io_outs_3)
  );
  Element ces_1_5 ( // @[MockArray.scala 37:53]
    .clock(ces_1_5_clock),
    .io_ins_0(ces_1_5_io_ins_0),
    .io_ins_1(ces_1_5_io_ins_1),
    .io_ins_2(ces_1_5_io_ins_2),
    .io_ins_3(ces_1_5_io_ins_3),
    .io_outs_0(ces_1_5_io_outs_0),
    .io_outs_1(ces_1_5_io_outs_1),
    .io_outs_2(ces_1_5_io_outs_2),
    .io_outs_3(ces_1_5_io_outs_3)
  );
  Element ces_1_6 ( // @[MockArray.scala 37:53]
    .clock(ces_1_6_clock),
    .io_ins_0(ces_1_6_io_ins_0),
    .io_ins_1(ces_1_6_io_ins_1),
    .io_ins_2(ces_1_6_io_ins_2),
    .io_ins_3(ces_1_6_io_ins_3),
    .io_outs_0(ces_1_6_io_outs_0),
    .io_outs_1(ces_1_6_io_outs_1),
    .io_outs_2(ces_1_6_io_outs_2),
    .io_outs_3(ces_1_6_io_outs_3)
  );
  Element ces_1_7 ( // @[MockArray.scala 37:53]
    .clock(ces_1_7_clock),
    .io_ins_0(ces_1_7_io_ins_0),
    .io_ins_1(ces_1_7_io_ins_1),
    .io_ins_2(ces_1_7_io_ins_2),
    .io_ins_3(ces_1_7_io_ins_3),
    .io_outs_0(ces_1_7_io_outs_0),
    .io_outs_1(ces_1_7_io_outs_1),
    .io_outs_2(ces_1_7_io_outs_2),
    .io_outs_3(ces_1_7_io_outs_3)
  );
  Element ces_1_8 ( // @[MockArray.scala 37:53]
    .clock(ces_1_8_clock),
    .io_ins_0(ces_1_8_io_ins_0),
    .io_ins_1(ces_1_8_io_ins_1),
    .io_ins_2(ces_1_8_io_ins_2),
    .io_ins_3(ces_1_8_io_ins_3),
    .io_outs_0(ces_1_8_io_outs_0),
    .io_outs_1(ces_1_8_io_outs_1),
    .io_outs_2(ces_1_8_io_outs_2),
    .io_outs_3(ces_1_8_io_outs_3)
  );
  Element ces_1_9 ( // @[MockArray.scala 37:53]
    .clock(ces_1_9_clock),
    .io_ins_0(ces_1_9_io_ins_0),
    .io_ins_1(ces_1_9_io_ins_1),
    .io_ins_2(ces_1_9_io_ins_2),
    .io_ins_3(ces_1_9_io_ins_3),
    .io_outs_0(ces_1_9_io_outs_0),
    .io_outs_1(ces_1_9_io_outs_1),
    .io_outs_2(ces_1_9_io_outs_2),
    .io_outs_3(ces_1_9_io_outs_3)
  );
  Element ces_1_10 ( // @[MockArray.scala 37:53]
    .clock(ces_1_10_clock),
    .io_ins_0(ces_1_10_io_ins_0),
    .io_ins_1(ces_1_10_io_ins_1),
    .io_ins_2(ces_1_10_io_ins_2),
    .io_ins_3(ces_1_10_io_ins_3),
    .io_outs_0(ces_1_10_io_outs_0),
    .io_outs_1(ces_1_10_io_outs_1),
    .io_outs_2(ces_1_10_io_outs_2),
    .io_outs_3(ces_1_10_io_outs_3)
  );
  Element ces_1_11 ( // @[MockArray.scala 37:53]
    .clock(ces_1_11_clock),
    .io_ins_0(ces_1_11_io_ins_0),
    .io_ins_1(ces_1_11_io_ins_1),
    .io_ins_2(ces_1_11_io_ins_2),
    .io_ins_3(ces_1_11_io_ins_3),
    .io_outs_0(ces_1_11_io_outs_0),
    .io_outs_1(ces_1_11_io_outs_1),
    .io_outs_2(ces_1_11_io_outs_2),
    .io_outs_3(ces_1_11_io_outs_3)
  );
  Element ces_1_12 ( // @[MockArray.scala 37:53]
    .clock(ces_1_12_clock),
    .io_ins_0(ces_1_12_io_ins_0),
    .io_ins_1(ces_1_12_io_ins_1),
    .io_ins_2(ces_1_12_io_ins_2),
    .io_ins_3(ces_1_12_io_ins_3),
    .io_outs_0(ces_1_12_io_outs_0),
    .io_outs_1(ces_1_12_io_outs_1),
    .io_outs_2(ces_1_12_io_outs_2),
    .io_outs_3(ces_1_12_io_outs_3)
  );
  Element ces_1_13 ( // @[MockArray.scala 37:53]
    .clock(ces_1_13_clock),
    .io_ins_0(ces_1_13_io_ins_0),
    .io_ins_1(ces_1_13_io_ins_1),
    .io_ins_2(ces_1_13_io_ins_2),
    .io_ins_3(ces_1_13_io_ins_3),
    .io_outs_0(ces_1_13_io_outs_0),
    .io_outs_1(ces_1_13_io_outs_1),
    .io_outs_2(ces_1_13_io_outs_2),
    .io_outs_3(ces_1_13_io_outs_3)
  );
  Element ces_1_14 ( // @[MockArray.scala 37:53]
    .clock(ces_1_14_clock),
    .io_ins_0(ces_1_14_io_ins_0),
    .io_ins_1(ces_1_14_io_ins_1),
    .io_ins_2(ces_1_14_io_ins_2),
    .io_ins_3(ces_1_14_io_ins_3),
    .io_outs_0(ces_1_14_io_outs_0),
    .io_outs_1(ces_1_14_io_outs_1),
    .io_outs_2(ces_1_14_io_outs_2),
    .io_outs_3(ces_1_14_io_outs_3)
  );
  Element ces_1_15 ( // @[MockArray.scala 37:53]
    .clock(ces_1_15_clock),
    .io_ins_0(ces_1_15_io_ins_0),
    .io_ins_1(ces_1_15_io_ins_1),
    .io_ins_2(ces_1_15_io_ins_2),
    .io_ins_3(ces_1_15_io_ins_3),
    .io_outs_0(ces_1_15_io_outs_0),
    .io_outs_1(ces_1_15_io_outs_1),
    .io_outs_2(ces_1_15_io_outs_2),
    .io_outs_3(ces_1_15_io_outs_3)
  );
  Element ces_2_0 ( // @[MockArray.scala 37:53]
    .clock(ces_2_0_clock),
    .io_ins_0(ces_2_0_io_ins_0),
    .io_ins_1(ces_2_0_io_ins_1),
    .io_ins_2(ces_2_0_io_ins_2),
    .io_ins_3(ces_2_0_io_ins_3),
    .io_outs_0(ces_2_0_io_outs_0),
    .io_outs_1(ces_2_0_io_outs_1),
    .io_outs_2(ces_2_0_io_outs_2),
    .io_outs_3(ces_2_0_io_outs_3)
  );
  Element ces_2_1 ( // @[MockArray.scala 37:53]
    .clock(ces_2_1_clock),
    .io_ins_0(ces_2_1_io_ins_0),
    .io_ins_1(ces_2_1_io_ins_1),
    .io_ins_2(ces_2_1_io_ins_2),
    .io_ins_3(ces_2_1_io_ins_3),
    .io_outs_0(ces_2_1_io_outs_0),
    .io_outs_1(ces_2_1_io_outs_1),
    .io_outs_2(ces_2_1_io_outs_2),
    .io_outs_3(ces_2_1_io_outs_3)
  );
  Element ces_2_2 ( // @[MockArray.scala 37:53]
    .clock(ces_2_2_clock),
    .io_ins_0(ces_2_2_io_ins_0),
    .io_ins_1(ces_2_2_io_ins_1),
    .io_ins_2(ces_2_2_io_ins_2),
    .io_ins_3(ces_2_2_io_ins_3),
    .io_outs_0(ces_2_2_io_outs_0),
    .io_outs_1(ces_2_2_io_outs_1),
    .io_outs_2(ces_2_2_io_outs_2),
    .io_outs_3(ces_2_2_io_outs_3)
  );
  Element ces_2_3 ( // @[MockArray.scala 37:53]
    .clock(ces_2_3_clock),
    .io_ins_0(ces_2_3_io_ins_0),
    .io_ins_1(ces_2_3_io_ins_1),
    .io_ins_2(ces_2_3_io_ins_2),
    .io_ins_3(ces_2_3_io_ins_3),
    .io_outs_0(ces_2_3_io_outs_0),
    .io_outs_1(ces_2_3_io_outs_1),
    .io_outs_2(ces_2_3_io_outs_2),
    .io_outs_3(ces_2_3_io_outs_3)
  );
  Element ces_2_4 ( // @[MockArray.scala 37:53]
    .clock(ces_2_4_clock),
    .io_ins_0(ces_2_4_io_ins_0),
    .io_ins_1(ces_2_4_io_ins_1),
    .io_ins_2(ces_2_4_io_ins_2),
    .io_ins_3(ces_2_4_io_ins_3),
    .io_outs_0(ces_2_4_io_outs_0),
    .io_outs_1(ces_2_4_io_outs_1),
    .io_outs_2(ces_2_4_io_outs_2),
    .io_outs_3(ces_2_4_io_outs_3)
  );
  Element ces_2_5 ( // @[MockArray.scala 37:53]
    .clock(ces_2_5_clock),
    .io_ins_0(ces_2_5_io_ins_0),
    .io_ins_1(ces_2_5_io_ins_1),
    .io_ins_2(ces_2_5_io_ins_2),
    .io_ins_3(ces_2_5_io_ins_3),
    .io_outs_0(ces_2_5_io_outs_0),
    .io_outs_1(ces_2_5_io_outs_1),
    .io_outs_2(ces_2_5_io_outs_2),
    .io_outs_3(ces_2_5_io_outs_3)
  );
  Element ces_2_6 ( // @[MockArray.scala 37:53]
    .clock(ces_2_6_clock),
    .io_ins_0(ces_2_6_io_ins_0),
    .io_ins_1(ces_2_6_io_ins_1),
    .io_ins_2(ces_2_6_io_ins_2),
    .io_ins_3(ces_2_6_io_ins_3),
    .io_outs_0(ces_2_6_io_outs_0),
    .io_outs_1(ces_2_6_io_outs_1),
    .io_outs_2(ces_2_6_io_outs_2),
    .io_outs_3(ces_2_6_io_outs_3)
  );
  Element ces_2_7 ( // @[MockArray.scala 37:53]
    .clock(ces_2_7_clock),
    .io_ins_0(ces_2_7_io_ins_0),
    .io_ins_1(ces_2_7_io_ins_1),
    .io_ins_2(ces_2_7_io_ins_2),
    .io_ins_3(ces_2_7_io_ins_3),
    .io_outs_0(ces_2_7_io_outs_0),
    .io_outs_1(ces_2_7_io_outs_1),
    .io_outs_2(ces_2_7_io_outs_2),
    .io_outs_3(ces_2_7_io_outs_3)
  );
  Element ces_2_8 ( // @[MockArray.scala 37:53]
    .clock(ces_2_8_clock),
    .io_ins_0(ces_2_8_io_ins_0),
    .io_ins_1(ces_2_8_io_ins_1),
    .io_ins_2(ces_2_8_io_ins_2),
    .io_ins_3(ces_2_8_io_ins_3),
    .io_outs_0(ces_2_8_io_outs_0),
    .io_outs_1(ces_2_8_io_outs_1),
    .io_outs_2(ces_2_8_io_outs_2),
    .io_outs_3(ces_2_8_io_outs_3)
  );
  Element ces_2_9 ( // @[MockArray.scala 37:53]
    .clock(ces_2_9_clock),
    .io_ins_0(ces_2_9_io_ins_0),
    .io_ins_1(ces_2_9_io_ins_1),
    .io_ins_2(ces_2_9_io_ins_2),
    .io_ins_3(ces_2_9_io_ins_3),
    .io_outs_0(ces_2_9_io_outs_0),
    .io_outs_1(ces_2_9_io_outs_1),
    .io_outs_2(ces_2_9_io_outs_2),
    .io_outs_3(ces_2_9_io_outs_3)
  );
  Element ces_2_10 ( // @[MockArray.scala 37:53]
    .clock(ces_2_10_clock),
    .io_ins_0(ces_2_10_io_ins_0),
    .io_ins_1(ces_2_10_io_ins_1),
    .io_ins_2(ces_2_10_io_ins_2),
    .io_ins_3(ces_2_10_io_ins_3),
    .io_outs_0(ces_2_10_io_outs_0),
    .io_outs_1(ces_2_10_io_outs_1),
    .io_outs_2(ces_2_10_io_outs_2),
    .io_outs_3(ces_2_10_io_outs_3)
  );
  Element ces_2_11 ( // @[MockArray.scala 37:53]
    .clock(ces_2_11_clock),
    .io_ins_0(ces_2_11_io_ins_0),
    .io_ins_1(ces_2_11_io_ins_1),
    .io_ins_2(ces_2_11_io_ins_2),
    .io_ins_3(ces_2_11_io_ins_3),
    .io_outs_0(ces_2_11_io_outs_0),
    .io_outs_1(ces_2_11_io_outs_1),
    .io_outs_2(ces_2_11_io_outs_2),
    .io_outs_3(ces_2_11_io_outs_3)
  );
  Element ces_2_12 ( // @[MockArray.scala 37:53]
    .clock(ces_2_12_clock),
    .io_ins_0(ces_2_12_io_ins_0),
    .io_ins_1(ces_2_12_io_ins_1),
    .io_ins_2(ces_2_12_io_ins_2),
    .io_ins_3(ces_2_12_io_ins_3),
    .io_outs_0(ces_2_12_io_outs_0),
    .io_outs_1(ces_2_12_io_outs_1),
    .io_outs_2(ces_2_12_io_outs_2),
    .io_outs_3(ces_2_12_io_outs_3)
  );
  Element ces_2_13 ( // @[MockArray.scala 37:53]
    .clock(ces_2_13_clock),
    .io_ins_0(ces_2_13_io_ins_0),
    .io_ins_1(ces_2_13_io_ins_1),
    .io_ins_2(ces_2_13_io_ins_2),
    .io_ins_3(ces_2_13_io_ins_3),
    .io_outs_0(ces_2_13_io_outs_0),
    .io_outs_1(ces_2_13_io_outs_1),
    .io_outs_2(ces_2_13_io_outs_2),
    .io_outs_3(ces_2_13_io_outs_3)
  );
  Element ces_2_14 ( // @[MockArray.scala 37:53]
    .clock(ces_2_14_clock),
    .io_ins_0(ces_2_14_io_ins_0),
    .io_ins_1(ces_2_14_io_ins_1),
    .io_ins_2(ces_2_14_io_ins_2),
    .io_ins_3(ces_2_14_io_ins_3),
    .io_outs_0(ces_2_14_io_outs_0),
    .io_outs_1(ces_2_14_io_outs_1),
    .io_outs_2(ces_2_14_io_outs_2),
    .io_outs_3(ces_2_14_io_outs_3)
  );
  Element ces_2_15 ( // @[MockArray.scala 37:53]
    .clock(ces_2_15_clock),
    .io_ins_0(ces_2_15_io_ins_0),
    .io_ins_1(ces_2_15_io_ins_1),
    .io_ins_2(ces_2_15_io_ins_2),
    .io_ins_3(ces_2_15_io_ins_3),
    .io_outs_0(ces_2_15_io_outs_0),
    .io_outs_1(ces_2_15_io_outs_1),
    .io_outs_2(ces_2_15_io_outs_2),
    .io_outs_3(ces_2_15_io_outs_3)
  );
  Element ces_3_0 ( // @[MockArray.scala 37:53]
    .clock(ces_3_0_clock),
    .io_ins_0(ces_3_0_io_ins_0),
    .io_ins_1(ces_3_0_io_ins_1),
    .io_ins_2(ces_3_0_io_ins_2),
    .io_ins_3(ces_3_0_io_ins_3),
    .io_outs_0(ces_3_0_io_outs_0),
    .io_outs_1(ces_3_0_io_outs_1),
    .io_outs_2(ces_3_0_io_outs_2),
    .io_outs_3(ces_3_0_io_outs_3)
  );
  Element ces_3_1 ( // @[MockArray.scala 37:53]
    .clock(ces_3_1_clock),
    .io_ins_0(ces_3_1_io_ins_0),
    .io_ins_1(ces_3_1_io_ins_1),
    .io_ins_2(ces_3_1_io_ins_2),
    .io_ins_3(ces_3_1_io_ins_3),
    .io_outs_0(ces_3_1_io_outs_0),
    .io_outs_1(ces_3_1_io_outs_1),
    .io_outs_2(ces_3_1_io_outs_2),
    .io_outs_3(ces_3_1_io_outs_3)
  );
  Element ces_3_2 ( // @[MockArray.scala 37:53]
    .clock(ces_3_2_clock),
    .io_ins_0(ces_3_2_io_ins_0),
    .io_ins_1(ces_3_2_io_ins_1),
    .io_ins_2(ces_3_2_io_ins_2),
    .io_ins_3(ces_3_2_io_ins_3),
    .io_outs_0(ces_3_2_io_outs_0),
    .io_outs_1(ces_3_2_io_outs_1),
    .io_outs_2(ces_3_2_io_outs_2),
    .io_outs_3(ces_3_2_io_outs_3)
  );
  Element ces_3_3 ( // @[MockArray.scala 37:53]
    .clock(ces_3_3_clock),
    .io_ins_0(ces_3_3_io_ins_0),
    .io_ins_1(ces_3_3_io_ins_1),
    .io_ins_2(ces_3_3_io_ins_2),
    .io_ins_3(ces_3_3_io_ins_3),
    .io_outs_0(ces_3_3_io_outs_0),
    .io_outs_1(ces_3_3_io_outs_1),
    .io_outs_2(ces_3_3_io_outs_2),
    .io_outs_3(ces_3_3_io_outs_3)
  );
  Element ces_3_4 ( // @[MockArray.scala 37:53]
    .clock(ces_3_4_clock),
    .io_ins_0(ces_3_4_io_ins_0),
    .io_ins_1(ces_3_4_io_ins_1),
    .io_ins_2(ces_3_4_io_ins_2),
    .io_ins_3(ces_3_4_io_ins_3),
    .io_outs_0(ces_3_4_io_outs_0),
    .io_outs_1(ces_3_4_io_outs_1),
    .io_outs_2(ces_3_4_io_outs_2),
    .io_outs_3(ces_3_4_io_outs_3)
  );
  Element ces_3_5 ( // @[MockArray.scala 37:53]
    .clock(ces_3_5_clock),
    .io_ins_0(ces_3_5_io_ins_0),
    .io_ins_1(ces_3_5_io_ins_1),
    .io_ins_2(ces_3_5_io_ins_2),
    .io_ins_3(ces_3_5_io_ins_3),
    .io_outs_0(ces_3_5_io_outs_0),
    .io_outs_1(ces_3_5_io_outs_1),
    .io_outs_2(ces_3_5_io_outs_2),
    .io_outs_3(ces_3_5_io_outs_3)
  );
  Element ces_3_6 ( // @[MockArray.scala 37:53]
    .clock(ces_3_6_clock),
    .io_ins_0(ces_3_6_io_ins_0),
    .io_ins_1(ces_3_6_io_ins_1),
    .io_ins_2(ces_3_6_io_ins_2),
    .io_ins_3(ces_3_6_io_ins_3),
    .io_outs_0(ces_3_6_io_outs_0),
    .io_outs_1(ces_3_6_io_outs_1),
    .io_outs_2(ces_3_6_io_outs_2),
    .io_outs_3(ces_3_6_io_outs_3)
  );
  Element ces_3_7 ( // @[MockArray.scala 37:53]
    .clock(ces_3_7_clock),
    .io_ins_0(ces_3_7_io_ins_0),
    .io_ins_1(ces_3_7_io_ins_1),
    .io_ins_2(ces_3_7_io_ins_2),
    .io_ins_3(ces_3_7_io_ins_3),
    .io_outs_0(ces_3_7_io_outs_0),
    .io_outs_1(ces_3_7_io_outs_1),
    .io_outs_2(ces_3_7_io_outs_2),
    .io_outs_3(ces_3_7_io_outs_3)
  );
  Element ces_3_8 ( // @[MockArray.scala 37:53]
    .clock(ces_3_8_clock),
    .io_ins_0(ces_3_8_io_ins_0),
    .io_ins_1(ces_3_8_io_ins_1),
    .io_ins_2(ces_3_8_io_ins_2),
    .io_ins_3(ces_3_8_io_ins_3),
    .io_outs_0(ces_3_8_io_outs_0),
    .io_outs_1(ces_3_8_io_outs_1),
    .io_outs_2(ces_3_8_io_outs_2),
    .io_outs_3(ces_3_8_io_outs_3)
  );
  Element ces_3_9 ( // @[MockArray.scala 37:53]
    .clock(ces_3_9_clock),
    .io_ins_0(ces_3_9_io_ins_0),
    .io_ins_1(ces_3_9_io_ins_1),
    .io_ins_2(ces_3_9_io_ins_2),
    .io_ins_3(ces_3_9_io_ins_3),
    .io_outs_0(ces_3_9_io_outs_0),
    .io_outs_1(ces_3_9_io_outs_1),
    .io_outs_2(ces_3_9_io_outs_2),
    .io_outs_3(ces_3_9_io_outs_3)
  );
  Element ces_3_10 ( // @[MockArray.scala 37:53]
    .clock(ces_3_10_clock),
    .io_ins_0(ces_3_10_io_ins_0),
    .io_ins_1(ces_3_10_io_ins_1),
    .io_ins_2(ces_3_10_io_ins_2),
    .io_ins_3(ces_3_10_io_ins_3),
    .io_outs_0(ces_3_10_io_outs_0),
    .io_outs_1(ces_3_10_io_outs_1),
    .io_outs_2(ces_3_10_io_outs_2),
    .io_outs_3(ces_3_10_io_outs_3)
  );
  Element ces_3_11 ( // @[MockArray.scala 37:53]
    .clock(ces_3_11_clock),
    .io_ins_0(ces_3_11_io_ins_0),
    .io_ins_1(ces_3_11_io_ins_1),
    .io_ins_2(ces_3_11_io_ins_2),
    .io_ins_3(ces_3_11_io_ins_3),
    .io_outs_0(ces_3_11_io_outs_0),
    .io_outs_1(ces_3_11_io_outs_1),
    .io_outs_2(ces_3_11_io_outs_2),
    .io_outs_3(ces_3_11_io_outs_3)
  );
  Element ces_3_12 ( // @[MockArray.scala 37:53]
    .clock(ces_3_12_clock),
    .io_ins_0(ces_3_12_io_ins_0),
    .io_ins_1(ces_3_12_io_ins_1),
    .io_ins_2(ces_3_12_io_ins_2),
    .io_ins_3(ces_3_12_io_ins_3),
    .io_outs_0(ces_3_12_io_outs_0),
    .io_outs_1(ces_3_12_io_outs_1),
    .io_outs_2(ces_3_12_io_outs_2),
    .io_outs_3(ces_3_12_io_outs_3)
  );
  Element ces_3_13 ( // @[MockArray.scala 37:53]
    .clock(ces_3_13_clock),
    .io_ins_0(ces_3_13_io_ins_0),
    .io_ins_1(ces_3_13_io_ins_1),
    .io_ins_2(ces_3_13_io_ins_2),
    .io_ins_3(ces_3_13_io_ins_3),
    .io_outs_0(ces_3_13_io_outs_0),
    .io_outs_1(ces_3_13_io_outs_1),
    .io_outs_2(ces_3_13_io_outs_2),
    .io_outs_3(ces_3_13_io_outs_3)
  );
  Element ces_3_14 ( // @[MockArray.scala 37:53]
    .clock(ces_3_14_clock),
    .io_ins_0(ces_3_14_io_ins_0),
    .io_ins_1(ces_3_14_io_ins_1),
    .io_ins_2(ces_3_14_io_ins_2),
    .io_ins_3(ces_3_14_io_ins_3),
    .io_outs_0(ces_3_14_io_outs_0),
    .io_outs_1(ces_3_14_io_outs_1),
    .io_outs_2(ces_3_14_io_outs_2),
    .io_outs_3(ces_3_14_io_outs_3)
  );
  Element ces_3_15 ( // @[MockArray.scala 37:53]
    .clock(ces_3_15_clock),
    .io_ins_0(ces_3_15_io_ins_0),
    .io_ins_1(ces_3_15_io_ins_1),
    .io_ins_2(ces_3_15_io_ins_2),
    .io_ins_3(ces_3_15_io_ins_3),
    .io_outs_0(ces_3_15_io_outs_0),
    .io_outs_1(ces_3_15_io_outs_1),
    .io_outs_2(ces_3_15_io_outs_2),
    .io_outs_3(ces_3_15_io_outs_3)
  );
  Element ces_4_0 ( // @[MockArray.scala 37:53]
    .clock(ces_4_0_clock),
    .io_ins_0(ces_4_0_io_ins_0),
    .io_ins_1(ces_4_0_io_ins_1),
    .io_ins_2(ces_4_0_io_ins_2),
    .io_ins_3(ces_4_0_io_ins_3),
    .io_outs_0(ces_4_0_io_outs_0),
    .io_outs_1(ces_4_0_io_outs_1),
    .io_outs_2(ces_4_0_io_outs_2),
    .io_outs_3(ces_4_0_io_outs_3)
  );
  Element ces_4_1 ( // @[MockArray.scala 37:53]
    .clock(ces_4_1_clock),
    .io_ins_0(ces_4_1_io_ins_0),
    .io_ins_1(ces_4_1_io_ins_1),
    .io_ins_2(ces_4_1_io_ins_2),
    .io_ins_3(ces_4_1_io_ins_3),
    .io_outs_0(ces_4_1_io_outs_0),
    .io_outs_1(ces_4_1_io_outs_1),
    .io_outs_2(ces_4_1_io_outs_2),
    .io_outs_3(ces_4_1_io_outs_3)
  );
  Element ces_4_2 ( // @[MockArray.scala 37:53]
    .clock(ces_4_2_clock),
    .io_ins_0(ces_4_2_io_ins_0),
    .io_ins_1(ces_4_2_io_ins_1),
    .io_ins_2(ces_4_2_io_ins_2),
    .io_ins_3(ces_4_2_io_ins_3),
    .io_outs_0(ces_4_2_io_outs_0),
    .io_outs_1(ces_4_2_io_outs_1),
    .io_outs_2(ces_4_2_io_outs_2),
    .io_outs_3(ces_4_2_io_outs_3)
  );
  Element ces_4_3 ( // @[MockArray.scala 37:53]
    .clock(ces_4_3_clock),
    .io_ins_0(ces_4_3_io_ins_0),
    .io_ins_1(ces_4_3_io_ins_1),
    .io_ins_2(ces_4_3_io_ins_2),
    .io_ins_3(ces_4_3_io_ins_3),
    .io_outs_0(ces_4_3_io_outs_0),
    .io_outs_1(ces_4_3_io_outs_1),
    .io_outs_2(ces_4_3_io_outs_2),
    .io_outs_3(ces_4_3_io_outs_3)
  );
  Element ces_4_4 ( // @[MockArray.scala 37:53]
    .clock(ces_4_4_clock),
    .io_ins_0(ces_4_4_io_ins_0),
    .io_ins_1(ces_4_4_io_ins_1),
    .io_ins_2(ces_4_4_io_ins_2),
    .io_ins_3(ces_4_4_io_ins_3),
    .io_outs_0(ces_4_4_io_outs_0),
    .io_outs_1(ces_4_4_io_outs_1),
    .io_outs_2(ces_4_4_io_outs_2),
    .io_outs_3(ces_4_4_io_outs_3)
  );
  Element ces_4_5 ( // @[MockArray.scala 37:53]
    .clock(ces_4_5_clock),
    .io_ins_0(ces_4_5_io_ins_0),
    .io_ins_1(ces_4_5_io_ins_1),
    .io_ins_2(ces_4_5_io_ins_2),
    .io_ins_3(ces_4_5_io_ins_3),
    .io_outs_0(ces_4_5_io_outs_0),
    .io_outs_1(ces_4_5_io_outs_1),
    .io_outs_2(ces_4_5_io_outs_2),
    .io_outs_3(ces_4_5_io_outs_3)
  );
  Element ces_4_6 ( // @[MockArray.scala 37:53]
    .clock(ces_4_6_clock),
    .io_ins_0(ces_4_6_io_ins_0),
    .io_ins_1(ces_4_6_io_ins_1),
    .io_ins_2(ces_4_6_io_ins_2),
    .io_ins_3(ces_4_6_io_ins_3),
    .io_outs_0(ces_4_6_io_outs_0),
    .io_outs_1(ces_4_6_io_outs_1),
    .io_outs_2(ces_4_6_io_outs_2),
    .io_outs_3(ces_4_6_io_outs_3)
  );
  Element ces_4_7 ( // @[MockArray.scala 37:53]
    .clock(ces_4_7_clock),
    .io_ins_0(ces_4_7_io_ins_0),
    .io_ins_1(ces_4_7_io_ins_1),
    .io_ins_2(ces_4_7_io_ins_2),
    .io_ins_3(ces_4_7_io_ins_3),
    .io_outs_0(ces_4_7_io_outs_0),
    .io_outs_1(ces_4_7_io_outs_1),
    .io_outs_2(ces_4_7_io_outs_2),
    .io_outs_3(ces_4_7_io_outs_3)
  );
  Element ces_4_8 ( // @[MockArray.scala 37:53]
    .clock(ces_4_8_clock),
    .io_ins_0(ces_4_8_io_ins_0),
    .io_ins_1(ces_4_8_io_ins_1),
    .io_ins_2(ces_4_8_io_ins_2),
    .io_ins_3(ces_4_8_io_ins_3),
    .io_outs_0(ces_4_8_io_outs_0),
    .io_outs_1(ces_4_8_io_outs_1),
    .io_outs_2(ces_4_8_io_outs_2),
    .io_outs_3(ces_4_8_io_outs_3)
  );
  Element ces_4_9 ( // @[MockArray.scala 37:53]
    .clock(ces_4_9_clock),
    .io_ins_0(ces_4_9_io_ins_0),
    .io_ins_1(ces_4_9_io_ins_1),
    .io_ins_2(ces_4_9_io_ins_2),
    .io_ins_3(ces_4_9_io_ins_3),
    .io_outs_0(ces_4_9_io_outs_0),
    .io_outs_1(ces_4_9_io_outs_1),
    .io_outs_2(ces_4_9_io_outs_2),
    .io_outs_3(ces_4_9_io_outs_3)
  );
  Element ces_4_10 ( // @[MockArray.scala 37:53]
    .clock(ces_4_10_clock),
    .io_ins_0(ces_4_10_io_ins_0),
    .io_ins_1(ces_4_10_io_ins_1),
    .io_ins_2(ces_4_10_io_ins_2),
    .io_ins_3(ces_4_10_io_ins_3),
    .io_outs_0(ces_4_10_io_outs_0),
    .io_outs_1(ces_4_10_io_outs_1),
    .io_outs_2(ces_4_10_io_outs_2),
    .io_outs_3(ces_4_10_io_outs_3)
  );
  Element ces_4_11 ( // @[MockArray.scala 37:53]
    .clock(ces_4_11_clock),
    .io_ins_0(ces_4_11_io_ins_0),
    .io_ins_1(ces_4_11_io_ins_1),
    .io_ins_2(ces_4_11_io_ins_2),
    .io_ins_3(ces_4_11_io_ins_3),
    .io_outs_0(ces_4_11_io_outs_0),
    .io_outs_1(ces_4_11_io_outs_1),
    .io_outs_2(ces_4_11_io_outs_2),
    .io_outs_3(ces_4_11_io_outs_3)
  );
  Element ces_4_12 ( // @[MockArray.scala 37:53]
    .clock(ces_4_12_clock),
    .io_ins_0(ces_4_12_io_ins_0),
    .io_ins_1(ces_4_12_io_ins_1),
    .io_ins_2(ces_4_12_io_ins_2),
    .io_ins_3(ces_4_12_io_ins_3),
    .io_outs_0(ces_4_12_io_outs_0),
    .io_outs_1(ces_4_12_io_outs_1),
    .io_outs_2(ces_4_12_io_outs_2),
    .io_outs_3(ces_4_12_io_outs_3)
  );
  Element ces_4_13 ( // @[MockArray.scala 37:53]
    .clock(ces_4_13_clock),
    .io_ins_0(ces_4_13_io_ins_0),
    .io_ins_1(ces_4_13_io_ins_1),
    .io_ins_2(ces_4_13_io_ins_2),
    .io_ins_3(ces_4_13_io_ins_3),
    .io_outs_0(ces_4_13_io_outs_0),
    .io_outs_1(ces_4_13_io_outs_1),
    .io_outs_2(ces_4_13_io_outs_2),
    .io_outs_3(ces_4_13_io_outs_3)
  );
  Element ces_4_14 ( // @[MockArray.scala 37:53]
    .clock(ces_4_14_clock),
    .io_ins_0(ces_4_14_io_ins_0),
    .io_ins_1(ces_4_14_io_ins_1),
    .io_ins_2(ces_4_14_io_ins_2),
    .io_ins_3(ces_4_14_io_ins_3),
    .io_outs_0(ces_4_14_io_outs_0),
    .io_outs_1(ces_4_14_io_outs_1),
    .io_outs_2(ces_4_14_io_outs_2),
    .io_outs_3(ces_4_14_io_outs_3)
  );
  Element ces_4_15 ( // @[MockArray.scala 37:53]
    .clock(ces_4_15_clock),
    .io_ins_0(ces_4_15_io_ins_0),
    .io_ins_1(ces_4_15_io_ins_1),
    .io_ins_2(ces_4_15_io_ins_2),
    .io_ins_3(ces_4_15_io_ins_3),
    .io_outs_0(ces_4_15_io_outs_0),
    .io_outs_1(ces_4_15_io_outs_1),
    .io_outs_2(ces_4_15_io_outs_2),
    .io_outs_3(ces_4_15_io_outs_3)
  );
  Element ces_5_0 ( // @[MockArray.scala 37:53]
    .clock(ces_5_0_clock),
    .io_ins_0(ces_5_0_io_ins_0),
    .io_ins_1(ces_5_0_io_ins_1),
    .io_ins_2(ces_5_0_io_ins_2),
    .io_ins_3(ces_5_0_io_ins_3),
    .io_outs_0(ces_5_0_io_outs_0),
    .io_outs_1(ces_5_0_io_outs_1),
    .io_outs_2(ces_5_0_io_outs_2),
    .io_outs_3(ces_5_0_io_outs_3)
  );
  Element ces_5_1 ( // @[MockArray.scala 37:53]
    .clock(ces_5_1_clock),
    .io_ins_0(ces_5_1_io_ins_0),
    .io_ins_1(ces_5_1_io_ins_1),
    .io_ins_2(ces_5_1_io_ins_2),
    .io_ins_3(ces_5_1_io_ins_3),
    .io_outs_0(ces_5_1_io_outs_0),
    .io_outs_1(ces_5_1_io_outs_1),
    .io_outs_2(ces_5_1_io_outs_2),
    .io_outs_3(ces_5_1_io_outs_3)
  );
  Element ces_5_2 ( // @[MockArray.scala 37:53]
    .clock(ces_5_2_clock),
    .io_ins_0(ces_5_2_io_ins_0),
    .io_ins_1(ces_5_2_io_ins_1),
    .io_ins_2(ces_5_2_io_ins_2),
    .io_ins_3(ces_5_2_io_ins_3),
    .io_outs_0(ces_5_2_io_outs_0),
    .io_outs_1(ces_5_2_io_outs_1),
    .io_outs_2(ces_5_2_io_outs_2),
    .io_outs_3(ces_5_2_io_outs_3)
  );
  Element ces_5_3 ( // @[MockArray.scala 37:53]
    .clock(ces_5_3_clock),
    .io_ins_0(ces_5_3_io_ins_0),
    .io_ins_1(ces_5_3_io_ins_1),
    .io_ins_2(ces_5_3_io_ins_2),
    .io_ins_3(ces_5_3_io_ins_3),
    .io_outs_0(ces_5_3_io_outs_0),
    .io_outs_1(ces_5_3_io_outs_1),
    .io_outs_2(ces_5_3_io_outs_2),
    .io_outs_3(ces_5_3_io_outs_3)
  );
  Element ces_5_4 ( // @[MockArray.scala 37:53]
    .clock(ces_5_4_clock),
    .io_ins_0(ces_5_4_io_ins_0),
    .io_ins_1(ces_5_4_io_ins_1),
    .io_ins_2(ces_5_4_io_ins_2),
    .io_ins_3(ces_5_4_io_ins_3),
    .io_outs_0(ces_5_4_io_outs_0),
    .io_outs_1(ces_5_4_io_outs_1),
    .io_outs_2(ces_5_4_io_outs_2),
    .io_outs_3(ces_5_4_io_outs_3)
  );
  Element ces_5_5 ( // @[MockArray.scala 37:53]
    .clock(ces_5_5_clock),
    .io_ins_0(ces_5_5_io_ins_0),
    .io_ins_1(ces_5_5_io_ins_1),
    .io_ins_2(ces_5_5_io_ins_2),
    .io_ins_3(ces_5_5_io_ins_3),
    .io_outs_0(ces_5_5_io_outs_0),
    .io_outs_1(ces_5_5_io_outs_1),
    .io_outs_2(ces_5_5_io_outs_2),
    .io_outs_3(ces_5_5_io_outs_3)
  );
  Element ces_5_6 ( // @[MockArray.scala 37:53]
    .clock(ces_5_6_clock),
    .io_ins_0(ces_5_6_io_ins_0),
    .io_ins_1(ces_5_6_io_ins_1),
    .io_ins_2(ces_5_6_io_ins_2),
    .io_ins_3(ces_5_6_io_ins_3),
    .io_outs_0(ces_5_6_io_outs_0),
    .io_outs_1(ces_5_6_io_outs_1),
    .io_outs_2(ces_5_6_io_outs_2),
    .io_outs_3(ces_5_6_io_outs_3)
  );
  Element ces_5_7 ( // @[MockArray.scala 37:53]
    .clock(ces_5_7_clock),
    .io_ins_0(ces_5_7_io_ins_0),
    .io_ins_1(ces_5_7_io_ins_1),
    .io_ins_2(ces_5_7_io_ins_2),
    .io_ins_3(ces_5_7_io_ins_3),
    .io_outs_0(ces_5_7_io_outs_0),
    .io_outs_1(ces_5_7_io_outs_1),
    .io_outs_2(ces_5_7_io_outs_2),
    .io_outs_3(ces_5_7_io_outs_3)
  );
  Element ces_5_8 ( // @[MockArray.scala 37:53]
    .clock(ces_5_8_clock),
    .io_ins_0(ces_5_8_io_ins_0),
    .io_ins_1(ces_5_8_io_ins_1),
    .io_ins_2(ces_5_8_io_ins_2),
    .io_ins_3(ces_5_8_io_ins_3),
    .io_outs_0(ces_5_8_io_outs_0),
    .io_outs_1(ces_5_8_io_outs_1),
    .io_outs_2(ces_5_8_io_outs_2),
    .io_outs_3(ces_5_8_io_outs_3)
  );
  Element ces_5_9 ( // @[MockArray.scala 37:53]
    .clock(ces_5_9_clock),
    .io_ins_0(ces_5_9_io_ins_0),
    .io_ins_1(ces_5_9_io_ins_1),
    .io_ins_2(ces_5_9_io_ins_2),
    .io_ins_3(ces_5_9_io_ins_3),
    .io_outs_0(ces_5_9_io_outs_0),
    .io_outs_1(ces_5_9_io_outs_1),
    .io_outs_2(ces_5_9_io_outs_2),
    .io_outs_3(ces_5_9_io_outs_3)
  );
  Element ces_5_10 ( // @[MockArray.scala 37:53]
    .clock(ces_5_10_clock),
    .io_ins_0(ces_5_10_io_ins_0),
    .io_ins_1(ces_5_10_io_ins_1),
    .io_ins_2(ces_5_10_io_ins_2),
    .io_ins_3(ces_5_10_io_ins_3),
    .io_outs_0(ces_5_10_io_outs_0),
    .io_outs_1(ces_5_10_io_outs_1),
    .io_outs_2(ces_5_10_io_outs_2),
    .io_outs_3(ces_5_10_io_outs_3)
  );
  Element ces_5_11 ( // @[MockArray.scala 37:53]
    .clock(ces_5_11_clock),
    .io_ins_0(ces_5_11_io_ins_0),
    .io_ins_1(ces_5_11_io_ins_1),
    .io_ins_2(ces_5_11_io_ins_2),
    .io_ins_3(ces_5_11_io_ins_3),
    .io_outs_0(ces_5_11_io_outs_0),
    .io_outs_1(ces_5_11_io_outs_1),
    .io_outs_2(ces_5_11_io_outs_2),
    .io_outs_3(ces_5_11_io_outs_3)
  );
  Element ces_5_12 ( // @[MockArray.scala 37:53]
    .clock(ces_5_12_clock),
    .io_ins_0(ces_5_12_io_ins_0),
    .io_ins_1(ces_5_12_io_ins_1),
    .io_ins_2(ces_5_12_io_ins_2),
    .io_ins_3(ces_5_12_io_ins_3),
    .io_outs_0(ces_5_12_io_outs_0),
    .io_outs_1(ces_5_12_io_outs_1),
    .io_outs_2(ces_5_12_io_outs_2),
    .io_outs_3(ces_5_12_io_outs_3)
  );
  Element ces_5_13 ( // @[MockArray.scala 37:53]
    .clock(ces_5_13_clock),
    .io_ins_0(ces_5_13_io_ins_0),
    .io_ins_1(ces_5_13_io_ins_1),
    .io_ins_2(ces_5_13_io_ins_2),
    .io_ins_3(ces_5_13_io_ins_3),
    .io_outs_0(ces_5_13_io_outs_0),
    .io_outs_1(ces_5_13_io_outs_1),
    .io_outs_2(ces_5_13_io_outs_2),
    .io_outs_3(ces_5_13_io_outs_3)
  );
  Element ces_5_14 ( // @[MockArray.scala 37:53]
    .clock(ces_5_14_clock),
    .io_ins_0(ces_5_14_io_ins_0),
    .io_ins_1(ces_5_14_io_ins_1),
    .io_ins_2(ces_5_14_io_ins_2),
    .io_ins_3(ces_5_14_io_ins_3),
    .io_outs_0(ces_5_14_io_outs_0),
    .io_outs_1(ces_5_14_io_outs_1),
    .io_outs_2(ces_5_14_io_outs_2),
    .io_outs_3(ces_5_14_io_outs_3)
  );
  Element ces_5_15 ( // @[MockArray.scala 37:53]
    .clock(ces_5_15_clock),
    .io_ins_0(ces_5_15_io_ins_0),
    .io_ins_1(ces_5_15_io_ins_1),
    .io_ins_2(ces_5_15_io_ins_2),
    .io_ins_3(ces_5_15_io_ins_3),
    .io_outs_0(ces_5_15_io_outs_0),
    .io_outs_1(ces_5_15_io_outs_1),
    .io_outs_2(ces_5_15_io_outs_2),
    .io_outs_3(ces_5_15_io_outs_3)
  );
  Element ces_6_0 ( // @[MockArray.scala 37:53]
    .clock(ces_6_0_clock),
    .io_ins_0(ces_6_0_io_ins_0),
    .io_ins_1(ces_6_0_io_ins_1),
    .io_ins_2(ces_6_0_io_ins_2),
    .io_ins_3(ces_6_0_io_ins_3),
    .io_outs_0(ces_6_0_io_outs_0),
    .io_outs_1(ces_6_0_io_outs_1),
    .io_outs_2(ces_6_0_io_outs_2),
    .io_outs_3(ces_6_0_io_outs_3)
  );
  Element ces_6_1 ( // @[MockArray.scala 37:53]
    .clock(ces_6_1_clock),
    .io_ins_0(ces_6_1_io_ins_0),
    .io_ins_1(ces_6_1_io_ins_1),
    .io_ins_2(ces_6_1_io_ins_2),
    .io_ins_3(ces_6_1_io_ins_3),
    .io_outs_0(ces_6_1_io_outs_0),
    .io_outs_1(ces_6_1_io_outs_1),
    .io_outs_2(ces_6_1_io_outs_2),
    .io_outs_3(ces_6_1_io_outs_3)
  );
  Element ces_6_2 ( // @[MockArray.scala 37:53]
    .clock(ces_6_2_clock),
    .io_ins_0(ces_6_2_io_ins_0),
    .io_ins_1(ces_6_2_io_ins_1),
    .io_ins_2(ces_6_2_io_ins_2),
    .io_ins_3(ces_6_2_io_ins_3),
    .io_outs_0(ces_6_2_io_outs_0),
    .io_outs_1(ces_6_2_io_outs_1),
    .io_outs_2(ces_6_2_io_outs_2),
    .io_outs_3(ces_6_2_io_outs_3)
  );
  Element ces_6_3 ( // @[MockArray.scala 37:53]
    .clock(ces_6_3_clock),
    .io_ins_0(ces_6_3_io_ins_0),
    .io_ins_1(ces_6_3_io_ins_1),
    .io_ins_2(ces_6_3_io_ins_2),
    .io_ins_3(ces_6_3_io_ins_3),
    .io_outs_0(ces_6_3_io_outs_0),
    .io_outs_1(ces_6_3_io_outs_1),
    .io_outs_2(ces_6_3_io_outs_2),
    .io_outs_3(ces_6_3_io_outs_3)
  );
  Element ces_6_4 ( // @[MockArray.scala 37:53]
    .clock(ces_6_4_clock),
    .io_ins_0(ces_6_4_io_ins_0),
    .io_ins_1(ces_6_4_io_ins_1),
    .io_ins_2(ces_6_4_io_ins_2),
    .io_ins_3(ces_6_4_io_ins_3),
    .io_outs_0(ces_6_4_io_outs_0),
    .io_outs_1(ces_6_4_io_outs_1),
    .io_outs_2(ces_6_4_io_outs_2),
    .io_outs_3(ces_6_4_io_outs_3)
  );
  Element ces_6_5 ( // @[MockArray.scala 37:53]
    .clock(ces_6_5_clock),
    .io_ins_0(ces_6_5_io_ins_0),
    .io_ins_1(ces_6_5_io_ins_1),
    .io_ins_2(ces_6_5_io_ins_2),
    .io_ins_3(ces_6_5_io_ins_3),
    .io_outs_0(ces_6_5_io_outs_0),
    .io_outs_1(ces_6_5_io_outs_1),
    .io_outs_2(ces_6_5_io_outs_2),
    .io_outs_3(ces_6_5_io_outs_3)
  );
  Element ces_6_6 ( // @[MockArray.scala 37:53]
    .clock(ces_6_6_clock),
    .io_ins_0(ces_6_6_io_ins_0),
    .io_ins_1(ces_6_6_io_ins_1),
    .io_ins_2(ces_6_6_io_ins_2),
    .io_ins_3(ces_6_6_io_ins_3),
    .io_outs_0(ces_6_6_io_outs_0),
    .io_outs_1(ces_6_6_io_outs_1),
    .io_outs_2(ces_6_6_io_outs_2),
    .io_outs_3(ces_6_6_io_outs_3)
  );
  Element ces_6_7 ( // @[MockArray.scala 37:53]
    .clock(ces_6_7_clock),
    .io_ins_0(ces_6_7_io_ins_0),
    .io_ins_1(ces_6_7_io_ins_1),
    .io_ins_2(ces_6_7_io_ins_2),
    .io_ins_3(ces_6_7_io_ins_3),
    .io_outs_0(ces_6_7_io_outs_0),
    .io_outs_1(ces_6_7_io_outs_1),
    .io_outs_2(ces_6_7_io_outs_2),
    .io_outs_3(ces_6_7_io_outs_3)
  );
  Element ces_6_8 ( // @[MockArray.scala 37:53]
    .clock(ces_6_8_clock),
    .io_ins_0(ces_6_8_io_ins_0),
    .io_ins_1(ces_6_8_io_ins_1),
    .io_ins_2(ces_6_8_io_ins_2),
    .io_ins_3(ces_6_8_io_ins_3),
    .io_outs_0(ces_6_8_io_outs_0),
    .io_outs_1(ces_6_8_io_outs_1),
    .io_outs_2(ces_6_8_io_outs_2),
    .io_outs_3(ces_6_8_io_outs_3)
  );
  Element ces_6_9 ( // @[MockArray.scala 37:53]
    .clock(ces_6_9_clock),
    .io_ins_0(ces_6_9_io_ins_0),
    .io_ins_1(ces_6_9_io_ins_1),
    .io_ins_2(ces_6_9_io_ins_2),
    .io_ins_3(ces_6_9_io_ins_3),
    .io_outs_0(ces_6_9_io_outs_0),
    .io_outs_1(ces_6_9_io_outs_1),
    .io_outs_2(ces_6_9_io_outs_2),
    .io_outs_3(ces_6_9_io_outs_3)
  );
  Element ces_6_10 ( // @[MockArray.scala 37:53]
    .clock(ces_6_10_clock),
    .io_ins_0(ces_6_10_io_ins_0),
    .io_ins_1(ces_6_10_io_ins_1),
    .io_ins_2(ces_6_10_io_ins_2),
    .io_ins_3(ces_6_10_io_ins_3),
    .io_outs_0(ces_6_10_io_outs_0),
    .io_outs_1(ces_6_10_io_outs_1),
    .io_outs_2(ces_6_10_io_outs_2),
    .io_outs_3(ces_6_10_io_outs_3)
  );
  Element ces_6_11 ( // @[MockArray.scala 37:53]
    .clock(ces_6_11_clock),
    .io_ins_0(ces_6_11_io_ins_0),
    .io_ins_1(ces_6_11_io_ins_1),
    .io_ins_2(ces_6_11_io_ins_2),
    .io_ins_3(ces_6_11_io_ins_3),
    .io_outs_0(ces_6_11_io_outs_0),
    .io_outs_1(ces_6_11_io_outs_1),
    .io_outs_2(ces_6_11_io_outs_2),
    .io_outs_3(ces_6_11_io_outs_3)
  );
  Element ces_6_12 ( // @[MockArray.scala 37:53]
    .clock(ces_6_12_clock),
    .io_ins_0(ces_6_12_io_ins_0),
    .io_ins_1(ces_6_12_io_ins_1),
    .io_ins_2(ces_6_12_io_ins_2),
    .io_ins_3(ces_6_12_io_ins_3),
    .io_outs_0(ces_6_12_io_outs_0),
    .io_outs_1(ces_6_12_io_outs_1),
    .io_outs_2(ces_6_12_io_outs_2),
    .io_outs_3(ces_6_12_io_outs_3)
  );
  Element ces_6_13 ( // @[MockArray.scala 37:53]
    .clock(ces_6_13_clock),
    .io_ins_0(ces_6_13_io_ins_0),
    .io_ins_1(ces_6_13_io_ins_1),
    .io_ins_2(ces_6_13_io_ins_2),
    .io_ins_3(ces_6_13_io_ins_3),
    .io_outs_0(ces_6_13_io_outs_0),
    .io_outs_1(ces_6_13_io_outs_1),
    .io_outs_2(ces_6_13_io_outs_2),
    .io_outs_3(ces_6_13_io_outs_3)
  );
  Element ces_6_14 ( // @[MockArray.scala 37:53]
    .clock(ces_6_14_clock),
    .io_ins_0(ces_6_14_io_ins_0),
    .io_ins_1(ces_6_14_io_ins_1),
    .io_ins_2(ces_6_14_io_ins_2),
    .io_ins_3(ces_6_14_io_ins_3),
    .io_outs_0(ces_6_14_io_outs_0),
    .io_outs_1(ces_6_14_io_outs_1),
    .io_outs_2(ces_6_14_io_outs_2),
    .io_outs_3(ces_6_14_io_outs_3)
  );
  Element ces_6_15 ( // @[MockArray.scala 37:53]
    .clock(ces_6_15_clock),
    .io_ins_0(ces_6_15_io_ins_0),
    .io_ins_1(ces_6_15_io_ins_1),
    .io_ins_2(ces_6_15_io_ins_2),
    .io_ins_3(ces_6_15_io_ins_3),
    .io_outs_0(ces_6_15_io_outs_0),
    .io_outs_1(ces_6_15_io_outs_1),
    .io_outs_2(ces_6_15_io_outs_2),
    .io_outs_3(ces_6_15_io_outs_3)
  );
  Element ces_7_0 ( // @[MockArray.scala 37:53]
    .clock(ces_7_0_clock),
    .io_ins_0(ces_7_0_io_ins_0),
    .io_ins_1(ces_7_0_io_ins_1),
    .io_ins_2(ces_7_0_io_ins_2),
    .io_ins_3(ces_7_0_io_ins_3),
    .io_outs_0(ces_7_0_io_outs_0),
    .io_outs_1(ces_7_0_io_outs_1),
    .io_outs_2(ces_7_0_io_outs_2),
    .io_outs_3(ces_7_0_io_outs_3)
  );
  Element ces_7_1 ( // @[MockArray.scala 37:53]
    .clock(ces_7_1_clock),
    .io_ins_0(ces_7_1_io_ins_0),
    .io_ins_1(ces_7_1_io_ins_1),
    .io_ins_2(ces_7_1_io_ins_2),
    .io_ins_3(ces_7_1_io_ins_3),
    .io_outs_0(ces_7_1_io_outs_0),
    .io_outs_1(ces_7_1_io_outs_1),
    .io_outs_2(ces_7_1_io_outs_2),
    .io_outs_3(ces_7_1_io_outs_3)
  );
  Element ces_7_2 ( // @[MockArray.scala 37:53]
    .clock(ces_7_2_clock),
    .io_ins_0(ces_7_2_io_ins_0),
    .io_ins_1(ces_7_2_io_ins_1),
    .io_ins_2(ces_7_2_io_ins_2),
    .io_ins_3(ces_7_2_io_ins_3),
    .io_outs_0(ces_7_2_io_outs_0),
    .io_outs_1(ces_7_2_io_outs_1),
    .io_outs_2(ces_7_2_io_outs_2),
    .io_outs_3(ces_7_2_io_outs_3)
  );
  Element ces_7_3 ( // @[MockArray.scala 37:53]
    .clock(ces_7_3_clock),
    .io_ins_0(ces_7_3_io_ins_0),
    .io_ins_1(ces_7_3_io_ins_1),
    .io_ins_2(ces_7_3_io_ins_2),
    .io_ins_3(ces_7_3_io_ins_3),
    .io_outs_0(ces_7_3_io_outs_0),
    .io_outs_1(ces_7_3_io_outs_1),
    .io_outs_2(ces_7_3_io_outs_2),
    .io_outs_3(ces_7_3_io_outs_3)
  );
  Element ces_7_4 ( // @[MockArray.scala 37:53]
    .clock(ces_7_4_clock),
    .io_ins_0(ces_7_4_io_ins_0),
    .io_ins_1(ces_7_4_io_ins_1),
    .io_ins_2(ces_7_4_io_ins_2),
    .io_ins_3(ces_7_4_io_ins_3),
    .io_outs_0(ces_7_4_io_outs_0),
    .io_outs_1(ces_7_4_io_outs_1),
    .io_outs_2(ces_7_4_io_outs_2),
    .io_outs_3(ces_7_4_io_outs_3)
  );
  Element ces_7_5 ( // @[MockArray.scala 37:53]
    .clock(ces_7_5_clock),
    .io_ins_0(ces_7_5_io_ins_0),
    .io_ins_1(ces_7_5_io_ins_1),
    .io_ins_2(ces_7_5_io_ins_2),
    .io_ins_3(ces_7_5_io_ins_3),
    .io_outs_0(ces_7_5_io_outs_0),
    .io_outs_1(ces_7_5_io_outs_1),
    .io_outs_2(ces_7_5_io_outs_2),
    .io_outs_3(ces_7_5_io_outs_3)
  );
  Element ces_7_6 ( // @[MockArray.scala 37:53]
    .clock(ces_7_6_clock),
    .io_ins_0(ces_7_6_io_ins_0),
    .io_ins_1(ces_7_6_io_ins_1),
    .io_ins_2(ces_7_6_io_ins_2),
    .io_ins_3(ces_7_6_io_ins_3),
    .io_outs_0(ces_7_6_io_outs_0),
    .io_outs_1(ces_7_6_io_outs_1),
    .io_outs_2(ces_7_6_io_outs_2),
    .io_outs_3(ces_7_6_io_outs_3)
  );
  Element ces_7_7 ( // @[MockArray.scala 37:53]
    .clock(ces_7_7_clock),
    .io_ins_0(ces_7_7_io_ins_0),
    .io_ins_1(ces_7_7_io_ins_1),
    .io_ins_2(ces_7_7_io_ins_2),
    .io_ins_3(ces_7_7_io_ins_3),
    .io_outs_0(ces_7_7_io_outs_0),
    .io_outs_1(ces_7_7_io_outs_1),
    .io_outs_2(ces_7_7_io_outs_2),
    .io_outs_3(ces_7_7_io_outs_3)
  );
  Element ces_7_8 ( // @[MockArray.scala 37:53]
    .clock(ces_7_8_clock),
    .io_ins_0(ces_7_8_io_ins_0),
    .io_ins_1(ces_7_8_io_ins_1),
    .io_ins_2(ces_7_8_io_ins_2),
    .io_ins_3(ces_7_8_io_ins_3),
    .io_outs_0(ces_7_8_io_outs_0),
    .io_outs_1(ces_7_8_io_outs_1),
    .io_outs_2(ces_7_8_io_outs_2),
    .io_outs_3(ces_7_8_io_outs_3)
  );
  Element ces_7_9 ( // @[MockArray.scala 37:53]
    .clock(ces_7_9_clock),
    .io_ins_0(ces_7_9_io_ins_0),
    .io_ins_1(ces_7_9_io_ins_1),
    .io_ins_2(ces_7_9_io_ins_2),
    .io_ins_3(ces_7_9_io_ins_3),
    .io_outs_0(ces_7_9_io_outs_0),
    .io_outs_1(ces_7_9_io_outs_1),
    .io_outs_2(ces_7_9_io_outs_2),
    .io_outs_3(ces_7_9_io_outs_3)
  );
  Element ces_7_10 ( // @[MockArray.scala 37:53]
    .clock(ces_7_10_clock),
    .io_ins_0(ces_7_10_io_ins_0),
    .io_ins_1(ces_7_10_io_ins_1),
    .io_ins_2(ces_7_10_io_ins_2),
    .io_ins_3(ces_7_10_io_ins_3),
    .io_outs_0(ces_7_10_io_outs_0),
    .io_outs_1(ces_7_10_io_outs_1),
    .io_outs_2(ces_7_10_io_outs_2),
    .io_outs_3(ces_7_10_io_outs_3)
  );
  Element ces_7_11 ( // @[MockArray.scala 37:53]
    .clock(ces_7_11_clock),
    .io_ins_0(ces_7_11_io_ins_0),
    .io_ins_1(ces_7_11_io_ins_1),
    .io_ins_2(ces_7_11_io_ins_2),
    .io_ins_3(ces_7_11_io_ins_3),
    .io_outs_0(ces_7_11_io_outs_0),
    .io_outs_1(ces_7_11_io_outs_1),
    .io_outs_2(ces_7_11_io_outs_2),
    .io_outs_3(ces_7_11_io_outs_3)
  );
  Element ces_7_12 ( // @[MockArray.scala 37:53]
    .clock(ces_7_12_clock),
    .io_ins_0(ces_7_12_io_ins_0),
    .io_ins_1(ces_7_12_io_ins_1),
    .io_ins_2(ces_7_12_io_ins_2),
    .io_ins_3(ces_7_12_io_ins_3),
    .io_outs_0(ces_7_12_io_outs_0),
    .io_outs_1(ces_7_12_io_outs_1),
    .io_outs_2(ces_7_12_io_outs_2),
    .io_outs_3(ces_7_12_io_outs_3)
  );
  Element ces_7_13 ( // @[MockArray.scala 37:53]
    .clock(ces_7_13_clock),
    .io_ins_0(ces_7_13_io_ins_0),
    .io_ins_1(ces_7_13_io_ins_1),
    .io_ins_2(ces_7_13_io_ins_2),
    .io_ins_3(ces_7_13_io_ins_3),
    .io_outs_0(ces_7_13_io_outs_0),
    .io_outs_1(ces_7_13_io_outs_1),
    .io_outs_2(ces_7_13_io_outs_2),
    .io_outs_3(ces_7_13_io_outs_3)
  );
  Element ces_7_14 ( // @[MockArray.scala 37:53]
    .clock(ces_7_14_clock),
    .io_ins_0(ces_7_14_io_ins_0),
    .io_ins_1(ces_7_14_io_ins_1),
    .io_ins_2(ces_7_14_io_ins_2),
    .io_ins_3(ces_7_14_io_ins_3),
    .io_outs_0(ces_7_14_io_outs_0),
    .io_outs_1(ces_7_14_io_outs_1),
    .io_outs_2(ces_7_14_io_outs_2),
    .io_outs_3(ces_7_14_io_outs_3)
  );
  Element ces_7_15 ( // @[MockArray.scala 37:53]
    .clock(ces_7_15_clock),
    .io_ins_0(ces_7_15_io_ins_0),
    .io_ins_1(ces_7_15_io_ins_1),
    .io_ins_2(ces_7_15_io_ins_2),
    .io_ins_3(ces_7_15_io_ins_3),
    .io_outs_0(ces_7_15_io_outs_0),
    .io_outs_1(ces_7_15_io_outs_1),
    .io_outs_2(ces_7_15_io_outs_2),
    .io_outs_3(ces_7_15_io_outs_3)
  );
  Element ces_8_0 ( // @[MockArray.scala 37:53]
    .clock(ces_8_0_clock),
    .io_ins_0(ces_8_0_io_ins_0),
    .io_ins_1(ces_8_0_io_ins_1),
    .io_ins_2(ces_8_0_io_ins_2),
    .io_ins_3(ces_8_0_io_ins_3),
    .io_outs_0(ces_8_0_io_outs_0),
    .io_outs_1(ces_8_0_io_outs_1),
    .io_outs_2(ces_8_0_io_outs_2),
    .io_outs_3(ces_8_0_io_outs_3)
  );
  Element ces_8_1 ( // @[MockArray.scala 37:53]
    .clock(ces_8_1_clock),
    .io_ins_0(ces_8_1_io_ins_0),
    .io_ins_1(ces_8_1_io_ins_1),
    .io_ins_2(ces_8_1_io_ins_2),
    .io_ins_3(ces_8_1_io_ins_3),
    .io_outs_0(ces_8_1_io_outs_0),
    .io_outs_1(ces_8_1_io_outs_1),
    .io_outs_2(ces_8_1_io_outs_2),
    .io_outs_3(ces_8_1_io_outs_3)
  );
  Element ces_8_2 ( // @[MockArray.scala 37:53]
    .clock(ces_8_2_clock),
    .io_ins_0(ces_8_2_io_ins_0),
    .io_ins_1(ces_8_2_io_ins_1),
    .io_ins_2(ces_8_2_io_ins_2),
    .io_ins_3(ces_8_2_io_ins_3),
    .io_outs_0(ces_8_2_io_outs_0),
    .io_outs_1(ces_8_2_io_outs_1),
    .io_outs_2(ces_8_2_io_outs_2),
    .io_outs_3(ces_8_2_io_outs_3)
  );
  Element ces_8_3 ( // @[MockArray.scala 37:53]
    .clock(ces_8_3_clock),
    .io_ins_0(ces_8_3_io_ins_0),
    .io_ins_1(ces_8_3_io_ins_1),
    .io_ins_2(ces_8_3_io_ins_2),
    .io_ins_3(ces_8_3_io_ins_3),
    .io_outs_0(ces_8_3_io_outs_0),
    .io_outs_1(ces_8_3_io_outs_1),
    .io_outs_2(ces_8_3_io_outs_2),
    .io_outs_3(ces_8_3_io_outs_3)
  );
  Element ces_8_4 ( // @[MockArray.scala 37:53]
    .clock(ces_8_4_clock),
    .io_ins_0(ces_8_4_io_ins_0),
    .io_ins_1(ces_8_4_io_ins_1),
    .io_ins_2(ces_8_4_io_ins_2),
    .io_ins_3(ces_8_4_io_ins_3),
    .io_outs_0(ces_8_4_io_outs_0),
    .io_outs_1(ces_8_4_io_outs_1),
    .io_outs_2(ces_8_4_io_outs_2),
    .io_outs_3(ces_8_4_io_outs_3)
  );
  Element ces_8_5 ( // @[MockArray.scala 37:53]
    .clock(ces_8_5_clock),
    .io_ins_0(ces_8_5_io_ins_0),
    .io_ins_1(ces_8_5_io_ins_1),
    .io_ins_2(ces_8_5_io_ins_2),
    .io_ins_3(ces_8_5_io_ins_3),
    .io_outs_0(ces_8_5_io_outs_0),
    .io_outs_1(ces_8_5_io_outs_1),
    .io_outs_2(ces_8_5_io_outs_2),
    .io_outs_3(ces_8_5_io_outs_3)
  );
  Element ces_8_6 ( // @[MockArray.scala 37:53]
    .clock(ces_8_6_clock),
    .io_ins_0(ces_8_6_io_ins_0),
    .io_ins_1(ces_8_6_io_ins_1),
    .io_ins_2(ces_8_6_io_ins_2),
    .io_ins_3(ces_8_6_io_ins_3),
    .io_outs_0(ces_8_6_io_outs_0),
    .io_outs_1(ces_8_6_io_outs_1),
    .io_outs_2(ces_8_6_io_outs_2),
    .io_outs_3(ces_8_6_io_outs_3)
  );
  Element ces_8_7 ( // @[MockArray.scala 37:53]
    .clock(ces_8_7_clock),
    .io_ins_0(ces_8_7_io_ins_0),
    .io_ins_1(ces_8_7_io_ins_1),
    .io_ins_2(ces_8_7_io_ins_2),
    .io_ins_3(ces_8_7_io_ins_3),
    .io_outs_0(ces_8_7_io_outs_0),
    .io_outs_1(ces_8_7_io_outs_1),
    .io_outs_2(ces_8_7_io_outs_2),
    .io_outs_3(ces_8_7_io_outs_3)
  );
  Element ces_8_8 ( // @[MockArray.scala 37:53]
    .clock(ces_8_8_clock),
    .io_ins_0(ces_8_8_io_ins_0),
    .io_ins_1(ces_8_8_io_ins_1),
    .io_ins_2(ces_8_8_io_ins_2),
    .io_ins_3(ces_8_8_io_ins_3),
    .io_outs_0(ces_8_8_io_outs_0),
    .io_outs_1(ces_8_8_io_outs_1),
    .io_outs_2(ces_8_8_io_outs_2),
    .io_outs_3(ces_8_8_io_outs_3)
  );
  Element ces_8_9 ( // @[MockArray.scala 37:53]
    .clock(ces_8_9_clock),
    .io_ins_0(ces_8_9_io_ins_0),
    .io_ins_1(ces_8_9_io_ins_1),
    .io_ins_2(ces_8_9_io_ins_2),
    .io_ins_3(ces_8_9_io_ins_3),
    .io_outs_0(ces_8_9_io_outs_0),
    .io_outs_1(ces_8_9_io_outs_1),
    .io_outs_2(ces_8_9_io_outs_2),
    .io_outs_3(ces_8_9_io_outs_3)
  );
  Element ces_8_10 ( // @[MockArray.scala 37:53]
    .clock(ces_8_10_clock),
    .io_ins_0(ces_8_10_io_ins_0),
    .io_ins_1(ces_8_10_io_ins_1),
    .io_ins_2(ces_8_10_io_ins_2),
    .io_ins_3(ces_8_10_io_ins_3),
    .io_outs_0(ces_8_10_io_outs_0),
    .io_outs_1(ces_8_10_io_outs_1),
    .io_outs_2(ces_8_10_io_outs_2),
    .io_outs_3(ces_8_10_io_outs_3)
  );
  Element ces_8_11 ( // @[MockArray.scala 37:53]
    .clock(ces_8_11_clock),
    .io_ins_0(ces_8_11_io_ins_0),
    .io_ins_1(ces_8_11_io_ins_1),
    .io_ins_2(ces_8_11_io_ins_2),
    .io_ins_3(ces_8_11_io_ins_3),
    .io_outs_0(ces_8_11_io_outs_0),
    .io_outs_1(ces_8_11_io_outs_1),
    .io_outs_2(ces_8_11_io_outs_2),
    .io_outs_3(ces_8_11_io_outs_3)
  );
  Element ces_8_12 ( // @[MockArray.scala 37:53]
    .clock(ces_8_12_clock),
    .io_ins_0(ces_8_12_io_ins_0),
    .io_ins_1(ces_8_12_io_ins_1),
    .io_ins_2(ces_8_12_io_ins_2),
    .io_ins_3(ces_8_12_io_ins_3),
    .io_outs_0(ces_8_12_io_outs_0),
    .io_outs_1(ces_8_12_io_outs_1),
    .io_outs_2(ces_8_12_io_outs_2),
    .io_outs_3(ces_8_12_io_outs_3)
  );
  Element ces_8_13 ( // @[MockArray.scala 37:53]
    .clock(ces_8_13_clock),
    .io_ins_0(ces_8_13_io_ins_0),
    .io_ins_1(ces_8_13_io_ins_1),
    .io_ins_2(ces_8_13_io_ins_2),
    .io_ins_3(ces_8_13_io_ins_3),
    .io_outs_0(ces_8_13_io_outs_0),
    .io_outs_1(ces_8_13_io_outs_1),
    .io_outs_2(ces_8_13_io_outs_2),
    .io_outs_3(ces_8_13_io_outs_3)
  );
  Element ces_8_14 ( // @[MockArray.scala 37:53]
    .clock(ces_8_14_clock),
    .io_ins_0(ces_8_14_io_ins_0),
    .io_ins_1(ces_8_14_io_ins_1),
    .io_ins_2(ces_8_14_io_ins_2),
    .io_ins_3(ces_8_14_io_ins_3),
    .io_outs_0(ces_8_14_io_outs_0),
    .io_outs_1(ces_8_14_io_outs_1),
    .io_outs_2(ces_8_14_io_outs_2),
    .io_outs_3(ces_8_14_io_outs_3)
  );
  Element ces_8_15 ( // @[MockArray.scala 37:53]
    .clock(ces_8_15_clock),
    .io_ins_0(ces_8_15_io_ins_0),
    .io_ins_1(ces_8_15_io_ins_1),
    .io_ins_2(ces_8_15_io_ins_2),
    .io_ins_3(ces_8_15_io_ins_3),
    .io_outs_0(ces_8_15_io_outs_0),
    .io_outs_1(ces_8_15_io_outs_1),
    .io_outs_2(ces_8_15_io_outs_2),
    .io_outs_3(ces_8_15_io_outs_3)
  );
  Element ces_9_0 ( // @[MockArray.scala 37:53]
    .clock(ces_9_0_clock),
    .io_ins_0(ces_9_0_io_ins_0),
    .io_ins_1(ces_9_0_io_ins_1),
    .io_ins_2(ces_9_0_io_ins_2),
    .io_ins_3(ces_9_0_io_ins_3),
    .io_outs_0(ces_9_0_io_outs_0),
    .io_outs_1(ces_9_0_io_outs_1),
    .io_outs_2(ces_9_0_io_outs_2),
    .io_outs_3(ces_9_0_io_outs_3)
  );
  Element ces_9_1 ( // @[MockArray.scala 37:53]
    .clock(ces_9_1_clock),
    .io_ins_0(ces_9_1_io_ins_0),
    .io_ins_1(ces_9_1_io_ins_1),
    .io_ins_2(ces_9_1_io_ins_2),
    .io_ins_3(ces_9_1_io_ins_3),
    .io_outs_0(ces_9_1_io_outs_0),
    .io_outs_1(ces_9_1_io_outs_1),
    .io_outs_2(ces_9_1_io_outs_2),
    .io_outs_3(ces_9_1_io_outs_3)
  );
  Element ces_9_2 ( // @[MockArray.scala 37:53]
    .clock(ces_9_2_clock),
    .io_ins_0(ces_9_2_io_ins_0),
    .io_ins_1(ces_9_2_io_ins_1),
    .io_ins_2(ces_9_2_io_ins_2),
    .io_ins_3(ces_9_2_io_ins_3),
    .io_outs_0(ces_9_2_io_outs_0),
    .io_outs_1(ces_9_2_io_outs_1),
    .io_outs_2(ces_9_2_io_outs_2),
    .io_outs_3(ces_9_2_io_outs_3)
  );
  Element ces_9_3 ( // @[MockArray.scala 37:53]
    .clock(ces_9_3_clock),
    .io_ins_0(ces_9_3_io_ins_0),
    .io_ins_1(ces_9_3_io_ins_1),
    .io_ins_2(ces_9_3_io_ins_2),
    .io_ins_3(ces_9_3_io_ins_3),
    .io_outs_0(ces_9_3_io_outs_0),
    .io_outs_1(ces_9_3_io_outs_1),
    .io_outs_2(ces_9_3_io_outs_2),
    .io_outs_3(ces_9_3_io_outs_3)
  );
  Element ces_9_4 ( // @[MockArray.scala 37:53]
    .clock(ces_9_4_clock),
    .io_ins_0(ces_9_4_io_ins_0),
    .io_ins_1(ces_9_4_io_ins_1),
    .io_ins_2(ces_9_4_io_ins_2),
    .io_ins_3(ces_9_4_io_ins_3),
    .io_outs_0(ces_9_4_io_outs_0),
    .io_outs_1(ces_9_4_io_outs_1),
    .io_outs_2(ces_9_4_io_outs_2),
    .io_outs_3(ces_9_4_io_outs_3)
  );
  Element ces_9_5 ( // @[MockArray.scala 37:53]
    .clock(ces_9_5_clock),
    .io_ins_0(ces_9_5_io_ins_0),
    .io_ins_1(ces_9_5_io_ins_1),
    .io_ins_2(ces_9_5_io_ins_2),
    .io_ins_3(ces_9_5_io_ins_3),
    .io_outs_0(ces_9_5_io_outs_0),
    .io_outs_1(ces_9_5_io_outs_1),
    .io_outs_2(ces_9_5_io_outs_2),
    .io_outs_3(ces_9_5_io_outs_3)
  );
  Element ces_9_6 ( // @[MockArray.scala 37:53]
    .clock(ces_9_6_clock),
    .io_ins_0(ces_9_6_io_ins_0),
    .io_ins_1(ces_9_6_io_ins_1),
    .io_ins_2(ces_9_6_io_ins_2),
    .io_ins_3(ces_9_6_io_ins_3),
    .io_outs_0(ces_9_6_io_outs_0),
    .io_outs_1(ces_9_6_io_outs_1),
    .io_outs_2(ces_9_6_io_outs_2),
    .io_outs_3(ces_9_6_io_outs_3)
  );
  Element ces_9_7 ( // @[MockArray.scala 37:53]
    .clock(ces_9_7_clock),
    .io_ins_0(ces_9_7_io_ins_0),
    .io_ins_1(ces_9_7_io_ins_1),
    .io_ins_2(ces_9_7_io_ins_2),
    .io_ins_3(ces_9_7_io_ins_3),
    .io_outs_0(ces_9_7_io_outs_0),
    .io_outs_1(ces_9_7_io_outs_1),
    .io_outs_2(ces_9_7_io_outs_2),
    .io_outs_3(ces_9_7_io_outs_3)
  );
  Element ces_9_8 ( // @[MockArray.scala 37:53]
    .clock(ces_9_8_clock),
    .io_ins_0(ces_9_8_io_ins_0),
    .io_ins_1(ces_9_8_io_ins_1),
    .io_ins_2(ces_9_8_io_ins_2),
    .io_ins_3(ces_9_8_io_ins_3),
    .io_outs_0(ces_9_8_io_outs_0),
    .io_outs_1(ces_9_8_io_outs_1),
    .io_outs_2(ces_9_8_io_outs_2),
    .io_outs_3(ces_9_8_io_outs_3)
  );
  Element ces_9_9 ( // @[MockArray.scala 37:53]
    .clock(ces_9_9_clock),
    .io_ins_0(ces_9_9_io_ins_0),
    .io_ins_1(ces_9_9_io_ins_1),
    .io_ins_2(ces_9_9_io_ins_2),
    .io_ins_3(ces_9_9_io_ins_3),
    .io_outs_0(ces_9_9_io_outs_0),
    .io_outs_1(ces_9_9_io_outs_1),
    .io_outs_2(ces_9_9_io_outs_2),
    .io_outs_3(ces_9_9_io_outs_3)
  );
  Element ces_9_10 ( // @[MockArray.scala 37:53]
    .clock(ces_9_10_clock),
    .io_ins_0(ces_9_10_io_ins_0),
    .io_ins_1(ces_9_10_io_ins_1),
    .io_ins_2(ces_9_10_io_ins_2),
    .io_ins_3(ces_9_10_io_ins_3),
    .io_outs_0(ces_9_10_io_outs_0),
    .io_outs_1(ces_9_10_io_outs_1),
    .io_outs_2(ces_9_10_io_outs_2),
    .io_outs_3(ces_9_10_io_outs_3)
  );
  Element ces_9_11 ( // @[MockArray.scala 37:53]
    .clock(ces_9_11_clock),
    .io_ins_0(ces_9_11_io_ins_0),
    .io_ins_1(ces_9_11_io_ins_1),
    .io_ins_2(ces_9_11_io_ins_2),
    .io_ins_3(ces_9_11_io_ins_3),
    .io_outs_0(ces_9_11_io_outs_0),
    .io_outs_1(ces_9_11_io_outs_1),
    .io_outs_2(ces_9_11_io_outs_2),
    .io_outs_3(ces_9_11_io_outs_3)
  );
  Element ces_9_12 ( // @[MockArray.scala 37:53]
    .clock(ces_9_12_clock),
    .io_ins_0(ces_9_12_io_ins_0),
    .io_ins_1(ces_9_12_io_ins_1),
    .io_ins_2(ces_9_12_io_ins_2),
    .io_ins_3(ces_9_12_io_ins_3),
    .io_outs_0(ces_9_12_io_outs_0),
    .io_outs_1(ces_9_12_io_outs_1),
    .io_outs_2(ces_9_12_io_outs_2),
    .io_outs_3(ces_9_12_io_outs_3)
  );
  Element ces_9_13 ( // @[MockArray.scala 37:53]
    .clock(ces_9_13_clock),
    .io_ins_0(ces_9_13_io_ins_0),
    .io_ins_1(ces_9_13_io_ins_1),
    .io_ins_2(ces_9_13_io_ins_2),
    .io_ins_3(ces_9_13_io_ins_3),
    .io_outs_0(ces_9_13_io_outs_0),
    .io_outs_1(ces_9_13_io_outs_1),
    .io_outs_2(ces_9_13_io_outs_2),
    .io_outs_3(ces_9_13_io_outs_3)
  );
  Element ces_9_14 ( // @[MockArray.scala 37:53]
    .clock(ces_9_14_clock),
    .io_ins_0(ces_9_14_io_ins_0),
    .io_ins_1(ces_9_14_io_ins_1),
    .io_ins_2(ces_9_14_io_ins_2),
    .io_ins_3(ces_9_14_io_ins_3),
    .io_outs_0(ces_9_14_io_outs_0),
    .io_outs_1(ces_9_14_io_outs_1),
    .io_outs_2(ces_9_14_io_outs_2),
    .io_outs_3(ces_9_14_io_outs_3)
  );
  Element ces_9_15 ( // @[MockArray.scala 37:53]
    .clock(ces_9_15_clock),
    .io_ins_0(ces_9_15_io_ins_0),
    .io_ins_1(ces_9_15_io_ins_1),
    .io_ins_2(ces_9_15_io_ins_2),
    .io_ins_3(ces_9_15_io_ins_3),
    .io_outs_0(ces_9_15_io_outs_0),
    .io_outs_1(ces_9_15_io_outs_1),
    .io_outs_2(ces_9_15_io_outs_2),
    .io_outs_3(ces_9_15_io_outs_3)
  );
  Element ces_10_0 ( // @[MockArray.scala 37:53]
    .clock(ces_10_0_clock),
    .io_ins_0(ces_10_0_io_ins_0),
    .io_ins_1(ces_10_0_io_ins_1),
    .io_ins_2(ces_10_0_io_ins_2),
    .io_ins_3(ces_10_0_io_ins_3),
    .io_outs_0(ces_10_0_io_outs_0),
    .io_outs_1(ces_10_0_io_outs_1),
    .io_outs_2(ces_10_0_io_outs_2),
    .io_outs_3(ces_10_0_io_outs_3)
  );
  Element ces_10_1 ( // @[MockArray.scala 37:53]
    .clock(ces_10_1_clock),
    .io_ins_0(ces_10_1_io_ins_0),
    .io_ins_1(ces_10_1_io_ins_1),
    .io_ins_2(ces_10_1_io_ins_2),
    .io_ins_3(ces_10_1_io_ins_3),
    .io_outs_0(ces_10_1_io_outs_0),
    .io_outs_1(ces_10_1_io_outs_1),
    .io_outs_2(ces_10_1_io_outs_2),
    .io_outs_3(ces_10_1_io_outs_3)
  );
  Element ces_10_2 ( // @[MockArray.scala 37:53]
    .clock(ces_10_2_clock),
    .io_ins_0(ces_10_2_io_ins_0),
    .io_ins_1(ces_10_2_io_ins_1),
    .io_ins_2(ces_10_2_io_ins_2),
    .io_ins_3(ces_10_2_io_ins_3),
    .io_outs_0(ces_10_2_io_outs_0),
    .io_outs_1(ces_10_2_io_outs_1),
    .io_outs_2(ces_10_2_io_outs_2),
    .io_outs_3(ces_10_2_io_outs_3)
  );
  Element ces_10_3 ( // @[MockArray.scala 37:53]
    .clock(ces_10_3_clock),
    .io_ins_0(ces_10_3_io_ins_0),
    .io_ins_1(ces_10_3_io_ins_1),
    .io_ins_2(ces_10_3_io_ins_2),
    .io_ins_3(ces_10_3_io_ins_3),
    .io_outs_0(ces_10_3_io_outs_0),
    .io_outs_1(ces_10_3_io_outs_1),
    .io_outs_2(ces_10_3_io_outs_2),
    .io_outs_3(ces_10_3_io_outs_3)
  );
  Element ces_10_4 ( // @[MockArray.scala 37:53]
    .clock(ces_10_4_clock),
    .io_ins_0(ces_10_4_io_ins_0),
    .io_ins_1(ces_10_4_io_ins_1),
    .io_ins_2(ces_10_4_io_ins_2),
    .io_ins_3(ces_10_4_io_ins_3),
    .io_outs_0(ces_10_4_io_outs_0),
    .io_outs_1(ces_10_4_io_outs_1),
    .io_outs_2(ces_10_4_io_outs_2),
    .io_outs_3(ces_10_4_io_outs_3)
  );
  Element ces_10_5 ( // @[MockArray.scala 37:53]
    .clock(ces_10_5_clock),
    .io_ins_0(ces_10_5_io_ins_0),
    .io_ins_1(ces_10_5_io_ins_1),
    .io_ins_2(ces_10_5_io_ins_2),
    .io_ins_3(ces_10_5_io_ins_3),
    .io_outs_0(ces_10_5_io_outs_0),
    .io_outs_1(ces_10_5_io_outs_1),
    .io_outs_2(ces_10_5_io_outs_2),
    .io_outs_3(ces_10_5_io_outs_3)
  );
  Element ces_10_6 ( // @[MockArray.scala 37:53]
    .clock(ces_10_6_clock),
    .io_ins_0(ces_10_6_io_ins_0),
    .io_ins_1(ces_10_6_io_ins_1),
    .io_ins_2(ces_10_6_io_ins_2),
    .io_ins_3(ces_10_6_io_ins_3),
    .io_outs_0(ces_10_6_io_outs_0),
    .io_outs_1(ces_10_6_io_outs_1),
    .io_outs_2(ces_10_6_io_outs_2),
    .io_outs_3(ces_10_6_io_outs_3)
  );
  Element ces_10_7 ( // @[MockArray.scala 37:53]
    .clock(ces_10_7_clock),
    .io_ins_0(ces_10_7_io_ins_0),
    .io_ins_1(ces_10_7_io_ins_1),
    .io_ins_2(ces_10_7_io_ins_2),
    .io_ins_3(ces_10_7_io_ins_3),
    .io_outs_0(ces_10_7_io_outs_0),
    .io_outs_1(ces_10_7_io_outs_1),
    .io_outs_2(ces_10_7_io_outs_2),
    .io_outs_3(ces_10_7_io_outs_3)
  );
  Element ces_10_8 ( // @[MockArray.scala 37:53]
    .clock(ces_10_8_clock),
    .io_ins_0(ces_10_8_io_ins_0),
    .io_ins_1(ces_10_8_io_ins_1),
    .io_ins_2(ces_10_8_io_ins_2),
    .io_ins_3(ces_10_8_io_ins_3),
    .io_outs_0(ces_10_8_io_outs_0),
    .io_outs_1(ces_10_8_io_outs_1),
    .io_outs_2(ces_10_8_io_outs_2),
    .io_outs_3(ces_10_8_io_outs_3)
  );
  Element ces_10_9 ( // @[MockArray.scala 37:53]
    .clock(ces_10_9_clock),
    .io_ins_0(ces_10_9_io_ins_0),
    .io_ins_1(ces_10_9_io_ins_1),
    .io_ins_2(ces_10_9_io_ins_2),
    .io_ins_3(ces_10_9_io_ins_3),
    .io_outs_0(ces_10_9_io_outs_0),
    .io_outs_1(ces_10_9_io_outs_1),
    .io_outs_2(ces_10_9_io_outs_2),
    .io_outs_3(ces_10_9_io_outs_3)
  );
  Element ces_10_10 ( // @[MockArray.scala 37:53]
    .clock(ces_10_10_clock),
    .io_ins_0(ces_10_10_io_ins_0),
    .io_ins_1(ces_10_10_io_ins_1),
    .io_ins_2(ces_10_10_io_ins_2),
    .io_ins_3(ces_10_10_io_ins_3),
    .io_outs_0(ces_10_10_io_outs_0),
    .io_outs_1(ces_10_10_io_outs_1),
    .io_outs_2(ces_10_10_io_outs_2),
    .io_outs_3(ces_10_10_io_outs_3)
  );
  Element ces_10_11 ( // @[MockArray.scala 37:53]
    .clock(ces_10_11_clock),
    .io_ins_0(ces_10_11_io_ins_0),
    .io_ins_1(ces_10_11_io_ins_1),
    .io_ins_2(ces_10_11_io_ins_2),
    .io_ins_3(ces_10_11_io_ins_3),
    .io_outs_0(ces_10_11_io_outs_0),
    .io_outs_1(ces_10_11_io_outs_1),
    .io_outs_2(ces_10_11_io_outs_2),
    .io_outs_3(ces_10_11_io_outs_3)
  );
  Element ces_10_12 ( // @[MockArray.scala 37:53]
    .clock(ces_10_12_clock),
    .io_ins_0(ces_10_12_io_ins_0),
    .io_ins_1(ces_10_12_io_ins_1),
    .io_ins_2(ces_10_12_io_ins_2),
    .io_ins_3(ces_10_12_io_ins_3),
    .io_outs_0(ces_10_12_io_outs_0),
    .io_outs_1(ces_10_12_io_outs_1),
    .io_outs_2(ces_10_12_io_outs_2),
    .io_outs_3(ces_10_12_io_outs_3)
  );
  Element ces_10_13 ( // @[MockArray.scala 37:53]
    .clock(ces_10_13_clock),
    .io_ins_0(ces_10_13_io_ins_0),
    .io_ins_1(ces_10_13_io_ins_1),
    .io_ins_2(ces_10_13_io_ins_2),
    .io_ins_3(ces_10_13_io_ins_3),
    .io_outs_0(ces_10_13_io_outs_0),
    .io_outs_1(ces_10_13_io_outs_1),
    .io_outs_2(ces_10_13_io_outs_2),
    .io_outs_3(ces_10_13_io_outs_3)
  );
  Element ces_10_14 ( // @[MockArray.scala 37:53]
    .clock(ces_10_14_clock),
    .io_ins_0(ces_10_14_io_ins_0),
    .io_ins_1(ces_10_14_io_ins_1),
    .io_ins_2(ces_10_14_io_ins_2),
    .io_ins_3(ces_10_14_io_ins_3),
    .io_outs_0(ces_10_14_io_outs_0),
    .io_outs_1(ces_10_14_io_outs_1),
    .io_outs_2(ces_10_14_io_outs_2),
    .io_outs_3(ces_10_14_io_outs_3)
  );
  Element ces_10_15 ( // @[MockArray.scala 37:53]
    .clock(ces_10_15_clock),
    .io_ins_0(ces_10_15_io_ins_0),
    .io_ins_1(ces_10_15_io_ins_1),
    .io_ins_2(ces_10_15_io_ins_2),
    .io_ins_3(ces_10_15_io_ins_3),
    .io_outs_0(ces_10_15_io_outs_0),
    .io_outs_1(ces_10_15_io_outs_1),
    .io_outs_2(ces_10_15_io_outs_2),
    .io_outs_3(ces_10_15_io_outs_3)
  );
  Element ces_11_0 ( // @[MockArray.scala 37:53]
    .clock(ces_11_0_clock),
    .io_ins_0(ces_11_0_io_ins_0),
    .io_ins_1(ces_11_0_io_ins_1),
    .io_ins_2(ces_11_0_io_ins_2),
    .io_ins_3(ces_11_0_io_ins_3),
    .io_outs_0(ces_11_0_io_outs_0),
    .io_outs_1(ces_11_0_io_outs_1),
    .io_outs_2(ces_11_0_io_outs_2),
    .io_outs_3(ces_11_0_io_outs_3)
  );
  Element ces_11_1 ( // @[MockArray.scala 37:53]
    .clock(ces_11_1_clock),
    .io_ins_0(ces_11_1_io_ins_0),
    .io_ins_1(ces_11_1_io_ins_1),
    .io_ins_2(ces_11_1_io_ins_2),
    .io_ins_3(ces_11_1_io_ins_3),
    .io_outs_0(ces_11_1_io_outs_0),
    .io_outs_1(ces_11_1_io_outs_1),
    .io_outs_2(ces_11_1_io_outs_2),
    .io_outs_3(ces_11_1_io_outs_3)
  );
  Element ces_11_2 ( // @[MockArray.scala 37:53]
    .clock(ces_11_2_clock),
    .io_ins_0(ces_11_2_io_ins_0),
    .io_ins_1(ces_11_2_io_ins_1),
    .io_ins_2(ces_11_2_io_ins_2),
    .io_ins_3(ces_11_2_io_ins_3),
    .io_outs_0(ces_11_2_io_outs_0),
    .io_outs_1(ces_11_2_io_outs_1),
    .io_outs_2(ces_11_2_io_outs_2),
    .io_outs_3(ces_11_2_io_outs_3)
  );
  Element ces_11_3 ( // @[MockArray.scala 37:53]
    .clock(ces_11_3_clock),
    .io_ins_0(ces_11_3_io_ins_0),
    .io_ins_1(ces_11_3_io_ins_1),
    .io_ins_2(ces_11_3_io_ins_2),
    .io_ins_3(ces_11_3_io_ins_3),
    .io_outs_0(ces_11_3_io_outs_0),
    .io_outs_1(ces_11_3_io_outs_1),
    .io_outs_2(ces_11_3_io_outs_2),
    .io_outs_3(ces_11_3_io_outs_3)
  );
  Element ces_11_4 ( // @[MockArray.scala 37:53]
    .clock(ces_11_4_clock),
    .io_ins_0(ces_11_4_io_ins_0),
    .io_ins_1(ces_11_4_io_ins_1),
    .io_ins_2(ces_11_4_io_ins_2),
    .io_ins_3(ces_11_4_io_ins_3),
    .io_outs_0(ces_11_4_io_outs_0),
    .io_outs_1(ces_11_4_io_outs_1),
    .io_outs_2(ces_11_4_io_outs_2),
    .io_outs_3(ces_11_4_io_outs_3)
  );
  Element ces_11_5 ( // @[MockArray.scala 37:53]
    .clock(ces_11_5_clock),
    .io_ins_0(ces_11_5_io_ins_0),
    .io_ins_1(ces_11_5_io_ins_1),
    .io_ins_2(ces_11_5_io_ins_2),
    .io_ins_3(ces_11_5_io_ins_3),
    .io_outs_0(ces_11_5_io_outs_0),
    .io_outs_1(ces_11_5_io_outs_1),
    .io_outs_2(ces_11_5_io_outs_2),
    .io_outs_3(ces_11_5_io_outs_3)
  );
  Element ces_11_6 ( // @[MockArray.scala 37:53]
    .clock(ces_11_6_clock),
    .io_ins_0(ces_11_6_io_ins_0),
    .io_ins_1(ces_11_6_io_ins_1),
    .io_ins_2(ces_11_6_io_ins_2),
    .io_ins_3(ces_11_6_io_ins_3),
    .io_outs_0(ces_11_6_io_outs_0),
    .io_outs_1(ces_11_6_io_outs_1),
    .io_outs_2(ces_11_6_io_outs_2),
    .io_outs_3(ces_11_6_io_outs_3)
  );
  Element ces_11_7 ( // @[MockArray.scala 37:53]
    .clock(ces_11_7_clock),
    .io_ins_0(ces_11_7_io_ins_0),
    .io_ins_1(ces_11_7_io_ins_1),
    .io_ins_2(ces_11_7_io_ins_2),
    .io_ins_3(ces_11_7_io_ins_3),
    .io_outs_0(ces_11_7_io_outs_0),
    .io_outs_1(ces_11_7_io_outs_1),
    .io_outs_2(ces_11_7_io_outs_2),
    .io_outs_3(ces_11_7_io_outs_3)
  );
  Element ces_11_8 ( // @[MockArray.scala 37:53]
    .clock(ces_11_8_clock),
    .io_ins_0(ces_11_8_io_ins_0),
    .io_ins_1(ces_11_8_io_ins_1),
    .io_ins_2(ces_11_8_io_ins_2),
    .io_ins_3(ces_11_8_io_ins_3),
    .io_outs_0(ces_11_8_io_outs_0),
    .io_outs_1(ces_11_8_io_outs_1),
    .io_outs_2(ces_11_8_io_outs_2),
    .io_outs_3(ces_11_8_io_outs_3)
  );
  Element ces_11_9 ( // @[MockArray.scala 37:53]
    .clock(ces_11_9_clock),
    .io_ins_0(ces_11_9_io_ins_0),
    .io_ins_1(ces_11_9_io_ins_1),
    .io_ins_2(ces_11_9_io_ins_2),
    .io_ins_3(ces_11_9_io_ins_3),
    .io_outs_0(ces_11_9_io_outs_0),
    .io_outs_1(ces_11_9_io_outs_1),
    .io_outs_2(ces_11_9_io_outs_2),
    .io_outs_3(ces_11_9_io_outs_3)
  );
  Element ces_11_10 ( // @[MockArray.scala 37:53]
    .clock(ces_11_10_clock),
    .io_ins_0(ces_11_10_io_ins_0),
    .io_ins_1(ces_11_10_io_ins_1),
    .io_ins_2(ces_11_10_io_ins_2),
    .io_ins_3(ces_11_10_io_ins_3),
    .io_outs_0(ces_11_10_io_outs_0),
    .io_outs_1(ces_11_10_io_outs_1),
    .io_outs_2(ces_11_10_io_outs_2),
    .io_outs_3(ces_11_10_io_outs_3)
  );
  Element ces_11_11 ( // @[MockArray.scala 37:53]
    .clock(ces_11_11_clock),
    .io_ins_0(ces_11_11_io_ins_0),
    .io_ins_1(ces_11_11_io_ins_1),
    .io_ins_2(ces_11_11_io_ins_2),
    .io_ins_3(ces_11_11_io_ins_3),
    .io_outs_0(ces_11_11_io_outs_0),
    .io_outs_1(ces_11_11_io_outs_1),
    .io_outs_2(ces_11_11_io_outs_2),
    .io_outs_3(ces_11_11_io_outs_3)
  );
  Element ces_11_12 ( // @[MockArray.scala 37:53]
    .clock(ces_11_12_clock),
    .io_ins_0(ces_11_12_io_ins_0),
    .io_ins_1(ces_11_12_io_ins_1),
    .io_ins_2(ces_11_12_io_ins_2),
    .io_ins_3(ces_11_12_io_ins_3),
    .io_outs_0(ces_11_12_io_outs_0),
    .io_outs_1(ces_11_12_io_outs_1),
    .io_outs_2(ces_11_12_io_outs_2),
    .io_outs_3(ces_11_12_io_outs_3)
  );
  Element ces_11_13 ( // @[MockArray.scala 37:53]
    .clock(ces_11_13_clock),
    .io_ins_0(ces_11_13_io_ins_0),
    .io_ins_1(ces_11_13_io_ins_1),
    .io_ins_2(ces_11_13_io_ins_2),
    .io_ins_3(ces_11_13_io_ins_3),
    .io_outs_0(ces_11_13_io_outs_0),
    .io_outs_1(ces_11_13_io_outs_1),
    .io_outs_2(ces_11_13_io_outs_2),
    .io_outs_3(ces_11_13_io_outs_3)
  );
  Element ces_11_14 ( // @[MockArray.scala 37:53]
    .clock(ces_11_14_clock),
    .io_ins_0(ces_11_14_io_ins_0),
    .io_ins_1(ces_11_14_io_ins_1),
    .io_ins_2(ces_11_14_io_ins_2),
    .io_ins_3(ces_11_14_io_ins_3),
    .io_outs_0(ces_11_14_io_outs_0),
    .io_outs_1(ces_11_14_io_outs_1),
    .io_outs_2(ces_11_14_io_outs_2),
    .io_outs_3(ces_11_14_io_outs_3)
  );
  Element ces_11_15 ( // @[MockArray.scala 37:53]
    .clock(ces_11_15_clock),
    .io_ins_0(ces_11_15_io_ins_0),
    .io_ins_1(ces_11_15_io_ins_1),
    .io_ins_2(ces_11_15_io_ins_2),
    .io_ins_3(ces_11_15_io_ins_3),
    .io_outs_0(ces_11_15_io_outs_0),
    .io_outs_1(ces_11_15_io_outs_1),
    .io_outs_2(ces_11_15_io_outs_2),
    .io_outs_3(ces_11_15_io_outs_3)
  );
  Element ces_12_0 ( // @[MockArray.scala 37:53]
    .clock(ces_12_0_clock),
    .io_ins_0(ces_12_0_io_ins_0),
    .io_ins_1(ces_12_0_io_ins_1),
    .io_ins_2(ces_12_0_io_ins_2),
    .io_ins_3(ces_12_0_io_ins_3),
    .io_outs_0(ces_12_0_io_outs_0),
    .io_outs_1(ces_12_0_io_outs_1),
    .io_outs_2(ces_12_0_io_outs_2),
    .io_outs_3(ces_12_0_io_outs_3)
  );
  Element ces_12_1 ( // @[MockArray.scala 37:53]
    .clock(ces_12_1_clock),
    .io_ins_0(ces_12_1_io_ins_0),
    .io_ins_1(ces_12_1_io_ins_1),
    .io_ins_2(ces_12_1_io_ins_2),
    .io_ins_3(ces_12_1_io_ins_3),
    .io_outs_0(ces_12_1_io_outs_0),
    .io_outs_1(ces_12_1_io_outs_1),
    .io_outs_2(ces_12_1_io_outs_2),
    .io_outs_3(ces_12_1_io_outs_3)
  );
  Element ces_12_2 ( // @[MockArray.scala 37:53]
    .clock(ces_12_2_clock),
    .io_ins_0(ces_12_2_io_ins_0),
    .io_ins_1(ces_12_2_io_ins_1),
    .io_ins_2(ces_12_2_io_ins_2),
    .io_ins_3(ces_12_2_io_ins_3),
    .io_outs_0(ces_12_2_io_outs_0),
    .io_outs_1(ces_12_2_io_outs_1),
    .io_outs_2(ces_12_2_io_outs_2),
    .io_outs_3(ces_12_2_io_outs_3)
  );
  Element ces_12_3 ( // @[MockArray.scala 37:53]
    .clock(ces_12_3_clock),
    .io_ins_0(ces_12_3_io_ins_0),
    .io_ins_1(ces_12_3_io_ins_1),
    .io_ins_2(ces_12_3_io_ins_2),
    .io_ins_3(ces_12_3_io_ins_3),
    .io_outs_0(ces_12_3_io_outs_0),
    .io_outs_1(ces_12_3_io_outs_1),
    .io_outs_2(ces_12_3_io_outs_2),
    .io_outs_3(ces_12_3_io_outs_3)
  );
  Element ces_12_4 ( // @[MockArray.scala 37:53]
    .clock(ces_12_4_clock),
    .io_ins_0(ces_12_4_io_ins_0),
    .io_ins_1(ces_12_4_io_ins_1),
    .io_ins_2(ces_12_4_io_ins_2),
    .io_ins_3(ces_12_4_io_ins_3),
    .io_outs_0(ces_12_4_io_outs_0),
    .io_outs_1(ces_12_4_io_outs_1),
    .io_outs_2(ces_12_4_io_outs_2),
    .io_outs_3(ces_12_4_io_outs_3)
  );
  Element ces_12_5 ( // @[MockArray.scala 37:53]
    .clock(ces_12_5_clock),
    .io_ins_0(ces_12_5_io_ins_0),
    .io_ins_1(ces_12_5_io_ins_1),
    .io_ins_2(ces_12_5_io_ins_2),
    .io_ins_3(ces_12_5_io_ins_3),
    .io_outs_0(ces_12_5_io_outs_0),
    .io_outs_1(ces_12_5_io_outs_1),
    .io_outs_2(ces_12_5_io_outs_2),
    .io_outs_3(ces_12_5_io_outs_3)
  );
  Element ces_12_6 ( // @[MockArray.scala 37:53]
    .clock(ces_12_6_clock),
    .io_ins_0(ces_12_6_io_ins_0),
    .io_ins_1(ces_12_6_io_ins_1),
    .io_ins_2(ces_12_6_io_ins_2),
    .io_ins_3(ces_12_6_io_ins_3),
    .io_outs_0(ces_12_6_io_outs_0),
    .io_outs_1(ces_12_6_io_outs_1),
    .io_outs_2(ces_12_6_io_outs_2),
    .io_outs_3(ces_12_6_io_outs_3)
  );
  Element ces_12_7 ( // @[MockArray.scala 37:53]
    .clock(ces_12_7_clock),
    .io_ins_0(ces_12_7_io_ins_0),
    .io_ins_1(ces_12_7_io_ins_1),
    .io_ins_2(ces_12_7_io_ins_2),
    .io_ins_3(ces_12_7_io_ins_3),
    .io_outs_0(ces_12_7_io_outs_0),
    .io_outs_1(ces_12_7_io_outs_1),
    .io_outs_2(ces_12_7_io_outs_2),
    .io_outs_3(ces_12_7_io_outs_3)
  );
  Element ces_12_8 ( // @[MockArray.scala 37:53]
    .clock(ces_12_8_clock),
    .io_ins_0(ces_12_8_io_ins_0),
    .io_ins_1(ces_12_8_io_ins_1),
    .io_ins_2(ces_12_8_io_ins_2),
    .io_ins_3(ces_12_8_io_ins_3),
    .io_outs_0(ces_12_8_io_outs_0),
    .io_outs_1(ces_12_8_io_outs_1),
    .io_outs_2(ces_12_8_io_outs_2),
    .io_outs_3(ces_12_8_io_outs_3)
  );
  Element ces_12_9 ( // @[MockArray.scala 37:53]
    .clock(ces_12_9_clock),
    .io_ins_0(ces_12_9_io_ins_0),
    .io_ins_1(ces_12_9_io_ins_1),
    .io_ins_2(ces_12_9_io_ins_2),
    .io_ins_3(ces_12_9_io_ins_3),
    .io_outs_0(ces_12_9_io_outs_0),
    .io_outs_1(ces_12_9_io_outs_1),
    .io_outs_2(ces_12_9_io_outs_2),
    .io_outs_3(ces_12_9_io_outs_3)
  );
  Element ces_12_10 ( // @[MockArray.scala 37:53]
    .clock(ces_12_10_clock),
    .io_ins_0(ces_12_10_io_ins_0),
    .io_ins_1(ces_12_10_io_ins_1),
    .io_ins_2(ces_12_10_io_ins_2),
    .io_ins_3(ces_12_10_io_ins_3),
    .io_outs_0(ces_12_10_io_outs_0),
    .io_outs_1(ces_12_10_io_outs_1),
    .io_outs_2(ces_12_10_io_outs_2),
    .io_outs_3(ces_12_10_io_outs_3)
  );
  Element ces_12_11 ( // @[MockArray.scala 37:53]
    .clock(ces_12_11_clock),
    .io_ins_0(ces_12_11_io_ins_0),
    .io_ins_1(ces_12_11_io_ins_1),
    .io_ins_2(ces_12_11_io_ins_2),
    .io_ins_3(ces_12_11_io_ins_3),
    .io_outs_0(ces_12_11_io_outs_0),
    .io_outs_1(ces_12_11_io_outs_1),
    .io_outs_2(ces_12_11_io_outs_2),
    .io_outs_3(ces_12_11_io_outs_3)
  );
  Element ces_12_12 ( // @[MockArray.scala 37:53]
    .clock(ces_12_12_clock),
    .io_ins_0(ces_12_12_io_ins_0),
    .io_ins_1(ces_12_12_io_ins_1),
    .io_ins_2(ces_12_12_io_ins_2),
    .io_ins_3(ces_12_12_io_ins_3),
    .io_outs_0(ces_12_12_io_outs_0),
    .io_outs_1(ces_12_12_io_outs_1),
    .io_outs_2(ces_12_12_io_outs_2),
    .io_outs_3(ces_12_12_io_outs_3)
  );
  Element ces_12_13 ( // @[MockArray.scala 37:53]
    .clock(ces_12_13_clock),
    .io_ins_0(ces_12_13_io_ins_0),
    .io_ins_1(ces_12_13_io_ins_1),
    .io_ins_2(ces_12_13_io_ins_2),
    .io_ins_3(ces_12_13_io_ins_3),
    .io_outs_0(ces_12_13_io_outs_0),
    .io_outs_1(ces_12_13_io_outs_1),
    .io_outs_2(ces_12_13_io_outs_2),
    .io_outs_3(ces_12_13_io_outs_3)
  );
  Element ces_12_14 ( // @[MockArray.scala 37:53]
    .clock(ces_12_14_clock),
    .io_ins_0(ces_12_14_io_ins_0),
    .io_ins_1(ces_12_14_io_ins_1),
    .io_ins_2(ces_12_14_io_ins_2),
    .io_ins_3(ces_12_14_io_ins_3),
    .io_outs_0(ces_12_14_io_outs_0),
    .io_outs_1(ces_12_14_io_outs_1),
    .io_outs_2(ces_12_14_io_outs_2),
    .io_outs_3(ces_12_14_io_outs_3)
  );
  Element ces_12_15 ( // @[MockArray.scala 37:53]
    .clock(ces_12_15_clock),
    .io_ins_0(ces_12_15_io_ins_0),
    .io_ins_1(ces_12_15_io_ins_1),
    .io_ins_2(ces_12_15_io_ins_2),
    .io_ins_3(ces_12_15_io_ins_3),
    .io_outs_0(ces_12_15_io_outs_0),
    .io_outs_1(ces_12_15_io_outs_1),
    .io_outs_2(ces_12_15_io_outs_2),
    .io_outs_3(ces_12_15_io_outs_3)
  );
  Element ces_13_0 ( // @[MockArray.scala 37:53]
    .clock(ces_13_0_clock),
    .io_ins_0(ces_13_0_io_ins_0),
    .io_ins_1(ces_13_0_io_ins_1),
    .io_ins_2(ces_13_0_io_ins_2),
    .io_ins_3(ces_13_0_io_ins_3),
    .io_outs_0(ces_13_0_io_outs_0),
    .io_outs_1(ces_13_0_io_outs_1),
    .io_outs_2(ces_13_0_io_outs_2),
    .io_outs_3(ces_13_0_io_outs_3)
  );
  Element ces_13_1 ( // @[MockArray.scala 37:53]
    .clock(ces_13_1_clock),
    .io_ins_0(ces_13_1_io_ins_0),
    .io_ins_1(ces_13_1_io_ins_1),
    .io_ins_2(ces_13_1_io_ins_2),
    .io_ins_3(ces_13_1_io_ins_3),
    .io_outs_0(ces_13_1_io_outs_0),
    .io_outs_1(ces_13_1_io_outs_1),
    .io_outs_2(ces_13_1_io_outs_2),
    .io_outs_3(ces_13_1_io_outs_3)
  );
  Element ces_13_2 ( // @[MockArray.scala 37:53]
    .clock(ces_13_2_clock),
    .io_ins_0(ces_13_2_io_ins_0),
    .io_ins_1(ces_13_2_io_ins_1),
    .io_ins_2(ces_13_2_io_ins_2),
    .io_ins_3(ces_13_2_io_ins_3),
    .io_outs_0(ces_13_2_io_outs_0),
    .io_outs_1(ces_13_2_io_outs_1),
    .io_outs_2(ces_13_2_io_outs_2),
    .io_outs_3(ces_13_2_io_outs_3)
  );
  Element ces_13_3 ( // @[MockArray.scala 37:53]
    .clock(ces_13_3_clock),
    .io_ins_0(ces_13_3_io_ins_0),
    .io_ins_1(ces_13_3_io_ins_1),
    .io_ins_2(ces_13_3_io_ins_2),
    .io_ins_3(ces_13_3_io_ins_3),
    .io_outs_0(ces_13_3_io_outs_0),
    .io_outs_1(ces_13_3_io_outs_1),
    .io_outs_2(ces_13_3_io_outs_2),
    .io_outs_3(ces_13_3_io_outs_3)
  );
  Element ces_13_4 ( // @[MockArray.scala 37:53]
    .clock(ces_13_4_clock),
    .io_ins_0(ces_13_4_io_ins_0),
    .io_ins_1(ces_13_4_io_ins_1),
    .io_ins_2(ces_13_4_io_ins_2),
    .io_ins_3(ces_13_4_io_ins_3),
    .io_outs_0(ces_13_4_io_outs_0),
    .io_outs_1(ces_13_4_io_outs_1),
    .io_outs_2(ces_13_4_io_outs_2),
    .io_outs_3(ces_13_4_io_outs_3)
  );
  Element ces_13_5 ( // @[MockArray.scala 37:53]
    .clock(ces_13_5_clock),
    .io_ins_0(ces_13_5_io_ins_0),
    .io_ins_1(ces_13_5_io_ins_1),
    .io_ins_2(ces_13_5_io_ins_2),
    .io_ins_3(ces_13_5_io_ins_3),
    .io_outs_0(ces_13_5_io_outs_0),
    .io_outs_1(ces_13_5_io_outs_1),
    .io_outs_2(ces_13_5_io_outs_2),
    .io_outs_3(ces_13_5_io_outs_3)
  );
  Element ces_13_6 ( // @[MockArray.scala 37:53]
    .clock(ces_13_6_clock),
    .io_ins_0(ces_13_6_io_ins_0),
    .io_ins_1(ces_13_6_io_ins_1),
    .io_ins_2(ces_13_6_io_ins_2),
    .io_ins_3(ces_13_6_io_ins_3),
    .io_outs_0(ces_13_6_io_outs_0),
    .io_outs_1(ces_13_6_io_outs_1),
    .io_outs_2(ces_13_6_io_outs_2),
    .io_outs_3(ces_13_6_io_outs_3)
  );
  Element ces_13_7 ( // @[MockArray.scala 37:53]
    .clock(ces_13_7_clock),
    .io_ins_0(ces_13_7_io_ins_0),
    .io_ins_1(ces_13_7_io_ins_1),
    .io_ins_2(ces_13_7_io_ins_2),
    .io_ins_3(ces_13_7_io_ins_3),
    .io_outs_0(ces_13_7_io_outs_0),
    .io_outs_1(ces_13_7_io_outs_1),
    .io_outs_2(ces_13_7_io_outs_2),
    .io_outs_3(ces_13_7_io_outs_3)
  );
  Element ces_13_8 ( // @[MockArray.scala 37:53]
    .clock(ces_13_8_clock),
    .io_ins_0(ces_13_8_io_ins_0),
    .io_ins_1(ces_13_8_io_ins_1),
    .io_ins_2(ces_13_8_io_ins_2),
    .io_ins_3(ces_13_8_io_ins_3),
    .io_outs_0(ces_13_8_io_outs_0),
    .io_outs_1(ces_13_8_io_outs_1),
    .io_outs_2(ces_13_8_io_outs_2),
    .io_outs_3(ces_13_8_io_outs_3)
  );
  Element ces_13_9 ( // @[MockArray.scala 37:53]
    .clock(ces_13_9_clock),
    .io_ins_0(ces_13_9_io_ins_0),
    .io_ins_1(ces_13_9_io_ins_1),
    .io_ins_2(ces_13_9_io_ins_2),
    .io_ins_3(ces_13_9_io_ins_3),
    .io_outs_0(ces_13_9_io_outs_0),
    .io_outs_1(ces_13_9_io_outs_1),
    .io_outs_2(ces_13_9_io_outs_2),
    .io_outs_3(ces_13_9_io_outs_3)
  );
  Element ces_13_10 ( // @[MockArray.scala 37:53]
    .clock(ces_13_10_clock),
    .io_ins_0(ces_13_10_io_ins_0),
    .io_ins_1(ces_13_10_io_ins_1),
    .io_ins_2(ces_13_10_io_ins_2),
    .io_ins_3(ces_13_10_io_ins_3),
    .io_outs_0(ces_13_10_io_outs_0),
    .io_outs_1(ces_13_10_io_outs_1),
    .io_outs_2(ces_13_10_io_outs_2),
    .io_outs_3(ces_13_10_io_outs_3)
  );
  Element ces_13_11 ( // @[MockArray.scala 37:53]
    .clock(ces_13_11_clock),
    .io_ins_0(ces_13_11_io_ins_0),
    .io_ins_1(ces_13_11_io_ins_1),
    .io_ins_2(ces_13_11_io_ins_2),
    .io_ins_3(ces_13_11_io_ins_3),
    .io_outs_0(ces_13_11_io_outs_0),
    .io_outs_1(ces_13_11_io_outs_1),
    .io_outs_2(ces_13_11_io_outs_2),
    .io_outs_3(ces_13_11_io_outs_3)
  );
  Element ces_13_12 ( // @[MockArray.scala 37:53]
    .clock(ces_13_12_clock),
    .io_ins_0(ces_13_12_io_ins_0),
    .io_ins_1(ces_13_12_io_ins_1),
    .io_ins_2(ces_13_12_io_ins_2),
    .io_ins_3(ces_13_12_io_ins_3),
    .io_outs_0(ces_13_12_io_outs_0),
    .io_outs_1(ces_13_12_io_outs_1),
    .io_outs_2(ces_13_12_io_outs_2),
    .io_outs_3(ces_13_12_io_outs_3)
  );
  Element ces_13_13 ( // @[MockArray.scala 37:53]
    .clock(ces_13_13_clock),
    .io_ins_0(ces_13_13_io_ins_0),
    .io_ins_1(ces_13_13_io_ins_1),
    .io_ins_2(ces_13_13_io_ins_2),
    .io_ins_3(ces_13_13_io_ins_3),
    .io_outs_0(ces_13_13_io_outs_0),
    .io_outs_1(ces_13_13_io_outs_1),
    .io_outs_2(ces_13_13_io_outs_2),
    .io_outs_3(ces_13_13_io_outs_3)
  );
  Element ces_13_14 ( // @[MockArray.scala 37:53]
    .clock(ces_13_14_clock),
    .io_ins_0(ces_13_14_io_ins_0),
    .io_ins_1(ces_13_14_io_ins_1),
    .io_ins_2(ces_13_14_io_ins_2),
    .io_ins_3(ces_13_14_io_ins_3),
    .io_outs_0(ces_13_14_io_outs_0),
    .io_outs_1(ces_13_14_io_outs_1),
    .io_outs_2(ces_13_14_io_outs_2),
    .io_outs_3(ces_13_14_io_outs_3)
  );
  Element ces_13_15 ( // @[MockArray.scala 37:53]
    .clock(ces_13_15_clock),
    .io_ins_0(ces_13_15_io_ins_0),
    .io_ins_1(ces_13_15_io_ins_1),
    .io_ins_2(ces_13_15_io_ins_2),
    .io_ins_3(ces_13_15_io_ins_3),
    .io_outs_0(ces_13_15_io_outs_0),
    .io_outs_1(ces_13_15_io_outs_1),
    .io_outs_2(ces_13_15_io_outs_2),
    .io_outs_3(ces_13_15_io_outs_3)
  );
  Element ces_14_0 ( // @[MockArray.scala 37:53]
    .clock(ces_14_0_clock),
    .io_ins_0(ces_14_0_io_ins_0),
    .io_ins_1(ces_14_0_io_ins_1),
    .io_ins_2(ces_14_0_io_ins_2),
    .io_ins_3(ces_14_0_io_ins_3),
    .io_outs_0(ces_14_0_io_outs_0),
    .io_outs_1(ces_14_0_io_outs_1),
    .io_outs_2(ces_14_0_io_outs_2),
    .io_outs_3(ces_14_0_io_outs_3)
  );
  Element ces_14_1 ( // @[MockArray.scala 37:53]
    .clock(ces_14_1_clock),
    .io_ins_0(ces_14_1_io_ins_0),
    .io_ins_1(ces_14_1_io_ins_1),
    .io_ins_2(ces_14_1_io_ins_2),
    .io_ins_3(ces_14_1_io_ins_3),
    .io_outs_0(ces_14_1_io_outs_0),
    .io_outs_1(ces_14_1_io_outs_1),
    .io_outs_2(ces_14_1_io_outs_2),
    .io_outs_3(ces_14_1_io_outs_3)
  );
  Element ces_14_2 ( // @[MockArray.scala 37:53]
    .clock(ces_14_2_clock),
    .io_ins_0(ces_14_2_io_ins_0),
    .io_ins_1(ces_14_2_io_ins_1),
    .io_ins_2(ces_14_2_io_ins_2),
    .io_ins_3(ces_14_2_io_ins_3),
    .io_outs_0(ces_14_2_io_outs_0),
    .io_outs_1(ces_14_2_io_outs_1),
    .io_outs_2(ces_14_2_io_outs_2),
    .io_outs_3(ces_14_2_io_outs_3)
  );
  Element ces_14_3 ( // @[MockArray.scala 37:53]
    .clock(ces_14_3_clock),
    .io_ins_0(ces_14_3_io_ins_0),
    .io_ins_1(ces_14_3_io_ins_1),
    .io_ins_2(ces_14_3_io_ins_2),
    .io_ins_3(ces_14_3_io_ins_3),
    .io_outs_0(ces_14_3_io_outs_0),
    .io_outs_1(ces_14_3_io_outs_1),
    .io_outs_2(ces_14_3_io_outs_2),
    .io_outs_3(ces_14_3_io_outs_3)
  );
  Element ces_14_4 ( // @[MockArray.scala 37:53]
    .clock(ces_14_4_clock),
    .io_ins_0(ces_14_4_io_ins_0),
    .io_ins_1(ces_14_4_io_ins_1),
    .io_ins_2(ces_14_4_io_ins_2),
    .io_ins_3(ces_14_4_io_ins_3),
    .io_outs_0(ces_14_4_io_outs_0),
    .io_outs_1(ces_14_4_io_outs_1),
    .io_outs_2(ces_14_4_io_outs_2),
    .io_outs_3(ces_14_4_io_outs_3)
  );
  Element ces_14_5 ( // @[MockArray.scala 37:53]
    .clock(ces_14_5_clock),
    .io_ins_0(ces_14_5_io_ins_0),
    .io_ins_1(ces_14_5_io_ins_1),
    .io_ins_2(ces_14_5_io_ins_2),
    .io_ins_3(ces_14_5_io_ins_3),
    .io_outs_0(ces_14_5_io_outs_0),
    .io_outs_1(ces_14_5_io_outs_1),
    .io_outs_2(ces_14_5_io_outs_2),
    .io_outs_3(ces_14_5_io_outs_3)
  );
  Element ces_14_6 ( // @[MockArray.scala 37:53]
    .clock(ces_14_6_clock),
    .io_ins_0(ces_14_6_io_ins_0),
    .io_ins_1(ces_14_6_io_ins_1),
    .io_ins_2(ces_14_6_io_ins_2),
    .io_ins_3(ces_14_6_io_ins_3),
    .io_outs_0(ces_14_6_io_outs_0),
    .io_outs_1(ces_14_6_io_outs_1),
    .io_outs_2(ces_14_6_io_outs_2),
    .io_outs_3(ces_14_6_io_outs_3)
  );
  Element ces_14_7 ( // @[MockArray.scala 37:53]
    .clock(ces_14_7_clock),
    .io_ins_0(ces_14_7_io_ins_0),
    .io_ins_1(ces_14_7_io_ins_1),
    .io_ins_2(ces_14_7_io_ins_2),
    .io_ins_3(ces_14_7_io_ins_3),
    .io_outs_0(ces_14_7_io_outs_0),
    .io_outs_1(ces_14_7_io_outs_1),
    .io_outs_2(ces_14_7_io_outs_2),
    .io_outs_3(ces_14_7_io_outs_3)
  );
  Element ces_14_8 ( // @[MockArray.scala 37:53]
    .clock(ces_14_8_clock),
    .io_ins_0(ces_14_8_io_ins_0),
    .io_ins_1(ces_14_8_io_ins_1),
    .io_ins_2(ces_14_8_io_ins_2),
    .io_ins_3(ces_14_8_io_ins_3),
    .io_outs_0(ces_14_8_io_outs_0),
    .io_outs_1(ces_14_8_io_outs_1),
    .io_outs_2(ces_14_8_io_outs_2),
    .io_outs_3(ces_14_8_io_outs_3)
  );
  Element ces_14_9 ( // @[MockArray.scala 37:53]
    .clock(ces_14_9_clock),
    .io_ins_0(ces_14_9_io_ins_0),
    .io_ins_1(ces_14_9_io_ins_1),
    .io_ins_2(ces_14_9_io_ins_2),
    .io_ins_3(ces_14_9_io_ins_3),
    .io_outs_0(ces_14_9_io_outs_0),
    .io_outs_1(ces_14_9_io_outs_1),
    .io_outs_2(ces_14_9_io_outs_2),
    .io_outs_3(ces_14_9_io_outs_3)
  );
  Element ces_14_10 ( // @[MockArray.scala 37:53]
    .clock(ces_14_10_clock),
    .io_ins_0(ces_14_10_io_ins_0),
    .io_ins_1(ces_14_10_io_ins_1),
    .io_ins_2(ces_14_10_io_ins_2),
    .io_ins_3(ces_14_10_io_ins_3),
    .io_outs_0(ces_14_10_io_outs_0),
    .io_outs_1(ces_14_10_io_outs_1),
    .io_outs_2(ces_14_10_io_outs_2),
    .io_outs_3(ces_14_10_io_outs_3)
  );
  Element ces_14_11 ( // @[MockArray.scala 37:53]
    .clock(ces_14_11_clock),
    .io_ins_0(ces_14_11_io_ins_0),
    .io_ins_1(ces_14_11_io_ins_1),
    .io_ins_2(ces_14_11_io_ins_2),
    .io_ins_3(ces_14_11_io_ins_3),
    .io_outs_0(ces_14_11_io_outs_0),
    .io_outs_1(ces_14_11_io_outs_1),
    .io_outs_2(ces_14_11_io_outs_2),
    .io_outs_3(ces_14_11_io_outs_3)
  );
  Element ces_14_12 ( // @[MockArray.scala 37:53]
    .clock(ces_14_12_clock),
    .io_ins_0(ces_14_12_io_ins_0),
    .io_ins_1(ces_14_12_io_ins_1),
    .io_ins_2(ces_14_12_io_ins_2),
    .io_ins_3(ces_14_12_io_ins_3),
    .io_outs_0(ces_14_12_io_outs_0),
    .io_outs_1(ces_14_12_io_outs_1),
    .io_outs_2(ces_14_12_io_outs_2),
    .io_outs_3(ces_14_12_io_outs_3)
  );
  Element ces_14_13 ( // @[MockArray.scala 37:53]
    .clock(ces_14_13_clock),
    .io_ins_0(ces_14_13_io_ins_0),
    .io_ins_1(ces_14_13_io_ins_1),
    .io_ins_2(ces_14_13_io_ins_2),
    .io_ins_3(ces_14_13_io_ins_3),
    .io_outs_0(ces_14_13_io_outs_0),
    .io_outs_1(ces_14_13_io_outs_1),
    .io_outs_2(ces_14_13_io_outs_2),
    .io_outs_3(ces_14_13_io_outs_3)
  );
  Element ces_14_14 ( // @[MockArray.scala 37:53]
    .clock(ces_14_14_clock),
    .io_ins_0(ces_14_14_io_ins_0),
    .io_ins_1(ces_14_14_io_ins_1),
    .io_ins_2(ces_14_14_io_ins_2),
    .io_ins_3(ces_14_14_io_ins_3),
    .io_outs_0(ces_14_14_io_outs_0),
    .io_outs_1(ces_14_14_io_outs_1),
    .io_outs_2(ces_14_14_io_outs_2),
    .io_outs_3(ces_14_14_io_outs_3)
  );
  Element ces_14_15 ( // @[MockArray.scala 37:53]
    .clock(ces_14_15_clock),
    .io_ins_0(ces_14_15_io_ins_0),
    .io_ins_1(ces_14_15_io_ins_1),
    .io_ins_2(ces_14_15_io_ins_2),
    .io_ins_3(ces_14_15_io_ins_3),
    .io_outs_0(ces_14_15_io_outs_0),
    .io_outs_1(ces_14_15_io_outs_1),
    .io_outs_2(ces_14_15_io_outs_2),
    .io_outs_3(ces_14_15_io_outs_3)
  );
  Element ces_15_0 ( // @[MockArray.scala 37:53]
    .clock(ces_15_0_clock),
    .io_ins_0(ces_15_0_io_ins_0),
    .io_ins_1(ces_15_0_io_ins_1),
    .io_ins_2(ces_15_0_io_ins_2),
    .io_ins_3(ces_15_0_io_ins_3),
    .io_outs_0(ces_15_0_io_outs_0),
    .io_outs_1(ces_15_0_io_outs_1),
    .io_outs_2(ces_15_0_io_outs_2),
    .io_outs_3(ces_15_0_io_outs_3)
  );
  Element ces_15_1 ( // @[MockArray.scala 37:53]
    .clock(ces_15_1_clock),
    .io_ins_0(ces_15_1_io_ins_0),
    .io_ins_1(ces_15_1_io_ins_1),
    .io_ins_2(ces_15_1_io_ins_2),
    .io_ins_3(ces_15_1_io_ins_3),
    .io_outs_0(ces_15_1_io_outs_0),
    .io_outs_1(ces_15_1_io_outs_1),
    .io_outs_2(ces_15_1_io_outs_2),
    .io_outs_3(ces_15_1_io_outs_3)
  );
  Element ces_15_2 ( // @[MockArray.scala 37:53]
    .clock(ces_15_2_clock),
    .io_ins_0(ces_15_2_io_ins_0),
    .io_ins_1(ces_15_2_io_ins_1),
    .io_ins_2(ces_15_2_io_ins_2),
    .io_ins_3(ces_15_2_io_ins_3),
    .io_outs_0(ces_15_2_io_outs_0),
    .io_outs_1(ces_15_2_io_outs_1),
    .io_outs_2(ces_15_2_io_outs_2),
    .io_outs_3(ces_15_2_io_outs_3)
  );
  Element ces_15_3 ( // @[MockArray.scala 37:53]
    .clock(ces_15_3_clock),
    .io_ins_0(ces_15_3_io_ins_0),
    .io_ins_1(ces_15_3_io_ins_1),
    .io_ins_2(ces_15_3_io_ins_2),
    .io_ins_3(ces_15_3_io_ins_3),
    .io_outs_0(ces_15_3_io_outs_0),
    .io_outs_1(ces_15_3_io_outs_1),
    .io_outs_2(ces_15_3_io_outs_2),
    .io_outs_3(ces_15_3_io_outs_3)
  );
  Element ces_15_4 ( // @[MockArray.scala 37:53]
    .clock(ces_15_4_clock),
    .io_ins_0(ces_15_4_io_ins_0),
    .io_ins_1(ces_15_4_io_ins_1),
    .io_ins_2(ces_15_4_io_ins_2),
    .io_ins_3(ces_15_4_io_ins_3),
    .io_outs_0(ces_15_4_io_outs_0),
    .io_outs_1(ces_15_4_io_outs_1),
    .io_outs_2(ces_15_4_io_outs_2),
    .io_outs_3(ces_15_4_io_outs_3)
  );
  Element ces_15_5 ( // @[MockArray.scala 37:53]
    .clock(ces_15_5_clock),
    .io_ins_0(ces_15_5_io_ins_0),
    .io_ins_1(ces_15_5_io_ins_1),
    .io_ins_2(ces_15_5_io_ins_2),
    .io_ins_3(ces_15_5_io_ins_3),
    .io_outs_0(ces_15_5_io_outs_0),
    .io_outs_1(ces_15_5_io_outs_1),
    .io_outs_2(ces_15_5_io_outs_2),
    .io_outs_3(ces_15_5_io_outs_3)
  );
  Element ces_15_6 ( // @[MockArray.scala 37:53]
    .clock(ces_15_6_clock),
    .io_ins_0(ces_15_6_io_ins_0),
    .io_ins_1(ces_15_6_io_ins_1),
    .io_ins_2(ces_15_6_io_ins_2),
    .io_ins_3(ces_15_6_io_ins_3),
    .io_outs_0(ces_15_6_io_outs_0),
    .io_outs_1(ces_15_6_io_outs_1),
    .io_outs_2(ces_15_6_io_outs_2),
    .io_outs_3(ces_15_6_io_outs_3)
  );
  Element ces_15_7 ( // @[MockArray.scala 37:53]
    .clock(ces_15_7_clock),
    .io_ins_0(ces_15_7_io_ins_0),
    .io_ins_1(ces_15_7_io_ins_1),
    .io_ins_2(ces_15_7_io_ins_2),
    .io_ins_3(ces_15_7_io_ins_3),
    .io_outs_0(ces_15_7_io_outs_0),
    .io_outs_1(ces_15_7_io_outs_1),
    .io_outs_2(ces_15_7_io_outs_2),
    .io_outs_3(ces_15_7_io_outs_3)
  );
  Element ces_15_8 ( // @[MockArray.scala 37:53]
    .clock(ces_15_8_clock),
    .io_ins_0(ces_15_8_io_ins_0),
    .io_ins_1(ces_15_8_io_ins_1),
    .io_ins_2(ces_15_8_io_ins_2),
    .io_ins_3(ces_15_8_io_ins_3),
    .io_outs_0(ces_15_8_io_outs_0),
    .io_outs_1(ces_15_8_io_outs_1),
    .io_outs_2(ces_15_8_io_outs_2),
    .io_outs_3(ces_15_8_io_outs_3)
  );
  Element ces_15_9 ( // @[MockArray.scala 37:53]
    .clock(ces_15_9_clock),
    .io_ins_0(ces_15_9_io_ins_0),
    .io_ins_1(ces_15_9_io_ins_1),
    .io_ins_2(ces_15_9_io_ins_2),
    .io_ins_3(ces_15_9_io_ins_3),
    .io_outs_0(ces_15_9_io_outs_0),
    .io_outs_1(ces_15_9_io_outs_1),
    .io_outs_2(ces_15_9_io_outs_2),
    .io_outs_3(ces_15_9_io_outs_3)
  );
  Element ces_15_10 ( // @[MockArray.scala 37:53]
    .clock(ces_15_10_clock),
    .io_ins_0(ces_15_10_io_ins_0),
    .io_ins_1(ces_15_10_io_ins_1),
    .io_ins_2(ces_15_10_io_ins_2),
    .io_ins_3(ces_15_10_io_ins_3),
    .io_outs_0(ces_15_10_io_outs_0),
    .io_outs_1(ces_15_10_io_outs_1),
    .io_outs_2(ces_15_10_io_outs_2),
    .io_outs_3(ces_15_10_io_outs_3)
  );
  Element ces_15_11 ( // @[MockArray.scala 37:53]
    .clock(ces_15_11_clock),
    .io_ins_0(ces_15_11_io_ins_0),
    .io_ins_1(ces_15_11_io_ins_1),
    .io_ins_2(ces_15_11_io_ins_2),
    .io_ins_3(ces_15_11_io_ins_3),
    .io_outs_0(ces_15_11_io_outs_0),
    .io_outs_1(ces_15_11_io_outs_1),
    .io_outs_2(ces_15_11_io_outs_2),
    .io_outs_3(ces_15_11_io_outs_3)
  );
  Element ces_15_12 ( // @[MockArray.scala 37:53]
    .clock(ces_15_12_clock),
    .io_ins_0(ces_15_12_io_ins_0),
    .io_ins_1(ces_15_12_io_ins_1),
    .io_ins_2(ces_15_12_io_ins_2),
    .io_ins_3(ces_15_12_io_ins_3),
    .io_outs_0(ces_15_12_io_outs_0),
    .io_outs_1(ces_15_12_io_outs_1),
    .io_outs_2(ces_15_12_io_outs_2),
    .io_outs_3(ces_15_12_io_outs_3)
  );
  Element ces_15_13 ( // @[MockArray.scala 37:53]
    .clock(ces_15_13_clock),
    .io_ins_0(ces_15_13_io_ins_0),
    .io_ins_1(ces_15_13_io_ins_1),
    .io_ins_2(ces_15_13_io_ins_2),
    .io_ins_3(ces_15_13_io_ins_3),
    .io_outs_0(ces_15_13_io_outs_0),
    .io_outs_1(ces_15_13_io_outs_1),
    .io_outs_2(ces_15_13_io_outs_2),
    .io_outs_3(ces_15_13_io_outs_3)
  );
  Element ces_15_14 ( // @[MockArray.scala 37:53]
    .clock(ces_15_14_clock),
    .io_ins_0(ces_15_14_io_ins_0),
    .io_ins_1(ces_15_14_io_ins_1),
    .io_ins_2(ces_15_14_io_ins_2),
    .io_ins_3(ces_15_14_io_ins_3),
    .io_outs_0(ces_15_14_io_outs_0),
    .io_outs_1(ces_15_14_io_outs_1),
    .io_outs_2(ces_15_14_io_outs_2),
    .io_outs_3(ces_15_14_io_outs_3)
  );
  Element ces_15_15 ( // @[MockArray.scala 37:53]
    .clock(ces_15_15_clock),
    .io_ins_0(ces_15_15_io_ins_0),
    .io_ins_1(ces_15_15_io_ins_1),
    .io_ins_2(ces_15_15_io_ins_2),
    .io_ins_3(ces_15_15_io_ins_3),
    .io_outs_0(ces_15_15_io_outs_0),
    .io_outs_1(ces_15_15_io_outs_1),
    .io_outs_2(ces_15_15_io_outs_2),
    .io_outs_3(ces_15_15_io_outs_3)
  );
  assign io_outsHorizontal_0_0 = ces_0_0_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_1 = ces_0_1_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_2 = ces_0_2_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_3 = ces_0_3_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_4 = ces_0_4_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_5 = ces_0_5_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_6 = ces_0_6_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_7 = ces_0_7_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_8 = ces_0_8_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_9 = ces_0_9_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_10 = ces_0_10_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_11 = ces_0_11_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_12 = ces_0_12_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_13 = ces_0_13_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_14 = ces_0_14_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_0_15 = ces_0_15_io_outs_0; // @[MockArray.scala 50:89]
  assign io_outsHorizontal_1_0 = ces_15_0_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_1 = ces_15_1_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_2 = ces_15_2_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_3 = ces_15_3_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_4 = ces_15_4_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_5 = ces_15_5_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_6 = ces_15_6_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_7 = ces_15_7_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_8 = ces_15_8_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_9 = ces_15_9_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_10 = ces_15_10_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_11 = ces_15_11_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_12 = ces_15_12_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_13 = ces_15_13_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_14 = ces_15_14_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsHorizontal_1_15 = ces_15_15_io_outs_2; // @[MockArray.scala 52:89]
  assign io_outsVertical_0_0 = ces_0_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_1 = ces_1_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_2 = ces_2_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_3 = ces_3_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_4 = ces_4_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_5 = ces_5_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_6 = ces_6_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_7 = ces_7_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_8 = ces_8_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_9 = ces_9_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_10 = ces_10_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_11 = ces_11_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_12 = ces_12_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_13 = ces_13_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_14 = ces_14_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_15 = ces_15_15_io_outs_1; // @[MockArray.scala 51:89]
  assign io_outsVertical_1_0 = ces_0_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_1 = ces_1_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_2 = ces_2_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_3 = ces_3_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_4 = ces_4_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_5 = ces_5_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_6 = ces_6_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_7 = ces_7_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_8 = ces_8_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_9 = ces_9_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_10 = ces_10_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_11 = ces_11_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_12 = ces_12_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_13 = ces_13_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_14 = ces_14_0_io_outs_3; // @[MockArray.scala 53:89]
  assign io_outsVertical_1_15 = ces_15_0_io_outs_3; // @[MockArray.scala 53:89]
  assign ces_0_0_clock = clock;
  assign ces_0_0_io_ins_0 = io_insHorizontal_0_0; // @[MockArray.scala 45:87]
  assign ces_0_0_io_ins_1 = ces_0_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_0_io_ins_2 = ces_1_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_0_io_ins_3 = io_insVertical_1_0; // @[MockArray.scala 48:87]
  assign ces_0_1_clock = clock;
  assign ces_0_1_io_ins_0 = io_insHorizontal_0_1; // @[MockArray.scala 45:87]
  assign ces_0_1_io_ins_1 = ces_0_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_1_io_ins_2 = ces_1_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_1_io_ins_3 = ces_0_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_2_clock = clock;
  assign ces_0_2_io_ins_0 = io_insHorizontal_0_2; // @[MockArray.scala 45:87]
  assign ces_0_2_io_ins_1 = ces_0_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_2_io_ins_2 = ces_1_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_2_io_ins_3 = ces_0_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_3_clock = clock;
  assign ces_0_3_io_ins_0 = io_insHorizontal_0_3; // @[MockArray.scala 45:87]
  assign ces_0_3_io_ins_1 = ces_0_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_3_io_ins_2 = ces_1_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_3_io_ins_3 = ces_0_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_4_clock = clock;
  assign ces_0_4_io_ins_0 = io_insHorizontal_0_4; // @[MockArray.scala 45:87]
  assign ces_0_4_io_ins_1 = ces_0_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_4_io_ins_2 = ces_1_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_4_io_ins_3 = ces_0_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_5_clock = clock;
  assign ces_0_5_io_ins_0 = io_insHorizontal_0_5; // @[MockArray.scala 45:87]
  assign ces_0_5_io_ins_1 = ces_0_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_5_io_ins_2 = ces_1_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_5_io_ins_3 = ces_0_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_6_clock = clock;
  assign ces_0_6_io_ins_0 = io_insHorizontal_0_6; // @[MockArray.scala 45:87]
  assign ces_0_6_io_ins_1 = ces_0_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_6_io_ins_2 = ces_1_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_6_io_ins_3 = ces_0_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_7_clock = clock;
  assign ces_0_7_io_ins_0 = io_insHorizontal_0_7; // @[MockArray.scala 45:87]
  assign ces_0_7_io_ins_1 = ces_0_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_7_io_ins_2 = ces_1_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_7_io_ins_3 = ces_0_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_8_clock = clock;
  assign ces_0_8_io_ins_0 = io_insHorizontal_0_8; // @[MockArray.scala 45:87]
  assign ces_0_8_io_ins_1 = ces_0_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_8_io_ins_2 = ces_1_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_8_io_ins_3 = ces_0_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_9_clock = clock;
  assign ces_0_9_io_ins_0 = io_insHorizontal_0_9; // @[MockArray.scala 45:87]
  assign ces_0_9_io_ins_1 = ces_0_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_9_io_ins_2 = ces_1_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_9_io_ins_3 = ces_0_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_10_clock = clock;
  assign ces_0_10_io_ins_0 = io_insHorizontal_0_10; // @[MockArray.scala 45:87]
  assign ces_0_10_io_ins_1 = ces_0_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_10_io_ins_2 = ces_1_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_10_io_ins_3 = ces_0_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_11_clock = clock;
  assign ces_0_11_io_ins_0 = io_insHorizontal_0_11; // @[MockArray.scala 45:87]
  assign ces_0_11_io_ins_1 = ces_0_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_11_io_ins_2 = ces_1_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_11_io_ins_3 = ces_0_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_12_clock = clock;
  assign ces_0_12_io_ins_0 = io_insHorizontal_0_12; // @[MockArray.scala 45:87]
  assign ces_0_12_io_ins_1 = ces_0_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_12_io_ins_2 = ces_1_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_12_io_ins_3 = ces_0_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_13_clock = clock;
  assign ces_0_13_io_ins_0 = io_insHorizontal_0_13; // @[MockArray.scala 45:87]
  assign ces_0_13_io_ins_1 = ces_0_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_13_io_ins_2 = ces_1_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_13_io_ins_3 = ces_0_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_14_clock = clock;
  assign ces_0_14_io_ins_0 = io_insHorizontal_0_14; // @[MockArray.scala 45:87]
  assign ces_0_14_io_ins_1 = ces_0_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_0_14_io_ins_2 = ces_1_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_14_io_ins_3 = ces_0_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_0_15_clock = clock;
  assign ces_0_15_io_ins_0 = io_insHorizontal_0_15; // @[MockArray.scala 45:87]
  assign ces_0_15_io_ins_1 = io_insVertical_0_0; // @[MockArray.scala 46:87]
  assign ces_0_15_io_ins_2 = ces_1_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_0_15_io_ins_3 = ces_0_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_0_clock = clock;
  assign ces_1_0_io_ins_0 = ces_0_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_0_io_ins_1 = ces_1_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_0_io_ins_2 = ces_2_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_0_io_ins_3 = io_insVertical_1_1; // @[MockArray.scala 48:87]
  assign ces_1_1_clock = clock;
  assign ces_1_1_io_ins_0 = ces_0_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_1_io_ins_1 = ces_1_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_1_io_ins_2 = ces_2_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_1_io_ins_3 = ces_1_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_2_clock = clock;
  assign ces_1_2_io_ins_0 = ces_0_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_2_io_ins_1 = ces_1_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_2_io_ins_2 = ces_2_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_2_io_ins_3 = ces_1_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_3_clock = clock;
  assign ces_1_3_io_ins_0 = ces_0_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_3_io_ins_1 = ces_1_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_3_io_ins_2 = ces_2_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_3_io_ins_3 = ces_1_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_4_clock = clock;
  assign ces_1_4_io_ins_0 = ces_0_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_4_io_ins_1 = ces_1_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_4_io_ins_2 = ces_2_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_4_io_ins_3 = ces_1_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_5_clock = clock;
  assign ces_1_5_io_ins_0 = ces_0_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_5_io_ins_1 = ces_1_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_5_io_ins_2 = ces_2_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_5_io_ins_3 = ces_1_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_6_clock = clock;
  assign ces_1_6_io_ins_0 = ces_0_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_6_io_ins_1 = ces_1_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_6_io_ins_2 = ces_2_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_6_io_ins_3 = ces_1_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_7_clock = clock;
  assign ces_1_7_io_ins_0 = ces_0_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_7_io_ins_1 = ces_1_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_7_io_ins_2 = ces_2_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_7_io_ins_3 = ces_1_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_8_clock = clock;
  assign ces_1_8_io_ins_0 = ces_0_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_8_io_ins_1 = ces_1_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_8_io_ins_2 = ces_2_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_8_io_ins_3 = ces_1_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_9_clock = clock;
  assign ces_1_9_io_ins_0 = ces_0_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_9_io_ins_1 = ces_1_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_9_io_ins_2 = ces_2_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_9_io_ins_3 = ces_1_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_10_clock = clock;
  assign ces_1_10_io_ins_0 = ces_0_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_10_io_ins_1 = ces_1_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_10_io_ins_2 = ces_2_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_10_io_ins_3 = ces_1_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_11_clock = clock;
  assign ces_1_11_io_ins_0 = ces_0_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_11_io_ins_1 = ces_1_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_11_io_ins_2 = ces_2_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_11_io_ins_3 = ces_1_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_12_clock = clock;
  assign ces_1_12_io_ins_0 = ces_0_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_12_io_ins_1 = ces_1_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_12_io_ins_2 = ces_2_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_12_io_ins_3 = ces_1_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_13_clock = clock;
  assign ces_1_13_io_ins_0 = ces_0_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_13_io_ins_1 = ces_1_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_13_io_ins_2 = ces_2_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_13_io_ins_3 = ces_1_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_14_clock = clock;
  assign ces_1_14_io_ins_0 = ces_0_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_14_io_ins_1 = ces_1_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_1_14_io_ins_2 = ces_2_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_14_io_ins_3 = ces_1_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_1_15_clock = clock;
  assign ces_1_15_io_ins_0 = ces_0_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_1_15_io_ins_1 = io_insVertical_0_1; // @[MockArray.scala 46:87]
  assign ces_1_15_io_ins_2 = ces_2_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_1_15_io_ins_3 = ces_1_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_0_clock = clock;
  assign ces_2_0_io_ins_0 = ces_1_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_0_io_ins_1 = ces_2_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_0_io_ins_2 = ces_3_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_0_io_ins_3 = io_insVertical_1_2; // @[MockArray.scala 48:87]
  assign ces_2_1_clock = clock;
  assign ces_2_1_io_ins_0 = ces_1_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_1_io_ins_1 = ces_2_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_1_io_ins_2 = ces_3_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_1_io_ins_3 = ces_2_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_2_clock = clock;
  assign ces_2_2_io_ins_0 = ces_1_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_2_io_ins_1 = ces_2_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_2_io_ins_2 = ces_3_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_2_io_ins_3 = ces_2_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_3_clock = clock;
  assign ces_2_3_io_ins_0 = ces_1_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_3_io_ins_1 = ces_2_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_3_io_ins_2 = ces_3_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_3_io_ins_3 = ces_2_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_4_clock = clock;
  assign ces_2_4_io_ins_0 = ces_1_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_4_io_ins_1 = ces_2_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_4_io_ins_2 = ces_3_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_4_io_ins_3 = ces_2_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_5_clock = clock;
  assign ces_2_5_io_ins_0 = ces_1_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_5_io_ins_1 = ces_2_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_5_io_ins_2 = ces_3_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_5_io_ins_3 = ces_2_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_6_clock = clock;
  assign ces_2_6_io_ins_0 = ces_1_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_6_io_ins_1 = ces_2_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_6_io_ins_2 = ces_3_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_6_io_ins_3 = ces_2_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_7_clock = clock;
  assign ces_2_7_io_ins_0 = ces_1_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_7_io_ins_1 = ces_2_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_7_io_ins_2 = ces_3_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_7_io_ins_3 = ces_2_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_8_clock = clock;
  assign ces_2_8_io_ins_0 = ces_1_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_8_io_ins_1 = ces_2_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_8_io_ins_2 = ces_3_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_8_io_ins_3 = ces_2_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_9_clock = clock;
  assign ces_2_9_io_ins_0 = ces_1_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_9_io_ins_1 = ces_2_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_9_io_ins_2 = ces_3_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_9_io_ins_3 = ces_2_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_10_clock = clock;
  assign ces_2_10_io_ins_0 = ces_1_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_10_io_ins_1 = ces_2_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_10_io_ins_2 = ces_3_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_10_io_ins_3 = ces_2_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_11_clock = clock;
  assign ces_2_11_io_ins_0 = ces_1_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_11_io_ins_1 = ces_2_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_11_io_ins_2 = ces_3_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_11_io_ins_3 = ces_2_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_12_clock = clock;
  assign ces_2_12_io_ins_0 = ces_1_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_12_io_ins_1 = ces_2_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_12_io_ins_2 = ces_3_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_12_io_ins_3 = ces_2_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_13_clock = clock;
  assign ces_2_13_io_ins_0 = ces_1_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_13_io_ins_1 = ces_2_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_13_io_ins_2 = ces_3_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_13_io_ins_3 = ces_2_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_14_clock = clock;
  assign ces_2_14_io_ins_0 = ces_1_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_14_io_ins_1 = ces_2_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_2_14_io_ins_2 = ces_3_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_14_io_ins_3 = ces_2_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_2_15_clock = clock;
  assign ces_2_15_io_ins_0 = ces_1_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_2_15_io_ins_1 = io_insVertical_0_2; // @[MockArray.scala 46:87]
  assign ces_2_15_io_ins_2 = ces_3_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_2_15_io_ins_3 = ces_2_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_0_clock = clock;
  assign ces_3_0_io_ins_0 = ces_2_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_0_io_ins_1 = ces_3_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_0_io_ins_2 = ces_4_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_0_io_ins_3 = io_insVertical_1_3; // @[MockArray.scala 48:87]
  assign ces_3_1_clock = clock;
  assign ces_3_1_io_ins_0 = ces_2_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_1_io_ins_1 = ces_3_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_1_io_ins_2 = ces_4_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_1_io_ins_3 = ces_3_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_2_clock = clock;
  assign ces_3_2_io_ins_0 = ces_2_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_2_io_ins_1 = ces_3_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_2_io_ins_2 = ces_4_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_2_io_ins_3 = ces_3_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_3_clock = clock;
  assign ces_3_3_io_ins_0 = ces_2_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_3_io_ins_1 = ces_3_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_3_io_ins_2 = ces_4_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_3_io_ins_3 = ces_3_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_4_clock = clock;
  assign ces_3_4_io_ins_0 = ces_2_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_4_io_ins_1 = ces_3_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_4_io_ins_2 = ces_4_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_4_io_ins_3 = ces_3_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_5_clock = clock;
  assign ces_3_5_io_ins_0 = ces_2_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_5_io_ins_1 = ces_3_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_5_io_ins_2 = ces_4_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_5_io_ins_3 = ces_3_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_6_clock = clock;
  assign ces_3_6_io_ins_0 = ces_2_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_6_io_ins_1 = ces_3_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_6_io_ins_2 = ces_4_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_6_io_ins_3 = ces_3_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_7_clock = clock;
  assign ces_3_7_io_ins_0 = ces_2_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_7_io_ins_1 = ces_3_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_7_io_ins_2 = ces_4_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_7_io_ins_3 = ces_3_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_8_clock = clock;
  assign ces_3_8_io_ins_0 = ces_2_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_8_io_ins_1 = ces_3_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_8_io_ins_2 = ces_4_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_8_io_ins_3 = ces_3_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_9_clock = clock;
  assign ces_3_9_io_ins_0 = ces_2_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_9_io_ins_1 = ces_3_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_9_io_ins_2 = ces_4_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_9_io_ins_3 = ces_3_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_10_clock = clock;
  assign ces_3_10_io_ins_0 = ces_2_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_10_io_ins_1 = ces_3_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_10_io_ins_2 = ces_4_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_10_io_ins_3 = ces_3_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_11_clock = clock;
  assign ces_3_11_io_ins_0 = ces_2_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_11_io_ins_1 = ces_3_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_11_io_ins_2 = ces_4_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_11_io_ins_3 = ces_3_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_12_clock = clock;
  assign ces_3_12_io_ins_0 = ces_2_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_12_io_ins_1 = ces_3_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_12_io_ins_2 = ces_4_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_12_io_ins_3 = ces_3_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_13_clock = clock;
  assign ces_3_13_io_ins_0 = ces_2_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_13_io_ins_1 = ces_3_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_13_io_ins_2 = ces_4_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_13_io_ins_3 = ces_3_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_14_clock = clock;
  assign ces_3_14_io_ins_0 = ces_2_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_14_io_ins_1 = ces_3_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_3_14_io_ins_2 = ces_4_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_14_io_ins_3 = ces_3_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_3_15_clock = clock;
  assign ces_3_15_io_ins_0 = ces_2_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_3_15_io_ins_1 = io_insVertical_0_3; // @[MockArray.scala 46:87]
  assign ces_3_15_io_ins_2 = ces_4_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_3_15_io_ins_3 = ces_3_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_0_clock = clock;
  assign ces_4_0_io_ins_0 = ces_3_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_0_io_ins_1 = ces_4_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_0_io_ins_2 = ces_5_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_0_io_ins_3 = io_insVertical_1_4; // @[MockArray.scala 48:87]
  assign ces_4_1_clock = clock;
  assign ces_4_1_io_ins_0 = ces_3_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_1_io_ins_1 = ces_4_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_1_io_ins_2 = ces_5_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_1_io_ins_3 = ces_4_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_2_clock = clock;
  assign ces_4_2_io_ins_0 = ces_3_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_2_io_ins_1 = ces_4_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_2_io_ins_2 = ces_5_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_2_io_ins_3 = ces_4_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_3_clock = clock;
  assign ces_4_3_io_ins_0 = ces_3_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_3_io_ins_1 = ces_4_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_3_io_ins_2 = ces_5_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_3_io_ins_3 = ces_4_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_4_clock = clock;
  assign ces_4_4_io_ins_0 = ces_3_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_4_io_ins_1 = ces_4_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_4_io_ins_2 = ces_5_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_4_io_ins_3 = ces_4_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_5_clock = clock;
  assign ces_4_5_io_ins_0 = ces_3_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_5_io_ins_1 = ces_4_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_5_io_ins_2 = ces_5_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_5_io_ins_3 = ces_4_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_6_clock = clock;
  assign ces_4_6_io_ins_0 = ces_3_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_6_io_ins_1 = ces_4_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_6_io_ins_2 = ces_5_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_6_io_ins_3 = ces_4_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_7_clock = clock;
  assign ces_4_7_io_ins_0 = ces_3_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_7_io_ins_1 = ces_4_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_7_io_ins_2 = ces_5_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_7_io_ins_3 = ces_4_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_8_clock = clock;
  assign ces_4_8_io_ins_0 = ces_3_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_8_io_ins_1 = ces_4_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_8_io_ins_2 = ces_5_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_8_io_ins_3 = ces_4_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_9_clock = clock;
  assign ces_4_9_io_ins_0 = ces_3_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_9_io_ins_1 = ces_4_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_9_io_ins_2 = ces_5_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_9_io_ins_3 = ces_4_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_10_clock = clock;
  assign ces_4_10_io_ins_0 = ces_3_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_10_io_ins_1 = ces_4_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_10_io_ins_2 = ces_5_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_10_io_ins_3 = ces_4_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_11_clock = clock;
  assign ces_4_11_io_ins_0 = ces_3_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_11_io_ins_1 = ces_4_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_11_io_ins_2 = ces_5_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_11_io_ins_3 = ces_4_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_12_clock = clock;
  assign ces_4_12_io_ins_0 = ces_3_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_12_io_ins_1 = ces_4_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_12_io_ins_2 = ces_5_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_12_io_ins_3 = ces_4_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_13_clock = clock;
  assign ces_4_13_io_ins_0 = ces_3_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_13_io_ins_1 = ces_4_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_13_io_ins_2 = ces_5_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_13_io_ins_3 = ces_4_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_14_clock = clock;
  assign ces_4_14_io_ins_0 = ces_3_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_14_io_ins_1 = ces_4_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_4_14_io_ins_2 = ces_5_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_14_io_ins_3 = ces_4_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_4_15_clock = clock;
  assign ces_4_15_io_ins_0 = ces_3_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_4_15_io_ins_1 = io_insVertical_0_4; // @[MockArray.scala 46:87]
  assign ces_4_15_io_ins_2 = ces_5_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_4_15_io_ins_3 = ces_4_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_0_clock = clock;
  assign ces_5_0_io_ins_0 = ces_4_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_0_io_ins_1 = ces_5_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_0_io_ins_2 = ces_6_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_0_io_ins_3 = io_insVertical_1_5; // @[MockArray.scala 48:87]
  assign ces_5_1_clock = clock;
  assign ces_5_1_io_ins_0 = ces_4_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_1_io_ins_1 = ces_5_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_1_io_ins_2 = ces_6_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_1_io_ins_3 = ces_5_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_2_clock = clock;
  assign ces_5_2_io_ins_0 = ces_4_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_2_io_ins_1 = ces_5_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_2_io_ins_2 = ces_6_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_2_io_ins_3 = ces_5_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_3_clock = clock;
  assign ces_5_3_io_ins_0 = ces_4_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_3_io_ins_1 = ces_5_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_3_io_ins_2 = ces_6_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_3_io_ins_3 = ces_5_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_4_clock = clock;
  assign ces_5_4_io_ins_0 = ces_4_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_4_io_ins_1 = ces_5_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_4_io_ins_2 = ces_6_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_4_io_ins_3 = ces_5_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_5_clock = clock;
  assign ces_5_5_io_ins_0 = ces_4_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_5_io_ins_1 = ces_5_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_5_io_ins_2 = ces_6_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_5_io_ins_3 = ces_5_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_6_clock = clock;
  assign ces_5_6_io_ins_0 = ces_4_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_6_io_ins_1 = ces_5_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_6_io_ins_2 = ces_6_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_6_io_ins_3 = ces_5_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_7_clock = clock;
  assign ces_5_7_io_ins_0 = ces_4_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_7_io_ins_1 = ces_5_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_7_io_ins_2 = ces_6_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_7_io_ins_3 = ces_5_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_8_clock = clock;
  assign ces_5_8_io_ins_0 = ces_4_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_8_io_ins_1 = ces_5_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_8_io_ins_2 = ces_6_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_8_io_ins_3 = ces_5_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_9_clock = clock;
  assign ces_5_9_io_ins_0 = ces_4_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_9_io_ins_1 = ces_5_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_9_io_ins_2 = ces_6_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_9_io_ins_3 = ces_5_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_10_clock = clock;
  assign ces_5_10_io_ins_0 = ces_4_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_10_io_ins_1 = ces_5_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_10_io_ins_2 = ces_6_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_10_io_ins_3 = ces_5_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_11_clock = clock;
  assign ces_5_11_io_ins_0 = ces_4_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_11_io_ins_1 = ces_5_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_11_io_ins_2 = ces_6_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_11_io_ins_3 = ces_5_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_12_clock = clock;
  assign ces_5_12_io_ins_0 = ces_4_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_12_io_ins_1 = ces_5_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_12_io_ins_2 = ces_6_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_12_io_ins_3 = ces_5_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_13_clock = clock;
  assign ces_5_13_io_ins_0 = ces_4_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_13_io_ins_1 = ces_5_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_13_io_ins_2 = ces_6_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_13_io_ins_3 = ces_5_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_14_clock = clock;
  assign ces_5_14_io_ins_0 = ces_4_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_14_io_ins_1 = ces_5_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_5_14_io_ins_2 = ces_6_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_14_io_ins_3 = ces_5_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_5_15_clock = clock;
  assign ces_5_15_io_ins_0 = ces_4_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_5_15_io_ins_1 = io_insVertical_0_5; // @[MockArray.scala 46:87]
  assign ces_5_15_io_ins_2 = ces_6_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_5_15_io_ins_3 = ces_5_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_0_clock = clock;
  assign ces_6_0_io_ins_0 = ces_5_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_0_io_ins_1 = ces_6_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_0_io_ins_2 = ces_7_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_0_io_ins_3 = io_insVertical_1_6; // @[MockArray.scala 48:87]
  assign ces_6_1_clock = clock;
  assign ces_6_1_io_ins_0 = ces_5_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_1_io_ins_1 = ces_6_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_1_io_ins_2 = ces_7_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_1_io_ins_3 = ces_6_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_2_clock = clock;
  assign ces_6_2_io_ins_0 = ces_5_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_2_io_ins_1 = ces_6_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_2_io_ins_2 = ces_7_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_2_io_ins_3 = ces_6_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_3_clock = clock;
  assign ces_6_3_io_ins_0 = ces_5_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_3_io_ins_1 = ces_6_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_3_io_ins_2 = ces_7_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_3_io_ins_3 = ces_6_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_4_clock = clock;
  assign ces_6_4_io_ins_0 = ces_5_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_4_io_ins_1 = ces_6_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_4_io_ins_2 = ces_7_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_4_io_ins_3 = ces_6_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_5_clock = clock;
  assign ces_6_5_io_ins_0 = ces_5_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_5_io_ins_1 = ces_6_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_5_io_ins_2 = ces_7_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_5_io_ins_3 = ces_6_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_6_clock = clock;
  assign ces_6_6_io_ins_0 = ces_5_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_6_io_ins_1 = ces_6_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_6_io_ins_2 = ces_7_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_6_io_ins_3 = ces_6_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_7_clock = clock;
  assign ces_6_7_io_ins_0 = ces_5_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_7_io_ins_1 = ces_6_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_7_io_ins_2 = ces_7_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_7_io_ins_3 = ces_6_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_8_clock = clock;
  assign ces_6_8_io_ins_0 = ces_5_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_8_io_ins_1 = ces_6_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_8_io_ins_2 = ces_7_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_8_io_ins_3 = ces_6_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_9_clock = clock;
  assign ces_6_9_io_ins_0 = ces_5_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_9_io_ins_1 = ces_6_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_9_io_ins_2 = ces_7_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_9_io_ins_3 = ces_6_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_10_clock = clock;
  assign ces_6_10_io_ins_0 = ces_5_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_10_io_ins_1 = ces_6_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_10_io_ins_2 = ces_7_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_10_io_ins_3 = ces_6_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_11_clock = clock;
  assign ces_6_11_io_ins_0 = ces_5_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_11_io_ins_1 = ces_6_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_11_io_ins_2 = ces_7_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_11_io_ins_3 = ces_6_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_12_clock = clock;
  assign ces_6_12_io_ins_0 = ces_5_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_12_io_ins_1 = ces_6_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_12_io_ins_2 = ces_7_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_12_io_ins_3 = ces_6_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_13_clock = clock;
  assign ces_6_13_io_ins_0 = ces_5_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_13_io_ins_1 = ces_6_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_13_io_ins_2 = ces_7_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_13_io_ins_3 = ces_6_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_14_clock = clock;
  assign ces_6_14_io_ins_0 = ces_5_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_14_io_ins_1 = ces_6_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_6_14_io_ins_2 = ces_7_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_14_io_ins_3 = ces_6_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_6_15_clock = clock;
  assign ces_6_15_io_ins_0 = ces_5_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_6_15_io_ins_1 = io_insVertical_0_6; // @[MockArray.scala 46:87]
  assign ces_6_15_io_ins_2 = ces_7_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_6_15_io_ins_3 = ces_6_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_0_clock = clock;
  assign ces_7_0_io_ins_0 = ces_6_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_0_io_ins_1 = ces_7_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_0_io_ins_2 = ces_8_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_0_io_ins_3 = io_insVertical_1_7; // @[MockArray.scala 48:87]
  assign ces_7_1_clock = clock;
  assign ces_7_1_io_ins_0 = ces_6_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_1_io_ins_1 = ces_7_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_1_io_ins_2 = ces_8_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_1_io_ins_3 = ces_7_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_2_clock = clock;
  assign ces_7_2_io_ins_0 = ces_6_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_2_io_ins_1 = ces_7_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_2_io_ins_2 = ces_8_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_2_io_ins_3 = ces_7_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_3_clock = clock;
  assign ces_7_3_io_ins_0 = ces_6_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_3_io_ins_1 = ces_7_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_3_io_ins_2 = ces_8_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_3_io_ins_3 = ces_7_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_4_clock = clock;
  assign ces_7_4_io_ins_0 = ces_6_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_4_io_ins_1 = ces_7_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_4_io_ins_2 = ces_8_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_4_io_ins_3 = ces_7_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_5_clock = clock;
  assign ces_7_5_io_ins_0 = ces_6_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_5_io_ins_1 = ces_7_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_5_io_ins_2 = ces_8_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_5_io_ins_3 = ces_7_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_6_clock = clock;
  assign ces_7_6_io_ins_0 = ces_6_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_6_io_ins_1 = ces_7_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_6_io_ins_2 = ces_8_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_6_io_ins_3 = ces_7_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_7_clock = clock;
  assign ces_7_7_io_ins_0 = ces_6_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_7_io_ins_1 = ces_7_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_7_io_ins_2 = ces_8_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_7_io_ins_3 = ces_7_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_8_clock = clock;
  assign ces_7_8_io_ins_0 = ces_6_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_8_io_ins_1 = ces_7_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_8_io_ins_2 = ces_8_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_8_io_ins_3 = ces_7_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_9_clock = clock;
  assign ces_7_9_io_ins_0 = ces_6_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_9_io_ins_1 = ces_7_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_9_io_ins_2 = ces_8_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_9_io_ins_3 = ces_7_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_10_clock = clock;
  assign ces_7_10_io_ins_0 = ces_6_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_10_io_ins_1 = ces_7_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_10_io_ins_2 = ces_8_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_10_io_ins_3 = ces_7_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_11_clock = clock;
  assign ces_7_11_io_ins_0 = ces_6_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_11_io_ins_1 = ces_7_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_11_io_ins_2 = ces_8_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_11_io_ins_3 = ces_7_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_12_clock = clock;
  assign ces_7_12_io_ins_0 = ces_6_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_12_io_ins_1 = ces_7_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_12_io_ins_2 = ces_8_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_12_io_ins_3 = ces_7_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_13_clock = clock;
  assign ces_7_13_io_ins_0 = ces_6_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_13_io_ins_1 = ces_7_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_13_io_ins_2 = ces_8_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_13_io_ins_3 = ces_7_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_14_clock = clock;
  assign ces_7_14_io_ins_0 = ces_6_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_14_io_ins_1 = ces_7_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_7_14_io_ins_2 = ces_8_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_14_io_ins_3 = ces_7_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_7_15_clock = clock;
  assign ces_7_15_io_ins_0 = ces_6_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_7_15_io_ins_1 = io_insVertical_0_7; // @[MockArray.scala 46:87]
  assign ces_7_15_io_ins_2 = ces_8_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_7_15_io_ins_3 = ces_7_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_0_clock = clock;
  assign ces_8_0_io_ins_0 = ces_7_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_0_io_ins_1 = ces_8_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_0_io_ins_2 = ces_9_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_0_io_ins_3 = io_insVertical_1_8; // @[MockArray.scala 48:87]
  assign ces_8_1_clock = clock;
  assign ces_8_1_io_ins_0 = ces_7_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_1_io_ins_1 = ces_8_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_1_io_ins_2 = ces_9_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_1_io_ins_3 = ces_8_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_2_clock = clock;
  assign ces_8_2_io_ins_0 = ces_7_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_2_io_ins_1 = ces_8_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_2_io_ins_2 = ces_9_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_2_io_ins_3 = ces_8_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_3_clock = clock;
  assign ces_8_3_io_ins_0 = ces_7_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_3_io_ins_1 = ces_8_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_3_io_ins_2 = ces_9_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_3_io_ins_3 = ces_8_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_4_clock = clock;
  assign ces_8_4_io_ins_0 = ces_7_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_4_io_ins_1 = ces_8_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_4_io_ins_2 = ces_9_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_4_io_ins_3 = ces_8_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_5_clock = clock;
  assign ces_8_5_io_ins_0 = ces_7_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_5_io_ins_1 = ces_8_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_5_io_ins_2 = ces_9_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_5_io_ins_3 = ces_8_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_6_clock = clock;
  assign ces_8_6_io_ins_0 = ces_7_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_6_io_ins_1 = ces_8_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_6_io_ins_2 = ces_9_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_6_io_ins_3 = ces_8_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_7_clock = clock;
  assign ces_8_7_io_ins_0 = ces_7_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_7_io_ins_1 = ces_8_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_7_io_ins_2 = ces_9_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_7_io_ins_3 = ces_8_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_8_clock = clock;
  assign ces_8_8_io_ins_0 = ces_7_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_8_io_ins_1 = ces_8_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_8_io_ins_2 = ces_9_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_8_io_ins_3 = ces_8_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_9_clock = clock;
  assign ces_8_9_io_ins_0 = ces_7_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_9_io_ins_1 = ces_8_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_9_io_ins_2 = ces_9_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_9_io_ins_3 = ces_8_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_10_clock = clock;
  assign ces_8_10_io_ins_0 = ces_7_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_10_io_ins_1 = ces_8_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_10_io_ins_2 = ces_9_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_10_io_ins_3 = ces_8_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_11_clock = clock;
  assign ces_8_11_io_ins_0 = ces_7_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_11_io_ins_1 = ces_8_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_11_io_ins_2 = ces_9_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_11_io_ins_3 = ces_8_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_12_clock = clock;
  assign ces_8_12_io_ins_0 = ces_7_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_12_io_ins_1 = ces_8_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_12_io_ins_2 = ces_9_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_12_io_ins_3 = ces_8_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_13_clock = clock;
  assign ces_8_13_io_ins_0 = ces_7_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_13_io_ins_1 = ces_8_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_13_io_ins_2 = ces_9_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_13_io_ins_3 = ces_8_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_14_clock = clock;
  assign ces_8_14_io_ins_0 = ces_7_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_14_io_ins_1 = ces_8_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_8_14_io_ins_2 = ces_9_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_14_io_ins_3 = ces_8_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_8_15_clock = clock;
  assign ces_8_15_io_ins_0 = ces_7_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_8_15_io_ins_1 = io_insVertical_0_8; // @[MockArray.scala 46:87]
  assign ces_8_15_io_ins_2 = ces_9_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_8_15_io_ins_3 = ces_8_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_0_clock = clock;
  assign ces_9_0_io_ins_0 = ces_8_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_0_io_ins_1 = ces_9_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_0_io_ins_2 = ces_10_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_0_io_ins_3 = io_insVertical_1_9; // @[MockArray.scala 48:87]
  assign ces_9_1_clock = clock;
  assign ces_9_1_io_ins_0 = ces_8_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_1_io_ins_1 = ces_9_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_1_io_ins_2 = ces_10_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_1_io_ins_3 = ces_9_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_2_clock = clock;
  assign ces_9_2_io_ins_0 = ces_8_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_2_io_ins_1 = ces_9_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_2_io_ins_2 = ces_10_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_2_io_ins_3 = ces_9_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_3_clock = clock;
  assign ces_9_3_io_ins_0 = ces_8_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_3_io_ins_1 = ces_9_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_3_io_ins_2 = ces_10_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_3_io_ins_3 = ces_9_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_4_clock = clock;
  assign ces_9_4_io_ins_0 = ces_8_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_4_io_ins_1 = ces_9_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_4_io_ins_2 = ces_10_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_4_io_ins_3 = ces_9_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_5_clock = clock;
  assign ces_9_5_io_ins_0 = ces_8_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_5_io_ins_1 = ces_9_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_5_io_ins_2 = ces_10_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_5_io_ins_3 = ces_9_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_6_clock = clock;
  assign ces_9_6_io_ins_0 = ces_8_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_6_io_ins_1 = ces_9_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_6_io_ins_2 = ces_10_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_6_io_ins_3 = ces_9_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_7_clock = clock;
  assign ces_9_7_io_ins_0 = ces_8_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_7_io_ins_1 = ces_9_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_7_io_ins_2 = ces_10_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_7_io_ins_3 = ces_9_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_8_clock = clock;
  assign ces_9_8_io_ins_0 = ces_8_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_8_io_ins_1 = ces_9_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_8_io_ins_2 = ces_10_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_8_io_ins_3 = ces_9_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_9_clock = clock;
  assign ces_9_9_io_ins_0 = ces_8_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_9_io_ins_1 = ces_9_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_9_io_ins_2 = ces_10_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_9_io_ins_3 = ces_9_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_10_clock = clock;
  assign ces_9_10_io_ins_0 = ces_8_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_10_io_ins_1 = ces_9_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_10_io_ins_2 = ces_10_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_10_io_ins_3 = ces_9_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_11_clock = clock;
  assign ces_9_11_io_ins_0 = ces_8_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_11_io_ins_1 = ces_9_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_11_io_ins_2 = ces_10_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_11_io_ins_3 = ces_9_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_12_clock = clock;
  assign ces_9_12_io_ins_0 = ces_8_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_12_io_ins_1 = ces_9_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_12_io_ins_2 = ces_10_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_12_io_ins_3 = ces_9_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_13_clock = clock;
  assign ces_9_13_io_ins_0 = ces_8_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_13_io_ins_1 = ces_9_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_13_io_ins_2 = ces_10_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_13_io_ins_3 = ces_9_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_14_clock = clock;
  assign ces_9_14_io_ins_0 = ces_8_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_14_io_ins_1 = ces_9_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_9_14_io_ins_2 = ces_10_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_14_io_ins_3 = ces_9_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_9_15_clock = clock;
  assign ces_9_15_io_ins_0 = ces_8_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_9_15_io_ins_1 = io_insVertical_0_9; // @[MockArray.scala 46:87]
  assign ces_9_15_io_ins_2 = ces_10_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_9_15_io_ins_3 = ces_9_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_0_clock = clock;
  assign ces_10_0_io_ins_0 = ces_9_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_0_io_ins_1 = ces_10_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_0_io_ins_2 = ces_11_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_0_io_ins_3 = io_insVertical_1_10; // @[MockArray.scala 48:87]
  assign ces_10_1_clock = clock;
  assign ces_10_1_io_ins_0 = ces_9_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_1_io_ins_1 = ces_10_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_1_io_ins_2 = ces_11_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_1_io_ins_3 = ces_10_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_2_clock = clock;
  assign ces_10_2_io_ins_0 = ces_9_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_2_io_ins_1 = ces_10_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_2_io_ins_2 = ces_11_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_2_io_ins_3 = ces_10_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_3_clock = clock;
  assign ces_10_3_io_ins_0 = ces_9_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_3_io_ins_1 = ces_10_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_3_io_ins_2 = ces_11_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_3_io_ins_3 = ces_10_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_4_clock = clock;
  assign ces_10_4_io_ins_0 = ces_9_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_4_io_ins_1 = ces_10_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_4_io_ins_2 = ces_11_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_4_io_ins_3 = ces_10_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_5_clock = clock;
  assign ces_10_5_io_ins_0 = ces_9_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_5_io_ins_1 = ces_10_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_5_io_ins_2 = ces_11_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_5_io_ins_3 = ces_10_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_6_clock = clock;
  assign ces_10_6_io_ins_0 = ces_9_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_6_io_ins_1 = ces_10_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_6_io_ins_2 = ces_11_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_6_io_ins_3 = ces_10_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_7_clock = clock;
  assign ces_10_7_io_ins_0 = ces_9_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_7_io_ins_1 = ces_10_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_7_io_ins_2 = ces_11_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_7_io_ins_3 = ces_10_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_8_clock = clock;
  assign ces_10_8_io_ins_0 = ces_9_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_8_io_ins_1 = ces_10_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_8_io_ins_2 = ces_11_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_8_io_ins_3 = ces_10_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_9_clock = clock;
  assign ces_10_9_io_ins_0 = ces_9_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_9_io_ins_1 = ces_10_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_9_io_ins_2 = ces_11_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_9_io_ins_3 = ces_10_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_10_clock = clock;
  assign ces_10_10_io_ins_0 = ces_9_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_10_io_ins_1 = ces_10_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_10_io_ins_2 = ces_11_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_10_io_ins_3 = ces_10_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_11_clock = clock;
  assign ces_10_11_io_ins_0 = ces_9_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_11_io_ins_1 = ces_10_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_11_io_ins_2 = ces_11_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_11_io_ins_3 = ces_10_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_12_clock = clock;
  assign ces_10_12_io_ins_0 = ces_9_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_12_io_ins_1 = ces_10_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_12_io_ins_2 = ces_11_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_12_io_ins_3 = ces_10_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_13_clock = clock;
  assign ces_10_13_io_ins_0 = ces_9_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_13_io_ins_1 = ces_10_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_13_io_ins_2 = ces_11_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_13_io_ins_3 = ces_10_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_14_clock = clock;
  assign ces_10_14_io_ins_0 = ces_9_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_14_io_ins_1 = ces_10_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_10_14_io_ins_2 = ces_11_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_14_io_ins_3 = ces_10_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_10_15_clock = clock;
  assign ces_10_15_io_ins_0 = ces_9_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_10_15_io_ins_1 = io_insVertical_0_10; // @[MockArray.scala 46:87]
  assign ces_10_15_io_ins_2 = ces_11_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_10_15_io_ins_3 = ces_10_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_0_clock = clock;
  assign ces_11_0_io_ins_0 = ces_10_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_0_io_ins_1 = ces_11_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_0_io_ins_2 = ces_12_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_0_io_ins_3 = io_insVertical_1_11; // @[MockArray.scala 48:87]
  assign ces_11_1_clock = clock;
  assign ces_11_1_io_ins_0 = ces_10_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_1_io_ins_1 = ces_11_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_1_io_ins_2 = ces_12_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_1_io_ins_3 = ces_11_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_2_clock = clock;
  assign ces_11_2_io_ins_0 = ces_10_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_2_io_ins_1 = ces_11_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_2_io_ins_2 = ces_12_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_2_io_ins_3 = ces_11_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_3_clock = clock;
  assign ces_11_3_io_ins_0 = ces_10_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_3_io_ins_1 = ces_11_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_3_io_ins_2 = ces_12_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_3_io_ins_3 = ces_11_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_4_clock = clock;
  assign ces_11_4_io_ins_0 = ces_10_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_4_io_ins_1 = ces_11_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_4_io_ins_2 = ces_12_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_4_io_ins_3 = ces_11_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_5_clock = clock;
  assign ces_11_5_io_ins_0 = ces_10_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_5_io_ins_1 = ces_11_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_5_io_ins_2 = ces_12_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_5_io_ins_3 = ces_11_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_6_clock = clock;
  assign ces_11_6_io_ins_0 = ces_10_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_6_io_ins_1 = ces_11_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_6_io_ins_2 = ces_12_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_6_io_ins_3 = ces_11_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_7_clock = clock;
  assign ces_11_7_io_ins_0 = ces_10_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_7_io_ins_1 = ces_11_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_7_io_ins_2 = ces_12_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_7_io_ins_3 = ces_11_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_8_clock = clock;
  assign ces_11_8_io_ins_0 = ces_10_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_8_io_ins_1 = ces_11_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_8_io_ins_2 = ces_12_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_8_io_ins_3 = ces_11_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_9_clock = clock;
  assign ces_11_9_io_ins_0 = ces_10_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_9_io_ins_1 = ces_11_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_9_io_ins_2 = ces_12_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_9_io_ins_3 = ces_11_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_10_clock = clock;
  assign ces_11_10_io_ins_0 = ces_10_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_10_io_ins_1 = ces_11_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_10_io_ins_2 = ces_12_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_10_io_ins_3 = ces_11_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_11_clock = clock;
  assign ces_11_11_io_ins_0 = ces_10_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_11_io_ins_1 = ces_11_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_11_io_ins_2 = ces_12_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_11_io_ins_3 = ces_11_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_12_clock = clock;
  assign ces_11_12_io_ins_0 = ces_10_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_12_io_ins_1 = ces_11_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_12_io_ins_2 = ces_12_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_12_io_ins_3 = ces_11_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_13_clock = clock;
  assign ces_11_13_io_ins_0 = ces_10_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_13_io_ins_1 = ces_11_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_13_io_ins_2 = ces_12_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_13_io_ins_3 = ces_11_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_14_clock = clock;
  assign ces_11_14_io_ins_0 = ces_10_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_14_io_ins_1 = ces_11_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_11_14_io_ins_2 = ces_12_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_14_io_ins_3 = ces_11_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_11_15_clock = clock;
  assign ces_11_15_io_ins_0 = ces_10_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_11_15_io_ins_1 = io_insVertical_0_11; // @[MockArray.scala 46:87]
  assign ces_11_15_io_ins_2 = ces_12_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_11_15_io_ins_3 = ces_11_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_0_clock = clock;
  assign ces_12_0_io_ins_0 = ces_11_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_0_io_ins_1 = ces_12_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_0_io_ins_2 = ces_13_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_0_io_ins_3 = io_insVertical_1_12; // @[MockArray.scala 48:87]
  assign ces_12_1_clock = clock;
  assign ces_12_1_io_ins_0 = ces_11_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_1_io_ins_1 = ces_12_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_1_io_ins_2 = ces_13_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_1_io_ins_3 = ces_12_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_2_clock = clock;
  assign ces_12_2_io_ins_0 = ces_11_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_2_io_ins_1 = ces_12_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_2_io_ins_2 = ces_13_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_2_io_ins_3 = ces_12_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_3_clock = clock;
  assign ces_12_3_io_ins_0 = ces_11_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_3_io_ins_1 = ces_12_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_3_io_ins_2 = ces_13_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_3_io_ins_3 = ces_12_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_4_clock = clock;
  assign ces_12_4_io_ins_0 = ces_11_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_4_io_ins_1 = ces_12_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_4_io_ins_2 = ces_13_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_4_io_ins_3 = ces_12_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_5_clock = clock;
  assign ces_12_5_io_ins_0 = ces_11_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_5_io_ins_1 = ces_12_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_5_io_ins_2 = ces_13_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_5_io_ins_3 = ces_12_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_6_clock = clock;
  assign ces_12_6_io_ins_0 = ces_11_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_6_io_ins_1 = ces_12_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_6_io_ins_2 = ces_13_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_6_io_ins_3 = ces_12_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_7_clock = clock;
  assign ces_12_7_io_ins_0 = ces_11_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_7_io_ins_1 = ces_12_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_7_io_ins_2 = ces_13_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_7_io_ins_3 = ces_12_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_8_clock = clock;
  assign ces_12_8_io_ins_0 = ces_11_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_8_io_ins_1 = ces_12_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_8_io_ins_2 = ces_13_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_8_io_ins_3 = ces_12_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_9_clock = clock;
  assign ces_12_9_io_ins_0 = ces_11_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_9_io_ins_1 = ces_12_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_9_io_ins_2 = ces_13_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_9_io_ins_3 = ces_12_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_10_clock = clock;
  assign ces_12_10_io_ins_0 = ces_11_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_10_io_ins_1 = ces_12_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_10_io_ins_2 = ces_13_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_10_io_ins_3 = ces_12_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_11_clock = clock;
  assign ces_12_11_io_ins_0 = ces_11_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_11_io_ins_1 = ces_12_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_11_io_ins_2 = ces_13_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_11_io_ins_3 = ces_12_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_12_clock = clock;
  assign ces_12_12_io_ins_0 = ces_11_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_12_io_ins_1 = ces_12_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_12_io_ins_2 = ces_13_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_12_io_ins_3 = ces_12_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_13_clock = clock;
  assign ces_12_13_io_ins_0 = ces_11_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_13_io_ins_1 = ces_12_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_13_io_ins_2 = ces_13_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_13_io_ins_3 = ces_12_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_14_clock = clock;
  assign ces_12_14_io_ins_0 = ces_11_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_14_io_ins_1 = ces_12_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_12_14_io_ins_2 = ces_13_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_14_io_ins_3 = ces_12_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_12_15_clock = clock;
  assign ces_12_15_io_ins_0 = ces_11_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_12_15_io_ins_1 = io_insVertical_0_12; // @[MockArray.scala 46:87]
  assign ces_12_15_io_ins_2 = ces_13_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_12_15_io_ins_3 = ces_12_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_0_clock = clock;
  assign ces_13_0_io_ins_0 = ces_12_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_0_io_ins_1 = ces_13_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_0_io_ins_2 = ces_14_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_0_io_ins_3 = io_insVertical_1_13; // @[MockArray.scala 48:87]
  assign ces_13_1_clock = clock;
  assign ces_13_1_io_ins_0 = ces_12_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_1_io_ins_1 = ces_13_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_1_io_ins_2 = ces_14_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_1_io_ins_3 = ces_13_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_2_clock = clock;
  assign ces_13_2_io_ins_0 = ces_12_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_2_io_ins_1 = ces_13_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_2_io_ins_2 = ces_14_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_2_io_ins_3 = ces_13_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_3_clock = clock;
  assign ces_13_3_io_ins_0 = ces_12_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_3_io_ins_1 = ces_13_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_3_io_ins_2 = ces_14_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_3_io_ins_3 = ces_13_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_4_clock = clock;
  assign ces_13_4_io_ins_0 = ces_12_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_4_io_ins_1 = ces_13_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_4_io_ins_2 = ces_14_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_4_io_ins_3 = ces_13_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_5_clock = clock;
  assign ces_13_5_io_ins_0 = ces_12_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_5_io_ins_1 = ces_13_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_5_io_ins_2 = ces_14_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_5_io_ins_3 = ces_13_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_6_clock = clock;
  assign ces_13_6_io_ins_0 = ces_12_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_6_io_ins_1 = ces_13_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_6_io_ins_2 = ces_14_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_6_io_ins_3 = ces_13_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_7_clock = clock;
  assign ces_13_7_io_ins_0 = ces_12_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_7_io_ins_1 = ces_13_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_7_io_ins_2 = ces_14_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_7_io_ins_3 = ces_13_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_8_clock = clock;
  assign ces_13_8_io_ins_0 = ces_12_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_8_io_ins_1 = ces_13_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_8_io_ins_2 = ces_14_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_8_io_ins_3 = ces_13_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_9_clock = clock;
  assign ces_13_9_io_ins_0 = ces_12_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_9_io_ins_1 = ces_13_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_9_io_ins_2 = ces_14_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_9_io_ins_3 = ces_13_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_10_clock = clock;
  assign ces_13_10_io_ins_0 = ces_12_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_10_io_ins_1 = ces_13_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_10_io_ins_2 = ces_14_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_10_io_ins_3 = ces_13_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_11_clock = clock;
  assign ces_13_11_io_ins_0 = ces_12_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_11_io_ins_1 = ces_13_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_11_io_ins_2 = ces_14_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_11_io_ins_3 = ces_13_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_12_clock = clock;
  assign ces_13_12_io_ins_0 = ces_12_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_12_io_ins_1 = ces_13_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_12_io_ins_2 = ces_14_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_12_io_ins_3 = ces_13_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_13_clock = clock;
  assign ces_13_13_io_ins_0 = ces_12_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_13_io_ins_1 = ces_13_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_13_io_ins_2 = ces_14_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_13_io_ins_3 = ces_13_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_14_clock = clock;
  assign ces_13_14_io_ins_0 = ces_12_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_14_io_ins_1 = ces_13_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_13_14_io_ins_2 = ces_14_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_14_io_ins_3 = ces_13_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_13_15_clock = clock;
  assign ces_13_15_io_ins_0 = ces_12_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_13_15_io_ins_1 = io_insVertical_0_13; // @[MockArray.scala 46:87]
  assign ces_13_15_io_ins_2 = ces_14_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_13_15_io_ins_3 = ces_13_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_0_clock = clock;
  assign ces_14_0_io_ins_0 = ces_13_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_0_io_ins_1 = ces_14_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_0_io_ins_2 = ces_15_0_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_0_io_ins_3 = io_insVertical_1_14; // @[MockArray.scala 48:87]
  assign ces_14_1_clock = clock;
  assign ces_14_1_io_ins_0 = ces_13_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_1_io_ins_1 = ces_14_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_1_io_ins_2 = ces_15_1_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_1_io_ins_3 = ces_14_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_2_clock = clock;
  assign ces_14_2_io_ins_0 = ces_13_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_2_io_ins_1 = ces_14_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_2_io_ins_2 = ces_15_2_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_2_io_ins_3 = ces_14_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_3_clock = clock;
  assign ces_14_3_io_ins_0 = ces_13_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_3_io_ins_1 = ces_14_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_3_io_ins_2 = ces_15_3_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_3_io_ins_3 = ces_14_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_4_clock = clock;
  assign ces_14_4_io_ins_0 = ces_13_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_4_io_ins_1 = ces_14_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_4_io_ins_2 = ces_15_4_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_4_io_ins_3 = ces_14_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_5_clock = clock;
  assign ces_14_5_io_ins_0 = ces_13_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_5_io_ins_1 = ces_14_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_5_io_ins_2 = ces_15_5_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_5_io_ins_3 = ces_14_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_6_clock = clock;
  assign ces_14_6_io_ins_0 = ces_13_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_6_io_ins_1 = ces_14_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_6_io_ins_2 = ces_15_6_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_6_io_ins_3 = ces_14_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_7_clock = clock;
  assign ces_14_7_io_ins_0 = ces_13_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_7_io_ins_1 = ces_14_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_7_io_ins_2 = ces_15_7_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_7_io_ins_3 = ces_14_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_8_clock = clock;
  assign ces_14_8_io_ins_0 = ces_13_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_8_io_ins_1 = ces_14_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_8_io_ins_2 = ces_15_8_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_8_io_ins_3 = ces_14_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_9_clock = clock;
  assign ces_14_9_io_ins_0 = ces_13_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_9_io_ins_1 = ces_14_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_9_io_ins_2 = ces_15_9_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_9_io_ins_3 = ces_14_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_10_clock = clock;
  assign ces_14_10_io_ins_0 = ces_13_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_10_io_ins_1 = ces_14_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_10_io_ins_2 = ces_15_10_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_10_io_ins_3 = ces_14_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_11_clock = clock;
  assign ces_14_11_io_ins_0 = ces_13_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_11_io_ins_1 = ces_14_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_11_io_ins_2 = ces_15_11_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_11_io_ins_3 = ces_14_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_12_clock = clock;
  assign ces_14_12_io_ins_0 = ces_13_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_12_io_ins_1 = ces_14_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_12_io_ins_2 = ces_15_12_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_12_io_ins_3 = ces_14_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_13_clock = clock;
  assign ces_14_13_io_ins_0 = ces_13_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_13_io_ins_1 = ces_14_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_13_io_ins_2 = ces_15_13_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_13_io_ins_3 = ces_14_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_14_clock = clock;
  assign ces_14_14_io_ins_0 = ces_13_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_14_io_ins_1 = ces_14_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_14_14_io_ins_2 = ces_15_14_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_14_io_ins_3 = ces_14_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_14_15_clock = clock;
  assign ces_14_15_io_ins_0 = ces_13_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_14_15_io_ins_1 = io_insVertical_0_14; // @[MockArray.scala 46:87]
  assign ces_14_15_io_ins_2 = ces_15_15_io_outs_0; // @[MockArray.scala 57:19]
  assign ces_14_15_io_ins_3 = ces_14_14_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_0_clock = clock;
  assign ces_15_0_io_ins_0 = ces_14_0_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_0_io_ins_1 = ces_15_1_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_0_io_ins_2 = io_insHorizontal_1_0; // @[MockArray.scala 47:87]
  assign ces_15_0_io_ins_3 = io_insVertical_1_15; // @[MockArray.scala 48:87]
  assign ces_15_1_clock = clock;
  assign ces_15_1_io_ins_0 = ces_14_1_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_1_io_ins_1 = ces_15_2_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_1_io_ins_2 = io_insHorizontal_1_1; // @[MockArray.scala 47:87]
  assign ces_15_1_io_ins_3 = ces_15_0_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_2_clock = clock;
  assign ces_15_2_io_ins_0 = ces_14_2_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_2_io_ins_1 = ces_15_3_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_2_io_ins_2 = io_insHorizontal_1_2; // @[MockArray.scala 47:87]
  assign ces_15_2_io_ins_3 = ces_15_1_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_3_clock = clock;
  assign ces_15_3_io_ins_0 = ces_14_3_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_3_io_ins_1 = ces_15_4_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_3_io_ins_2 = io_insHorizontal_1_3; // @[MockArray.scala 47:87]
  assign ces_15_3_io_ins_3 = ces_15_2_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_4_clock = clock;
  assign ces_15_4_io_ins_0 = ces_14_4_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_4_io_ins_1 = ces_15_5_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_4_io_ins_2 = io_insHorizontal_1_4; // @[MockArray.scala 47:87]
  assign ces_15_4_io_ins_3 = ces_15_3_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_5_clock = clock;
  assign ces_15_5_io_ins_0 = ces_14_5_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_5_io_ins_1 = ces_15_6_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_5_io_ins_2 = io_insHorizontal_1_5; // @[MockArray.scala 47:87]
  assign ces_15_5_io_ins_3 = ces_15_4_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_6_clock = clock;
  assign ces_15_6_io_ins_0 = ces_14_6_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_6_io_ins_1 = ces_15_7_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_6_io_ins_2 = io_insHorizontal_1_6; // @[MockArray.scala 47:87]
  assign ces_15_6_io_ins_3 = ces_15_5_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_7_clock = clock;
  assign ces_15_7_io_ins_0 = ces_14_7_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_7_io_ins_1 = ces_15_8_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_7_io_ins_2 = io_insHorizontal_1_7; // @[MockArray.scala 47:87]
  assign ces_15_7_io_ins_3 = ces_15_6_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_8_clock = clock;
  assign ces_15_8_io_ins_0 = ces_14_8_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_8_io_ins_1 = ces_15_9_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_8_io_ins_2 = io_insHorizontal_1_8; // @[MockArray.scala 47:87]
  assign ces_15_8_io_ins_3 = ces_15_7_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_9_clock = clock;
  assign ces_15_9_io_ins_0 = ces_14_9_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_9_io_ins_1 = ces_15_10_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_9_io_ins_2 = io_insHorizontal_1_9; // @[MockArray.scala 47:87]
  assign ces_15_9_io_ins_3 = ces_15_8_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_10_clock = clock;
  assign ces_15_10_io_ins_0 = ces_14_10_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_10_io_ins_1 = ces_15_11_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_10_io_ins_2 = io_insHorizontal_1_10; // @[MockArray.scala 47:87]
  assign ces_15_10_io_ins_3 = ces_15_9_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_11_clock = clock;
  assign ces_15_11_io_ins_0 = ces_14_11_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_11_io_ins_1 = ces_15_12_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_11_io_ins_2 = io_insHorizontal_1_11; // @[MockArray.scala 47:87]
  assign ces_15_11_io_ins_3 = ces_15_10_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_12_clock = clock;
  assign ces_15_12_io_ins_0 = ces_14_12_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_12_io_ins_1 = ces_15_13_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_12_io_ins_2 = io_insHorizontal_1_12; // @[MockArray.scala 47:87]
  assign ces_15_12_io_ins_3 = ces_15_11_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_13_clock = clock;
  assign ces_15_13_io_ins_0 = ces_14_13_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_13_io_ins_1 = ces_15_14_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_13_io_ins_2 = io_insHorizontal_1_13; // @[MockArray.scala 47:87]
  assign ces_15_13_io_ins_3 = ces_15_12_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_14_clock = clock;
  assign ces_15_14_io_ins_0 = ces_14_14_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_14_io_ins_1 = ces_15_15_io_outs_3; // @[MockArray.scala 63:19]
  assign ces_15_14_io_ins_2 = io_insHorizontal_1_14; // @[MockArray.scala 47:87]
  assign ces_15_14_io_ins_3 = ces_15_13_io_outs_1; // @[MockArray.scala 64:19]
  assign ces_15_15_clock = clock;
  assign ces_15_15_io_ins_0 = ces_14_15_io_outs_2; // @[MockArray.scala 58:19]
  assign ces_15_15_io_ins_1 = io_insVertical_0_15; // @[MockArray.scala 46:87]
  assign ces_15_15_io_ins_2 = io_insHorizontal_1_15; // @[MockArray.scala 47:87]
  assign ces_15_15_io_ins_3 = ces_15_14_io_outs_1; // @[MockArray.scala 64:19]
endmodule
