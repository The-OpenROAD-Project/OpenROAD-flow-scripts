module fakeram45_64x64 (
   output reg [63:0] rd_out,
   input logic [5:0] addr_in,
   input logic we_in,
   input logic [63:0] wd_in,
   input logic clk,
   input logic ce_in
);
endmodule
