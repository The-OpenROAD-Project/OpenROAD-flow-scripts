VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO apb_sys_0
  CLASS BLOCK ;
  FOREIGN apb_sys_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 448.090 BY 700.000 ;
  PIN HADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 4.000 ;
    END
  END HADDR[0]
  PIN HADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.720 0.000 44.000 4.000 ;
    END
  END HADDR[10]
  PIN HADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.320 0.000 48.600 4.000 ;
    END
  END HADDR[11]
  PIN HADDR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.920 0.000 53.200 4.000 ;
    END
  END HADDR[12]
  PIN HADDR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.060 0.000 57.340 4.000 ;
    END
  END HADDR[13]
  PIN HADDR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.660 0.000 61.940 4.000 ;
    END
  END HADDR[14]
  PIN HADDR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.800 0.000 66.080 4.000 ;
    END
  END HADDR[15]
  PIN HADDR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.400 0.000 70.680 4.000 ;
    END
  END HADDR[16]
  PIN HADDR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.000 0.000 75.280 4.000 ;
    END
  END HADDR[17]
  PIN HADDR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.140 0.000 79.420 4.000 ;
    END
  END HADDR[18]
  PIN HADDR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.740 0.000 84.020 4.000 ;
    END
  END HADDR[19]
  PIN HADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.160 0.000 4.440 4.000 ;
    END
  END HADDR[1]
  PIN HADDR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.880 0.000 88.160 4.000 ;
    END
  END HADDR[20]
  PIN HADDR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.480 0.000 92.760 4.000 ;
    END
  END HADDR[21]
  PIN HADDR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.620 0.000 96.900 4.000 ;
    END
  END HADDR[22]
  PIN HADDR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.220 0.000 101.500 4.000 ;
    END
  END HADDR[23]
  PIN HADDR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.820 0.000 106.100 4.000 ;
    END
  END HADDR[24]
  PIN HADDR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.960 0.000 110.240 4.000 ;
    END
  END HADDR[25]
  PIN HADDR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.560 0.000 114.840 4.000 ;
    END
  END HADDR[26]
  PIN HADDR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.700 0.000 118.980 4.000 ;
    END
  END HADDR[27]
  PIN HADDR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.300 0.000 123.580 4.000 ;
    END
  END HADDR[28]
  PIN HADDR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.900 0.000 128.180 4.000 ;
    END
  END HADDR[29]
  PIN HADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.760 0.000 9.040 4.000 ;
    END
  END HADDR[2]
  PIN HADDR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.040 0.000 132.320 4.000 ;
    END
  END HADDR[30]
  PIN HADDR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.640 0.000 136.920 4.000 ;
    END
  END HADDR[31]
  PIN HADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.900 0.000 13.180 4.000 ;
    END
  END HADDR[3]
  PIN HADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.500 0.000 17.780 4.000 ;
    END
  END HADDR[4]
  PIN HADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.640 0.000 21.920 4.000 ;
    END
  END HADDR[5]
  PIN HADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.240 0.000 26.520 4.000 ;
    END
  END HADDR[6]
  PIN HADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.840 0.000 31.120 4.000 ;
    END
  END HADDR[7]
  PIN HADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.980 0.000 35.260 4.000 ;
    END
  END HADDR[8]
  PIN HADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.580 0.000 39.860 4.000 ;
    END
  END HADDR[9]
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 19.080 448.090 19.680 ;
    END
  END HCLK
  PIN HRDATA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.780 0.000 141.060 4.000 ;
    END
  END HRDATA[0]
  PIN HRDATA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.940 0.000 185.220 4.000 ;
    END
  END HRDATA[10]
  PIN HRDATA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.540 0.000 189.820 4.000 ;
    END
  END HRDATA[11]
  PIN HRDATA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.680 0.000 193.960 4.000 ;
    END
  END HRDATA[12]
  PIN HRDATA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.280 0.000 198.560 4.000 ;
    END
  END HRDATA[13]
  PIN HRDATA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.880 0.000 203.160 4.000 ;
    END
  END HRDATA[14]
  PIN HRDATA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.020 0.000 207.300 4.000 ;
    END
  END HRDATA[15]
  PIN HRDATA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.620 0.000 211.900 4.000 ;
    END
  END HRDATA[16]
  PIN HRDATA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.760 0.000 216.040 4.000 ;
    END
  END HRDATA[17]
  PIN HRDATA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.360 0.000 220.640 4.000 ;
    END
  END HRDATA[18]
  PIN HRDATA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.960 0.000 225.240 4.000 ;
    END
  END HRDATA[19]
  PIN HRDATA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.380 0.000 145.660 4.000 ;
    END
  END HRDATA[1]
  PIN HRDATA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.100 0.000 229.380 4.000 ;
    END
  END HRDATA[20]
  PIN HRDATA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.700 0.000 233.980 4.000 ;
    END
  END HRDATA[21]
  PIN HRDATA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.840 0.000 238.120 4.000 ;
    END
  END HRDATA[22]
  PIN HRDATA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.440 0.000 242.720 4.000 ;
    END
  END HRDATA[23]
  PIN HRDATA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.580 0.000 246.860 4.000 ;
    END
  END HRDATA[24]
  PIN HRDATA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.180 0.000 251.460 4.000 ;
    END
  END HRDATA[25]
  PIN HRDATA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.780 0.000 256.060 4.000 ;
    END
  END HRDATA[26]
  PIN HRDATA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.920 0.000 260.200 4.000 ;
    END
  END HRDATA[27]
  PIN HRDATA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.520 0.000 264.800 4.000 ;
    END
  END HRDATA[28]
  PIN HRDATA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.660 0.000 268.940 4.000 ;
    END
  END HRDATA[29]
  PIN HRDATA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.980 0.000 150.260 4.000 ;
    END
  END HRDATA[2]
  PIN HRDATA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.260 0.000 273.540 4.000 ;
    END
  END HRDATA[30]
  PIN HRDATA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.860 0.000 278.140 4.000 ;
    END
  END HRDATA[31]
  PIN HRDATA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.120 0.000 154.400 4.000 ;
    END
  END HRDATA[3]
  PIN HRDATA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.720 0.000 159.000 4.000 ;
    END
  END HRDATA[4]
  PIN HRDATA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.860 0.000 163.140 4.000 ;
    END
  END HRDATA[5]
  PIN HRDATA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.460 0.000 167.740 4.000 ;
    END
  END HRDATA[6]
  PIN HRDATA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.600 0.000 171.880 4.000 ;
    END
  END HRDATA[7]
  PIN HRDATA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.200 0.000 176.480 4.000 ;
    END
  END HRDATA[8]
  PIN HRDATA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.800 0.000 181.080 4.000 ;
    END
  END HRDATA[9]
  PIN HREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.560 0.000 436.840 4.000 ;
    END
  END HREADY
  PIN HREADYOUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.300 0.000 445.580 4.000 ;
    END
  END HREADYOUT
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 57.840 448.090 58.440 ;
    END
  END HRESETn
  PIN HSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.700 0.000 440.980 4.000 ;
    END
  END HSEL
  PIN HTRANS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.220 0.000 423.500 4.000 ;
    END
  END HTRANS[0]
  PIN HTRANS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.820 0.000 428.100 4.000 ;
    END
  END HTRANS[1]
  PIN HWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.000 0.000 282.280 4.000 ;
    END
  END HWDATA[0]
  PIN HWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.160 0.000 326.440 4.000 ;
    END
  END HWDATA[10]
  PIN HWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.760 0.000 331.040 4.000 ;
    END
  END HWDATA[11]
  PIN HWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.900 0.000 335.180 4.000 ;
    END
  END HWDATA[12]
  PIN HWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.500 0.000 339.780 4.000 ;
    END
  END HWDATA[13]
  PIN HWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.640 0.000 343.920 4.000 ;
    END
  END HWDATA[14]
  PIN HWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.240 0.000 348.520 4.000 ;
    END
  END HWDATA[15]
  PIN HWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.840 0.000 353.120 4.000 ;
    END
  END HWDATA[16]
  PIN HWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.980 0.000 357.260 4.000 ;
    END
  END HWDATA[17]
  PIN HWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.580 0.000 361.860 4.000 ;
    END
  END HWDATA[18]
  PIN HWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.720 0.000 366.000 4.000 ;
    END
  END HWDATA[19]
  PIN HWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.600 0.000 286.880 4.000 ;
    END
  END HWDATA[1]
  PIN HWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.320 0.000 370.600 4.000 ;
    END
  END HWDATA[20]
  PIN HWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.920 0.000 375.200 4.000 ;
    END
  END HWDATA[21]
  PIN HWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.060 0.000 379.340 4.000 ;
    END
  END HWDATA[22]
  PIN HWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.660 0.000 383.940 4.000 ;
    END
  END HWDATA[23]
  PIN HWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.800 0.000 388.080 4.000 ;
    END
  END HWDATA[24]
  PIN HWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.400 0.000 392.680 4.000 ;
    END
  END HWDATA[25]
  PIN HWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.540 0.000 396.820 4.000 ;
    END
  END HWDATA[26]
  PIN HWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.140 0.000 401.420 4.000 ;
    END
  END HWDATA[27]
  PIN HWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.740 0.000 406.020 4.000 ;
    END
  END HWDATA[28]
  PIN HWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.880 0.000 410.160 4.000 ;
    END
  END HWDATA[29]
  PIN HWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.740 0.000 291.020 4.000 ;
    END
  END HWDATA[2]
  PIN HWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.480 0.000 414.760 4.000 ;
    END
  END HWDATA[30]
  PIN HWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.620 0.000 418.900 4.000 ;
    END
  END HWDATA[31]
  PIN HWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.340 0.000 295.620 4.000 ;
    END
  END HWDATA[3]
  PIN HWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.940 0.000 300.220 4.000 ;
    END
  END HWDATA[4]
  PIN HWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.080 0.000 304.360 4.000 ;
    END
  END HWDATA[5]
  PIN HWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.680 0.000 308.960 4.000 ;
    END
  END HWDATA[6]
  PIN HWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.820 0.000 313.100 4.000 ;
    END
  END HWDATA[7]
  PIN HWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.420 0.000 317.700 4.000 ;
    END
  END HWDATA[8]
  PIN HWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.560 0.000 321.840 4.000 ;
    END
  END HWDATA[9]
  PIN HWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.960 0.000 432.240 4.000 ;
    END
  END HWRITE
  PIN IRQ[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 96.600 448.090 97.200 ;
    END
  END IRQ[0]
  PIN IRQ[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 485.560 448.090 486.160 ;
    END
  END IRQ[10]
  PIN IRQ[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 524.320 448.090 524.920 ;
    END
  END IRQ[11]
  PIN IRQ[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 563.080 448.090 563.680 ;
    END
  END IRQ[12]
  PIN IRQ[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 601.840 448.090 602.440 ;
    END
  END IRQ[13]
  PIN IRQ[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 640.600 448.090 641.200 ;
    END
  END IRQ[14]
  PIN IRQ[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 679.360 448.090 679.960 ;
    END
  END IRQ[15]
  PIN IRQ[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 135.360 448.090 135.960 ;
    END
  END IRQ[1]
  PIN IRQ[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 174.120 448.090 174.720 ;
    END
  END IRQ[2]
  PIN IRQ[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 212.880 448.090 213.480 ;
    END
  END IRQ[3]
  PIN IRQ[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 252.320 448.090 252.920 ;
    END
  END IRQ[4]
  PIN IRQ[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 291.080 448.090 291.680 ;
    END
  END IRQ[5]
  PIN IRQ[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 329.840 448.090 330.440 ;
    END
  END IRQ[6]
  PIN IRQ[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 368.600 448.090 369.200 ;
    END
  END IRQ[7]
  PIN IRQ[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 407.360 448.090 407.960 ;
    END
  END IRQ[8]
  PIN IRQ[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 444.090 446.120 448.090 446.720 ;
    END
  END IRQ[9]
  PIN MSI_S2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.460 696.000 75.740 700.000 ;
    END
  END MSI_S2
  PIN MSI_S3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.460 696.000 144.740 700.000 ;
    END
  END MSI_S3
  PIN MSO_S2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.940 696.000 93.220 700.000 ;
    END
  END MSO_S2
  PIN MSO_S3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.940 696.000 162.220 700.000 ;
    END
  END MSO_S3
  PIN RsRx_S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.460 696.000 6.740 700.000 ;
    END
  END RsRx_S0
  PIN RsRx_S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.960 696.000 41.240 700.000 ;
    END
  END RsRx_S1
  PIN RsTx_S0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.480 696.000 23.760 700.000 ;
    END
  END RsTx_S0
  PIN RsTx_S1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.980 696.000 58.260 700.000 ;
    END
  END RsTx_S1
  PIN SCLK_S2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.440 696.000 127.720 700.000 ;
    END
  END SCLK_S2
  PIN SCLK_S3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.440 696.000 196.720 700.000 ;
    END
  END SCLK_S3
  PIN SSn_S2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.960 696.000 110.240 700.000 ;
    END
  END SSn_S2
  PIN SSn_S3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.420 696.000 179.700 700.000 ;
    END
  END SSn_S3
  PIN pwm_S6
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.380 696.000 421.660 700.000 ;
    END
  END pwm_S6
  PIN pwm_S7
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.860 696.000 439.140 700.000 ;
    END
  END pwm_S7
  PIN scl_i_S4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.920 696.000 214.200 700.000 ;
    END
  END scl_i_S4
  PIN scl_i_S5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.880 696.000 318.160 700.000 ;
    END
  END scl_i_S5
  PIN scl_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.400 696.000 231.680 700.000 ;
    END
  END scl_o_S4
  PIN scl_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.900 696.000 335.180 700.000 ;
    END
  END scl_o_S5
  PIN scl_oen_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.420 696.000 248.700 700.000 ;
    END
  END scl_oen_o_S4
  PIN scl_oen_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.380 696.000 352.660 700.000 ;
    END
  END scl_oen_o_S5
  PIN sda_i_S4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.900 696.000 266.180 700.000 ;
    END
  END sda_i_S4
  PIN sda_i_S5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.400 696.000 369.680 700.000 ;
    END
  END sda_i_S5
  PIN sda_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.920 696.000 283.200 700.000 ;
    END
  END sda_o_S4
  PIN sda_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.880 696.000 387.160 700.000 ;
    END
  END sda_o_S5
  PIN sda_oen_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.400 696.000 300.680 700.000 ;
    END
  END sda_oen_o_S4
  PIN sda_oen_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.360 696.000 404.640 700.000 ;
    END
  END sda_oen_o_S5
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 326.330 10.640 327.930 688.400 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 172.730 10.640 174.330 688.400 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.130 10.640 20.730 688.400 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 403.130 10.640 404.730 688.400 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 249.530 10.640 251.130 688.400 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.930 10.640 97.530 688.400 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 3.610 10.795 443.685 688.245 ;
      LAYER met1 ;
        RECT 0.000 9.220 446.060 688.400 ;
      LAYER met2 ;
        RECT 0.030 695.720 6.180 696.050 ;
        RECT 7.020 695.720 23.200 696.050 ;
        RECT 24.040 695.720 40.680 696.050 ;
        RECT 41.520 695.720 57.700 696.050 ;
        RECT 58.540 695.720 75.180 696.050 ;
        RECT 76.020 695.720 92.660 696.050 ;
        RECT 93.500 695.720 109.680 696.050 ;
        RECT 110.520 695.720 127.160 696.050 ;
        RECT 128.000 695.720 144.180 696.050 ;
        RECT 145.020 695.720 161.660 696.050 ;
        RECT 162.500 695.720 179.140 696.050 ;
        RECT 179.980 695.720 196.160 696.050 ;
        RECT 197.000 695.720 213.640 696.050 ;
        RECT 214.480 695.720 231.120 696.050 ;
        RECT 231.960 695.720 248.140 696.050 ;
        RECT 248.980 695.720 265.620 696.050 ;
        RECT 266.460 695.720 282.640 696.050 ;
        RECT 283.480 695.720 300.120 696.050 ;
        RECT 300.960 695.720 317.600 696.050 ;
        RECT 318.440 695.720 334.620 696.050 ;
        RECT 335.460 695.720 352.100 696.050 ;
        RECT 352.940 695.720 369.120 696.050 ;
        RECT 369.960 695.720 386.600 696.050 ;
        RECT 387.440 695.720 404.080 696.050 ;
        RECT 404.920 695.720 421.100 696.050 ;
        RECT 421.940 695.720 438.580 696.050 ;
        RECT 439.420 695.720 446.040 696.050 ;
        RECT 0.030 4.280 446.040 695.720 ;
        RECT 0.580 4.000 3.880 4.280 ;
        RECT 4.720 4.000 8.480 4.280 ;
        RECT 9.320 4.000 12.620 4.280 ;
        RECT 13.460 4.000 17.220 4.280 ;
        RECT 18.060 4.000 21.360 4.280 ;
        RECT 22.200 4.000 25.960 4.280 ;
        RECT 26.800 4.000 30.560 4.280 ;
        RECT 31.400 4.000 34.700 4.280 ;
        RECT 35.540 4.000 39.300 4.280 ;
        RECT 40.140 4.000 43.440 4.280 ;
        RECT 44.280 4.000 48.040 4.280 ;
        RECT 48.880 4.000 52.640 4.280 ;
        RECT 53.480 4.000 56.780 4.280 ;
        RECT 57.620 4.000 61.380 4.280 ;
        RECT 62.220 4.000 65.520 4.280 ;
        RECT 66.360 4.000 70.120 4.280 ;
        RECT 70.960 4.000 74.720 4.280 ;
        RECT 75.560 4.000 78.860 4.280 ;
        RECT 79.700 4.000 83.460 4.280 ;
        RECT 84.300 4.000 87.600 4.280 ;
        RECT 88.440 4.000 92.200 4.280 ;
        RECT 93.040 4.000 96.340 4.280 ;
        RECT 97.180 4.000 100.940 4.280 ;
        RECT 101.780 4.000 105.540 4.280 ;
        RECT 106.380 4.000 109.680 4.280 ;
        RECT 110.520 4.000 114.280 4.280 ;
        RECT 115.120 4.000 118.420 4.280 ;
        RECT 119.260 4.000 123.020 4.280 ;
        RECT 123.860 4.000 127.620 4.280 ;
        RECT 128.460 4.000 131.760 4.280 ;
        RECT 132.600 4.000 136.360 4.280 ;
        RECT 137.200 4.000 140.500 4.280 ;
        RECT 141.340 4.000 145.100 4.280 ;
        RECT 145.940 4.000 149.700 4.280 ;
        RECT 150.540 4.000 153.840 4.280 ;
        RECT 154.680 4.000 158.440 4.280 ;
        RECT 159.280 4.000 162.580 4.280 ;
        RECT 163.420 4.000 167.180 4.280 ;
        RECT 168.020 4.000 171.320 4.280 ;
        RECT 172.160 4.000 175.920 4.280 ;
        RECT 176.760 4.000 180.520 4.280 ;
        RECT 181.360 4.000 184.660 4.280 ;
        RECT 185.500 4.000 189.260 4.280 ;
        RECT 190.100 4.000 193.400 4.280 ;
        RECT 194.240 4.000 198.000 4.280 ;
        RECT 198.840 4.000 202.600 4.280 ;
        RECT 203.440 4.000 206.740 4.280 ;
        RECT 207.580 4.000 211.340 4.280 ;
        RECT 212.180 4.000 215.480 4.280 ;
        RECT 216.320 4.000 220.080 4.280 ;
        RECT 220.920 4.000 224.680 4.280 ;
        RECT 225.520 4.000 228.820 4.280 ;
        RECT 229.660 4.000 233.420 4.280 ;
        RECT 234.260 4.000 237.560 4.280 ;
        RECT 238.400 4.000 242.160 4.280 ;
        RECT 243.000 4.000 246.300 4.280 ;
        RECT 247.140 4.000 250.900 4.280 ;
        RECT 251.740 4.000 255.500 4.280 ;
        RECT 256.340 4.000 259.640 4.280 ;
        RECT 260.480 4.000 264.240 4.280 ;
        RECT 265.080 4.000 268.380 4.280 ;
        RECT 269.220 4.000 272.980 4.280 ;
        RECT 273.820 4.000 277.580 4.280 ;
        RECT 278.420 4.000 281.720 4.280 ;
        RECT 282.560 4.000 286.320 4.280 ;
        RECT 287.160 4.000 290.460 4.280 ;
        RECT 291.300 4.000 295.060 4.280 ;
        RECT 295.900 4.000 299.660 4.280 ;
        RECT 300.500 4.000 303.800 4.280 ;
        RECT 304.640 4.000 308.400 4.280 ;
        RECT 309.240 4.000 312.540 4.280 ;
        RECT 313.380 4.000 317.140 4.280 ;
        RECT 317.980 4.000 321.280 4.280 ;
        RECT 322.120 4.000 325.880 4.280 ;
        RECT 326.720 4.000 330.480 4.280 ;
        RECT 331.320 4.000 334.620 4.280 ;
        RECT 335.460 4.000 339.220 4.280 ;
        RECT 340.060 4.000 343.360 4.280 ;
        RECT 344.200 4.000 347.960 4.280 ;
        RECT 348.800 4.000 352.560 4.280 ;
        RECT 353.400 4.000 356.700 4.280 ;
        RECT 357.540 4.000 361.300 4.280 ;
        RECT 362.140 4.000 365.440 4.280 ;
        RECT 366.280 4.000 370.040 4.280 ;
        RECT 370.880 4.000 374.640 4.280 ;
        RECT 375.480 4.000 378.780 4.280 ;
        RECT 379.620 4.000 383.380 4.280 ;
        RECT 384.220 4.000 387.520 4.280 ;
        RECT 388.360 4.000 392.120 4.280 ;
        RECT 392.960 4.000 396.260 4.280 ;
        RECT 397.100 4.000 400.860 4.280 ;
        RECT 401.700 4.000 405.460 4.280 ;
        RECT 406.300 4.000 409.600 4.280 ;
        RECT 410.440 4.000 414.200 4.280 ;
        RECT 415.040 4.000 418.340 4.280 ;
        RECT 419.180 4.000 422.940 4.280 ;
        RECT 423.780 4.000 427.540 4.280 ;
        RECT 428.380 4.000 431.680 4.280 ;
        RECT 432.520 4.000 436.280 4.280 ;
        RECT 437.120 4.000 440.420 4.280 ;
        RECT 441.260 4.000 445.020 4.280 ;
        RECT 445.860 4.000 446.040 4.280 ;
      LAYER met3 ;
        RECT 4.135 680.360 446.065 688.325 ;
        RECT 4.135 678.960 443.690 680.360 ;
        RECT 4.135 641.600 446.065 678.960 ;
        RECT 4.135 640.200 443.690 641.600 ;
        RECT 4.135 602.840 446.065 640.200 ;
        RECT 4.135 601.440 443.690 602.840 ;
        RECT 4.135 564.080 446.065 601.440 ;
        RECT 4.135 562.680 443.690 564.080 ;
        RECT 4.135 525.320 446.065 562.680 ;
        RECT 4.135 523.920 443.690 525.320 ;
        RECT 4.135 486.560 446.065 523.920 ;
        RECT 4.135 485.160 443.690 486.560 ;
        RECT 4.135 447.120 446.065 485.160 ;
        RECT 4.135 445.720 443.690 447.120 ;
        RECT 4.135 408.360 446.065 445.720 ;
        RECT 4.135 406.960 443.690 408.360 ;
        RECT 4.135 369.600 446.065 406.960 ;
        RECT 4.135 368.200 443.690 369.600 ;
        RECT 4.135 330.840 446.065 368.200 ;
        RECT 4.135 329.440 443.690 330.840 ;
        RECT 4.135 292.080 446.065 329.440 ;
        RECT 4.135 290.680 443.690 292.080 ;
        RECT 4.135 253.320 446.065 290.680 ;
        RECT 4.135 251.920 443.690 253.320 ;
        RECT 4.135 213.880 446.065 251.920 ;
        RECT 4.135 212.480 443.690 213.880 ;
        RECT 4.135 175.120 446.065 212.480 ;
        RECT 4.135 173.720 443.690 175.120 ;
        RECT 4.135 136.360 446.065 173.720 ;
        RECT 4.135 134.960 443.690 136.360 ;
        RECT 4.135 97.600 446.065 134.960 ;
        RECT 4.135 96.200 443.690 97.600 ;
        RECT 4.135 58.840 446.065 96.200 ;
        RECT 4.135 57.440 443.690 58.840 ;
        RECT 4.135 20.080 446.065 57.440 ;
        RECT 4.135 18.680 443.690 20.080 ;
        RECT 4.135 10.715 446.065 18.680 ;
      LAYER met4 ;
        RECT 21.385 12.415 95.530 680.505 ;
        RECT 97.930 12.415 172.330 680.505 ;
        RECT 174.730 12.415 249.130 680.505 ;
        RECT 251.530 12.415 325.930 680.505 ;
        RECT 328.330 12.415 402.730 680.505 ;
        RECT 405.130 12.415 438.475 680.505 ;
  END
END apb_sys_0
END LIBRARY

