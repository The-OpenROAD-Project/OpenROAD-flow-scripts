module MuxTest_width_256_inputs_4_outputs_8_pipeline_5( // @[:@3.2]
  input          clock, // @[:@4.4]
  input          reset, // @[:@5.4]
  input  [1:0]   io_selects_0_0, // @[:@6.4]
  input  [1:0]   io_selects_0_1, // @[:@6.4]
  input  [1:0]   io_selects_1_0, // @[:@6.4]
  input  [1:0]   io_selects_1_1, // @[:@6.4]
  input  [1:0]   io_selects_2_0, // @[:@6.4]
  input  [1:0]   io_selects_2_1, // @[:@6.4]
  input  [1:0]   io_selects_3_0, // @[:@6.4]
  input  [1:0]   io_selects_3_1, // @[:@6.4]
  input  [1:0]   io_selects_4_0, // @[:@6.4]
  input  [1:0]   io_selects_4_1, // @[:@6.4]
  input  [1:0]   io_selects_5_0, // @[:@6.4]
  input  [1:0]   io_selects_5_1, // @[:@6.4]
  input  [1:0]   io_selects_6_0, // @[:@6.4]
  input  [1:0]   io_selects_6_1, // @[:@6.4]
  input  [1:0]   io_selects_7_0, // @[:@6.4]
  input  [1:0]   io_selects_7_1, // @[:@6.4]
  input  [2:0]   io_operation_0, // @[:@6.4]
  input  [2:0]   io_operation_1, // @[:@6.4]
  input  [2:0]   io_operation_2, // @[:@6.4]
  input  [2:0]   io_operation_3, // @[:@6.4]
  input  [2:0]   io_operation_4, // @[:@6.4]
  input  [2:0]   io_operation_5, // @[:@6.4]
  input  [2:0]   io_operation_6, // @[:@6.4]
  input  [2:0]   io_operation_7, // @[:@6.4]
  input  [255:0] io_inputs_0, // @[:@6.4]
  input  [255:0] io_inputs_1, // @[:@6.4]
  input  [255:0] io_inputs_2, // @[:@6.4]
  input  [255:0] io_inputs_3, // @[:@6.4]
  output [255:0] io_outputs_0, // @[:@6.4]
  output [255:0] io_outputs_1, // @[:@6.4]
  output [255:0] io_outputs_2, // @[:@6.4]
  output [255:0] io_outputs_3, // @[:@6.4]
  output [255:0] io_outputs_4, // @[:@6.4]
  output [255:0] io_outputs_5, // @[:@6.4]
  output [255:0] io_outputs_6, // @[:@6.4]
  output [255:0] io_outputs_7 // @[:@6.4]
);
  wire [255:0] _GEN_1; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _GEN_2; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _GEN_3; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _GEN_5; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _GEN_6; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _GEN_7; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [256:0] _T_394; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  wire [255:0] _T_395; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@9.4]
  wire [511:0] _T_397; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@10.4]
  wire [255:0] _T_399; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@11.4]
  wire  _T_400; // @[Mux.scala 46:19:@12.4]
  wire [255:0] _T_401; // @[Mux.scala 46:16:@13.4]
  wire  _T_402; // @[Mux.scala 46:19:@14.4]
  wire [511:0] _T_403; // @[Mux.scala 46:16:@15.4]
  wire  _T_404; // @[Mux.scala 46:19:@16.4]
  wire [511:0] _T_405; // @[Mux.scala 46:16:@17.4]
  wire  _T_406; // @[Mux.scala 46:19:@18.4]
  wire [255:0] _GEN_9; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _GEN_10; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _GEN_11; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _GEN_13; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _GEN_14; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _GEN_15; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [256:0] _T_411; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  wire [255:0] _T_412; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@21.4]
  wire [511:0] _T_414; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@22.4]
  wire [255:0] _T_416; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@23.4]
  wire  _T_417; // @[Mux.scala 46:19:@24.4]
  wire [255:0] _T_418; // @[Mux.scala 46:16:@25.4]
  wire  _T_419; // @[Mux.scala 46:19:@26.4]
  wire [511:0] _T_420; // @[Mux.scala 46:16:@27.4]
  wire  _T_421; // @[Mux.scala 46:19:@28.4]
  wire [511:0] _T_422; // @[Mux.scala 46:16:@29.4]
  wire  _T_423; // @[Mux.scala 46:19:@30.4]
  wire [255:0] _GEN_17; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _GEN_18; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _GEN_19; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _GEN_21; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _GEN_22; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _GEN_23; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [256:0] _T_428; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  wire [255:0] _T_429; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@33.4]
  wire [511:0] _T_431; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@34.4]
  wire [255:0] _T_433; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@35.4]
  wire  _T_434; // @[Mux.scala 46:19:@36.4]
  wire [255:0] _T_435; // @[Mux.scala 46:16:@37.4]
  wire  _T_436; // @[Mux.scala 46:19:@38.4]
  wire [511:0] _T_437; // @[Mux.scala 46:16:@39.4]
  wire  _T_438; // @[Mux.scala 46:19:@40.4]
  wire [511:0] _T_439; // @[Mux.scala 46:16:@41.4]
  wire  _T_440; // @[Mux.scala 46:19:@42.4]
  wire [255:0] _GEN_25; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _GEN_26; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _GEN_27; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _GEN_29; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _GEN_30; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _GEN_31; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [256:0] _T_445; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  wire [255:0] _T_446; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@45.4]
  wire [511:0] _T_448; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@46.4]
  wire [255:0] _T_450; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@47.4]
  wire  _T_451; // @[Mux.scala 46:19:@48.4]
  wire [255:0] _T_452; // @[Mux.scala 46:16:@49.4]
  wire  _T_453; // @[Mux.scala 46:19:@50.4]
  wire [511:0] _T_454; // @[Mux.scala 46:16:@51.4]
  wire  _T_455; // @[Mux.scala 46:19:@52.4]
  wire [511:0] _T_456; // @[Mux.scala 46:16:@53.4]
  wire  _T_457; // @[Mux.scala 46:19:@54.4]
  wire [255:0] _GEN_33; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _GEN_34; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _GEN_35; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _GEN_37; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _GEN_38; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _GEN_39; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [256:0] _T_462; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  wire [255:0] _T_463; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@57.4]
  wire [511:0] _T_465; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@58.4]
  wire [255:0] _T_467; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@59.4]
  wire  _T_468; // @[Mux.scala 46:19:@60.4]
  wire [255:0] _T_469; // @[Mux.scala 46:16:@61.4]
  wire  _T_470; // @[Mux.scala 46:19:@62.4]
  wire [511:0] _T_471; // @[Mux.scala 46:16:@63.4]
  wire  _T_472; // @[Mux.scala 46:19:@64.4]
  wire [511:0] _T_473; // @[Mux.scala 46:16:@65.4]
  wire  _T_474; // @[Mux.scala 46:19:@66.4]
  wire [255:0] _GEN_41; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _GEN_42; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _GEN_43; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _GEN_45; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _GEN_46; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _GEN_47; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [256:0] _T_479; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  wire [255:0] _T_480; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@69.4]
  wire [511:0] _T_482; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@70.4]
  wire [255:0] _T_484; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@71.4]
  wire  _T_485; // @[Mux.scala 46:19:@72.4]
  wire [255:0] _T_486; // @[Mux.scala 46:16:@73.4]
  wire  _T_487; // @[Mux.scala 46:19:@74.4]
  wire [511:0] _T_488; // @[Mux.scala 46:16:@75.4]
  wire  _T_489; // @[Mux.scala 46:19:@76.4]
  wire [511:0] _T_490; // @[Mux.scala 46:16:@77.4]
  wire  _T_491; // @[Mux.scala 46:19:@78.4]
  wire [255:0] _GEN_49; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _GEN_50; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _GEN_51; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _GEN_53; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _GEN_54; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _GEN_55; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [256:0] _T_496; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  wire [255:0] _T_497; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@81.4]
  wire [511:0] _T_499; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@82.4]
  wire [255:0] _T_501; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@83.4]
  wire  _T_502; // @[Mux.scala 46:19:@84.4]
  wire [255:0] _T_503; // @[Mux.scala 46:16:@85.4]
  wire  _T_504; // @[Mux.scala 46:19:@86.4]
  wire [511:0] _T_505; // @[Mux.scala 46:16:@87.4]
  wire  _T_506; // @[Mux.scala 46:19:@88.4]
  wire [511:0] _T_507; // @[Mux.scala 46:16:@89.4]
  wire  _T_508; // @[Mux.scala 46:19:@90.4]
  wire [255:0] _GEN_57; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _GEN_58; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _GEN_59; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _GEN_61; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _GEN_62; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _GEN_63; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [256:0] _T_513; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  wire [255:0] _T_514; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@93.4]
  wire [511:0] _T_516; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@94.4]
  wire [255:0] _T_518; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@95.4]
  wire  _T_519; // @[Mux.scala 46:19:@96.4]
  wire [255:0] _T_520; // @[Mux.scala 46:16:@97.4]
  wire  _T_521; // @[Mux.scala 46:19:@98.4]
  wire [511:0] _T_522; // @[Mux.scala 46:16:@99.4]
  wire  _T_523; // @[Mux.scala 46:19:@100.4]
  wire [511:0] _T_524; // @[Mux.scala 46:16:@101.4]
  wire  _T_525; // @[Mux.scala 46:19:@102.4]
  reg [511:0] _T_529; // @[Reg.scala 11:16:@104.4]
  reg [511:0] _RAND_0;
  reg [511:0] _T_531; // @[Reg.scala 11:16:@108.4]
  reg [511:0] _RAND_1;
  reg [511:0] _T_533; // @[Reg.scala 11:16:@112.4]
  reg [511:0] _RAND_2;
  reg [511:0] _T_535; // @[Reg.scala 11:16:@116.4]
  reg [511:0] _RAND_3;
  reg [511:0] _T_537; // @[Reg.scala 11:16:@120.4]
  reg [511:0] _RAND_4;
  reg [511:0] _T_540; // @[Reg.scala 11:16:@124.4]
  reg [511:0] _RAND_5;
  reg [511:0] _T_542; // @[Reg.scala 11:16:@128.4]
  reg [511:0] _RAND_6;
  reg [511:0] _T_544; // @[Reg.scala 11:16:@132.4]
  reg [511:0] _RAND_7;
  reg [511:0] _T_546; // @[Reg.scala 11:16:@136.4]
  reg [511:0] _RAND_8;
  reg [511:0] _T_548; // @[Reg.scala 11:16:@140.4]
  reg [511:0] _RAND_9;
  reg [511:0] _T_551; // @[Reg.scala 11:16:@144.4]
  reg [511:0] _RAND_10;
  reg [511:0] _T_553; // @[Reg.scala 11:16:@148.4]
  reg [511:0] _RAND_11;
  reg [511:0] _T_555; // @[Reg.scala 11:16:@152.4]
  reg [511:0] _RAND_12;
  reg [511:0] _T_557; // @[Reg.scala 11:16:@156.4]
  reg [511:0] _RAND_13;
  reg [511:0] _T_559; // @[Reg.scala 11:16:@160.4]
  reg [511:0] _RAND_14;
  reg [511:0] _T_562; // @[Reg.scala 11:16:@164.4]
  reg [511:0] _RAND_15;
  reg [511:0] _T_564; // @[Reg.scala 11:16:@168.4]
  reg [511:0] _RAND_16;
  reg [511:0] _T_566; // @[Reg.scala 11:16:@172.4]
  reg [511:0] _RAND_17;
  reg [511:0] _T_568; // @[Reg.scala 11:16:@176.4]
  reg [511:0] _RAND_18;
  reg [511:0] _T_570; // @[Reg.scala 11:16:@180.4]
  reg [511:0] _RAND_19;
  reg [511:0] _T_573; // @[Reg.scala 11:16:@184.4]
  reg [511:0] _RAND_20;
  reg [511:0] _T_575; // @[Reg.scala 11:16:@188.4]
  reg [511:0] _RAND_21;
  reg [511:0] _T_577; // @[Reg.scala 11:16:@192.4]
  reg [511:0] _RAND_22;
  reg [511:0] _T_579; // @[Reg.scala 11:16:@196.4]
  reg [511:0] _RAND_23;
  reg [511:0] _T_581; // @[Reg.scala 11:16:@200.4]
  reg [511:0] _RAND_24;
  reg [511:0] _T_584; // @[Reg.scala 11:16:@204.4]
  reg [511:0] _RAND_25;
  reg [511:0] _T_586; // @[Reg.scala 11:16:@208.4]
  reg [511:0] _RAND_26;
  reg [511:0] _T_588; // @[Reg.scala 11:16:@212.4]
  reg [511:0] _RAND_27;
  reg [511:0] _T_590; // @[Reg.scala 11:16:@216.4]
  reg [511:0] _RAND_28;
  reg [511:0] _T_592; // @[Reg.scala 11:16:@220.4]
  reg [511:0] _RAND_29;
  reg [511:0] _T_595; // @[Reg.scala 11:16:@224.4]
  reg [511:0] _RAND_30;
  reg [511:0] _T_597; // @[Reg.scala 11:16:@228.4]
  reg [511:0] _RAND_31;
  reg [511:0] _T_599; // @[Reg.scala 11:16:@232.4]
  reg [511:0] _RAND_32;
  reg [511:0] _T_601; // @[Reg.scala 11:16:@236.4]
  reg [511:0] _RAND_33;
  reg [511:0] _T_603; // @[Reg.scala 11:16:@240.4]
  reg [511:0] _RAND_34;
  reg [511:0] _T_606; // @[Reg.scala 11:16:@244.4]
  reg [511:0] _RAND_35;
  reg [511:0] _T_608; // @[Reg.scala 11:16:@248.4]
  reg [511:0] _RAND_36;
  reg [511:0] _T_610; // @[Reg.scala 11:16:@252.4]
  reg [511:0] _RAND_37;
  reg [511:0] _T_612; // @[Reg.scala 11:16:@256.4]
  reg [511:0] _RAND_38;
  reg [511:0] _T_614; // @[Reg.scala 11:16:@260.4]
  reg [511:0] _RAND_39;
  assign _GEN_1 = 2'h1 == io_selects_0_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_2 = 2'h2 == io_selects_0_0 ? io_inputs_2 : _GEN_1; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_3 = 2'h3 == io_selects_0_0 ? io_inputs_3 : _GEN_2; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_5 = 2'h1 == io_selects_0_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_6 = 2'h2 == io_selects_0_1 ? io_inputs_2 : _GEN_5; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _GEN_7 = 2'h3 == io_selects_0_1 ? io_inputs_3 : _GEN_6; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _T_394 = _GEN_3 + _GEN_7; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@8.4]
  assign _T_395 = _GEN_3 + _GEN_7; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@9.4]
  assign _T_397 = _GEN_3 * _GEN_7; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@10.4]
  assign _T_399 = _GEN_3 / _GEN_7; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@11.4]
  assign _T_400 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_401 = _T_400 ? _T_399 : 256'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_402 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_403 = _T_402 ? _T_397 : {{256'd0}, _T_401}; // @[Mux.scala 46:16:@15.4]
  assign _T_404 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_405 = _T_404 ? {{256'd0}, _T_395} : _T_403; // @[Mux.scala 46:16:@17.4]
  assign _T_406 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _GEN_9 = 2'h1 == io_selects_1_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_10 = 2'h2 == io_selects_1_0 ? io_inputs_2 : _GEN_9; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_11 = 2'h3 == io_selects_1_0 ? io_inputs_3 : _GEN_10; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_13 = 2'h1 == io_selects_1_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_14 = 2'h2 == io_selects_1_1 ? io_inputs_2 : _GEN_13; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _GEN_15 = 2'h3 == io_selects_1_1 ? io_inputs_3 : _GEN_14; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _T_411 = _GEN_11 + _GEN_15; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@20.4]
  assign _T_412 = _GEN_11 + _GEN_15; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@21.4]
  assign _T_414 = _GEN_11 * _GEN_15; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@22.4]
  assign _T_416 = _GEN_11 / _GEN_15; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@23.4]
  assign _T_417 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_418 = _T_417 ? _T_416 : 256'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_419 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_420 = _T_419 ? _T_414 : {{256'd0}, _T_418}; // @[Mux.scala 46:16:@27.4]
  assign _T_421 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_422 = _T_421 ? {{256'd0}, _T_412} : _T_420; // @[Mux.scala 46:16:@29.4]
  assign _T_423 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _GEN_17 = 2'h1 == io_selects_2_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_18 = 2'h2 == io_selects_2_0 ? io_inputs_2 : _GEN_17; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_19 = 2'h3 == io_selects_2_0 ? io_inputs_3 : _GEN_18; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_21 = 2'h1 == io_selects_2_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_22 = 2'h2 == io_selects_2_1 ? io_inputs_2 : _GEN_21; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _GEN_23 = 2'h3 == io_selects_2_1 ? io_inputs_3 : _GEN_22; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _T_428 = _GEN_19 + _GEN_23; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@32.4]
  assign _T_429 = _GEN_19 + _GEN_23; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@33.4]
  assign _T_431 = _GEN_19 * _GEN_23; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@34.4]
  assign _T_433 = _GEN_19 / _GEN_23; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@35.4]
  assign _T_434 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_435 = _T_434 ? _T_433 : 256'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_436 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_437 = _T_436 ? _T_431 : {{256'd0}, _T_435}; // @[Mux.scala 46:16:@39.4]
  assign _T_438 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_439 = _T_438 ? {{256'd0}, _T_429} : _T_437; // @[Mux.scala 46:16:@41.4]
  assign _T_440 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _GEN_25 = 2'h1 == io_selects_3_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_26 = 2'h2 == io_selects_3_0 ? io_inputs_2 : _GEN_25; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_27 = 2'h3 == io_selects_3_0 ? io_inputs_3 : _GEN_26; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_29 = 2'h1 == io_selects_3_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_30 = 2'h2 == io_selects_3_1 ? io_inputs_2 : _GEN_29; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _GEN_31 = 2'h3 == io_selects_3_1 ? io_inputs_3 : _GEN_30; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _T_445 = _GEN_27 + _GEN_31; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@44.4]
  assign _T_446 = _GEN_27 + _GEN_31; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@45.4]
  assign _T_448 = _GEN_27 * _GEN_31; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@46.4]
  assign _T_450 = _GEN_27 / _GEN_31; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@47.4]
  assign _T_451 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_452 = _T_451 ? _T_450 : 256'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_453 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_454 = _T_453 ? _T_448 : {{256'd0}, _T_452}; // @[Mux.scala 46:16:@51.4]
  assign _T_455 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_456 = _T_455 ? {{256'd0}, _T_446} : _T_454; // @[Mux.scala 46:16:@53.4]
  assign _T_457 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _GEN_33 = 2'h1 == io_selects_4_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_34 = 2'h2 == io_selects_4_0 ? io_inputs_2 : _GEN_33; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_35 = 2'h3 == io_selects_4_0 ? io_inputs_3 : _GEN_34; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_37 = 2'h1 == io_selects_4_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_38 = 2'h2 == io_selects_4_1 ? io_inputs_2 : _GEN_37; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _GEN_39 = 2'h3 == io_selects_4_1 ? io_inputs_3 : _GEN_38; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _T_462 = _GEN_35 + _GEN_39; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@56.4]
  assign _T_463 = _GEN_35 + _GEN_39; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@57.4]
  assign _T_465 = _GEN_35 * _GEN_39; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@58.4]
  assign _T_467 = _GEN_35 / _GEN_39; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@59.4]
  assign _T_468 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_469 = _T_468 ? _T_467 : 256'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_470 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_471 = _T_470 ? _T_465 : {{256'd0}, _T_469}; // @[Mux.scala 46:16:@63.4]
  assign _T_472 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_473 = _T_472 ? {{256'd0}, _T_463} : _T_471; // @[Mux.scala 46:16:@65.4]
  assign _T_474 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _GEN_41 = 2'h1 == io_selects_5_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_42 = 2'h2 == io_selects_5_0 ? io_inputs_2 : _GEN_41; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_43 = 2'h3 == io_selects_5_0 ? io_inputs_3 : _GEN_42; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_45 = 2'h1 == io_selects_5_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_46 = 2'h2 == io_selects_5_1 ? io_inputs_2 : _GEN_45; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _GEN_47 = 2'h3 == io_selects_5_1 ? io_inputs_3 : _GEN_46; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _T_479 = _GEN_43 + _GEN_47; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@68.4]
  assign _T_480 = _GEN_43 + _GEN_47; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@69.4]
  assign _T_482 = _GEN_43 * _GEN_47; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@70.4]
  assign _T_484 = _GEN_43 / _GEN_47; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@71.4]
  assign _T_485 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_486 = _T_485 ? _T_484 : 256'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_487 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_488 = _T_487 ? _T_482 : {{256'd0}, _T_486}; // @[Mux.scala 46:16:@75.4]
  assign _T_489 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_490 = _T_489 ? {{256'd0}, _T_480} : _T_488; // @[Mux.scala 46:16:@77.4]
  assign _T_491 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _GEN_49 = 2'h1 == io_selects_6_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_50 = 2'h2 == io_selects_6_0 ? io_inputs_2 : _GEN_49; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_51 = 2'h3 == io_selects_6_0 ? io_inputs_3 : _GEN_50; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_53 = 2'h1 == io_selects_6_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_54 = 2'h2 == io_selects_6_1 ? io_inputs_2 : _GEN_53; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _GEN_55 = 2'h3 == io_selects_6_1 ? io_inputs_3 : _GEN_54; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _T_496 = _GEN_51 + _GEN_55; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@80.4]
  assign _T_497 = _GEN_51 + _GEN_55; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@81.4]
  assign _T_499 = _GEN_51 * _GEN_55; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@82.4]
  assign _T_501 = _GEN_51 / _GEN_55; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@83.4]
  assign _T_502 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_503 = _T_502 ? _T_501 : 256'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_504 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_505 = _T_504 ? _T_499 : {{256'd0}, _T_503}; // @[Mux.scala 46:16:@87.4]
  assign _T_506 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_507 = _T_506 ? {{256'd0}, _T_497} : _T_505; // @[Mux.scala 46:16:@89.4]
  assign _T_508 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _GEN_57 = 2'h1 == io_selects_7_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_58 = 2'h2 == io_selects_7_0 ? io_inputs_2 : _GEN_57; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_59 = 2'h3 == io_selects_7_0 ? io_inputs_3 : _GEN_58; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_61 = 2'h1 == io_selects_7_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_62 = 2'h2 == io_selects_7_1 ? io_inputs_2 : _GEN_61; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _GEN_63 = 2'h3 == io_selects_7_1 ? io_inputs_3 : _GEN_62; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _T_513 = _GEN_59 + _GEN_63; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@92.4]
  assign _T_514 = _GEN_59 + _GEN_63; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 32:53:@93.4]
  assign _T_516 = _GEN_59 * _GEN_63; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 33:58:@94.4]
  assign _T_518 = _GEN_59 / _GEN_63; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 34:56:@95.4]
  assign _T_519 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_520 = _T_519 ? _T_518 : 256'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_521 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_522 = _T_521 ? _T_516 : {{256'd0}, _T_520}; // @[Mux.scala 46:16:@99.4]
  assign _T_523 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_524 = _T_523 ? {{256'd0}, _T_514} : _T_522; // @[Mux.scala 46:16:@101.4]
  assign _T_525 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign io_outputs_0 = _T_537[255:0]; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 23:14:@264.4]
  assign io_outputs_1 = _T_548[255:0]; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 23:14:@265.4]
  assign io_outputs_2 = _T_559[255:0]; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 23:14:@266.4]
  assign io_outputs_3 = _T_570[255:0]; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 23:14:@267.4]
  assign io_outputs_4 = _T_581[255:0]; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 23:14:@268.4]
  assign io_outputs_5 = _T_592[255:0]; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 23:14:@269.4]
  assign io_outputs_6 = _T_603[255:0]; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 23:14:@270.4]
  assign io_outputs_7 = _T_614[255:0]; // @[MuxTest_width_256_inputs_4_outputs_8_pipeline_5s.scala 23:14:@271.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {16{`RANDOM}};
  _T_529 = _RAND_0[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {16{`RANDOM}};
  _T_531 = _RAND_1[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {16{`RANDOM}};
  _T_533 = _RAND_2[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {16{`RANDOM}};
  _T_535 = _RAND_3[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {16{`RANDOM}};
  _T_537 = _RAND_4[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {16{`RANDOM}};
  _T_540 = _RAND_5[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {16{`RANDOM}};
  _T_542 = _RAND_6[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {16{`RANDOM}};
  _T_544 = _RAND_7[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {16{`RANDOM}};
  _T_546 = _RAND_8[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {16{`RANDOM}};
  _T_548 = _RAND_9[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {16{`RANDOM}};
  _T_551 = _RAND_10[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {16{`RANDOM}};
  _T_553 = _RAND_11[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {16{`RANDOM}};
  _T_555 = _RAND_12[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {16{`RANDOM}};
  _T_557 = _RAND_13[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {16{`RANDOM}};
  _T_559 = _RAND_14[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {16{`RANDOM}};
  _T_562 = _RAND_15[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {16{`RANDOM}};
  _T_564 = _RAND_16[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {16{`RANDOM}};
  _T_566 = _RAND_17[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {16{`RANDOM}};
  _T_568 = _RAND_18[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {16{`RANDOM}};
  _T_570 = _RAND_19[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {16{`RANDOM}};
  _T_573 = _RAND_20[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {16{`RANDOM}};
  _T_575 = _RAND_21[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {16{`RANDOM}};
  _T_577 = _RAND_22[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {16{`RANDOM}};
  _T_579 = _RAND_23[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {16{`RANDOM}};
  _T_581 = _RAND_24[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {16{`RANDOM}};
  _T_584 = _RAND_25[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {16{`RANDOM}};
  _T_586 = _RAND_26[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {16{`RANDOM}};
  _T_588 = _RAND_27[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {16{`RANDOM}};
  _T_590 = _RAND_28[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {16{`RANDOM}};
  _T_592 = _RAND_29[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {16{`RANDOM}};
  _T_595 = _RAND_30[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {16{`RANDOM}};
  _T_597 = _RAND_31[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {16{`RANDOM}};
  _T_599 = _RAND_32[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {16{`RANDOM}};
  _T_601 = _RAND_33[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {16{`RANDOM}};
  _T_603 = _RAND_34[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {16{`RANDOM}};
  _T_606 = _RAND_35[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {16{`RANDOM}};
  _T_608 = _RAND_36[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {16{`RANDOM}};
  _T_610 = _RAND_37[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {16{`RANDOM}};
  _T_612 = _RAND_38[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {16{`RANDOM}};
  _T_614 = _RAND_39[511:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_406) begin
      _T_529 <= {{256'd0}, _GEN_3};
    end else begin
      _T_529 <= _T_405;
    end
    _T_531 <= _T_529;
    _T_533 <= _T_531;
    _T_535 <= _T_533;
    _T_537 <= _T_535;
    if (_T_423) begin
      _T_540 <= {{256'd0}, _GEN_11};
    end else begin
      _T_540 <= _T_422;
    end
    _T_542 <= _T_540;
    _T_544 <= _T_542;
    _T_546 <= _T_544;
    _T_548 <= _T_546;
    if (_T_440) begin
      _T_551 <= {{256'd0}, _GEN_19};
    end else begin
      _T_551 <= _T_439;
    end
    _T_553 <= _T_551;
    _T_555 <= _T_553;
    _T_557 <= _T_555;
    _T_559 <= _T_557;
    if (_T_457) begin
      _T_562 <= {{256'd0}, _GEN_27};
    end else begin
      _T_562 <= _T_456;
    end
    _T_564 <= _T_562;
    _T_566 <= _T_564;
    _T_568 <= _T_566;
    _T_570 <= _T_568;
    if (_T_474) begin
      _T_573 <= {{256'd0}, _GEN_35};
    end else begin
      _T_573 <= _T_473;
    end
    _T_575 <= _T_573;
    _T_577 <= _T_575;
    _T_579 <= _T_577;
    _T_581 <= _T_579;
    if (_T_491) begin
      _T_584 <= {{256'd0}, _GEN_43};
    end else begin
      _T_584 <= _T_490;
    end
    _T_586 <= _T_584;
    _T_588 <= _T_586;
    _T_590 <= _T_588;
    _T_592 <= _T_590;
    if (_T_508) begin
      _T_595 <= {{256'd0}, _GEN_51};
    end else begin
      _T_595 <= _T_507;
    end
    _T_597 <= _T_595;
    _T_599 <= _T_597;
    _T_601 <= _T_599;
    _T_603 <= _T_601;
    if (_T_525) begin
      _T_606 <= {{256'd0}, _GEN_59};
    end else begin
      _T_606 <= _T_524;
    end
    _T_608 <= _T_606;
    _T_610 <= _T_608;
    _T_612 <= _T_610;
    _T_614 <= _T_612;
  end
endmodule
