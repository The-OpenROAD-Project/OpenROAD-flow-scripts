../../nangate45/lef/NangateOpenCellLibrary.macro.rect.lef