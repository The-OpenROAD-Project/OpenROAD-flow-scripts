../../nangate45/lef/fakeram45_512x64.lef