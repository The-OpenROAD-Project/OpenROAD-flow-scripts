// Used to silence warnings.
module TAPCELL_ASAP7_75t_R;
endmodule
module FILLERxp5_ASAP7_75t_R;
endmodule
module FILLER_ASAP7_75t_R;
endmodule
module DECAPx1_ASAP7_75t_R;
endmodule
module DECAPx2_ASAP7_75t_R;
endmodule
module DECAPx4_ASAP7_75t_R;
endmodule
module DECAPx6_ASAP7_75t_R;
endmodule
module DECAPx10_ASAP7_75t_R;
endmodule
