../../nangate45/lef/NangateOpenCellLibrary.tech.lef