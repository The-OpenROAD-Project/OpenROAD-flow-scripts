VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram7_256x32
  FOREIGN fakeram7_256x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 4.180 BY 67.200 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.576 0.024 0.600 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.440 0.024 1.464 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.304 0.024 2.328 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.168 0.024 3.192 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.032 0.024 4.056 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.896 0.024 4.920 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.760 0.024 5.784 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.624 0.024 6.648 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.488 0.024 7.512 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.352 0.024 8.376 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.216 0.024 9.240 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.080 0.024 10.104 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.944 0.024 10.968 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.808 0.024 11.832 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.672 0.024 12.696 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.536 0.024 13.560 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.400 0.024 14.424 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.264 0.024 15.288 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.128 0.024 16.152 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 16.992 0.024 17.016 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.856 0.024 17.880 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 18.720 0.024 18.744 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 19.584 0.024 19.608 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 20.448 0.024 20.472 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 21.312 0.024 21.336 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 22.176 0.024 22.200 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.040 0.024 23.064 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.904 0.024 23.928 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 24.768 0.024 24.792 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 25.632 0.024 25.656 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 26.496 0.024 26.520 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.360 0.024 27.384 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 27.648 0.024 27.672 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.512 0.024 28.536 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 29.376 0.024 29.400 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 30.240 0.024 30.264 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.104 0.024 31.128 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 31.968 0.024 31.992 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 32.832 0.024 32.856 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 33.696 0.024 33.720 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 34.560 0.024 34.584 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 35.424 0.024 35.448 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 36.288 0.024 36.312 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 37.152 0.024 37.176 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 38.016 0.024 38.040 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 38.880 0.024 38.904 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 39.744 0.024 39.768 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 40.608 0.024 40.632 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 41.472 0.024 41.496 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 42.336 0.024 42.360 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 43.200 0.024 43.224 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 44.064 0.024 44.088 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 44.928 0.024 44.952 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 45.792 0.024 45.816 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 46.656 0.024 46.680 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 47.520 0.024 47.544 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 48.384 0.024 48.408 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 49.248 0.024 49.272 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 50.112 0.024 50.136 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 50.976 0.024 51.000 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.840 0.024 51.864 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 52.704 0.024 52.728 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 53.568 0.024 53.592 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.432 0.024 54.456 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 54.720 0.024 54.744 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 55.584 0.024 55.608 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 56.448 0.024 56.472 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 57.312 0.024 57.336 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 58.176 0.024 58.200 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.040 0.024 59.064 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 59.904 0.024 59.928 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 60.768 0.024 60.792 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 61.056 0.024 61.080 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 61.920 0.024 61.944 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 62.784 0.024 62.808 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.576 0.528 3.604 0.624 ;
      RECT 0.576 1.296 3.604 1.392 ;
      RECT 0.576 2.064 3.604 2.160 ;
      RECT 0.576 2.832 3.604 2.928 ;
      RECT 0.576 3.600 3.604 3.696 ;
      RECT 0.576 4.368 3.604 4.464 ;
      RECT 0.576 5.136 3.604 5.232 ;
      RECT 0.576 5.904 3.604 6.000 ;
      RECT 0.576 6.672 3.604 6.768 ;
      RECT 0.576 7.440 3.604 7.536 ;
      RECT 0.576 8.208 3.604 8.304 ;
      RECT 0.576 8.976 3.604 9.072 ;
      RECT 0.576 9.744 3.604 9.840 ;
      RECT 0.576 10.512 3.604 10.608 ;
      RECT 0.576 11.280 3.604 11.376 ;
      RECT 0.576 12.048 3.604 12.144 ;
      RECT 0.576 12.816 3.604 12.912 ;
      RECT 0.576 13.584 3.604 13.680 ;
      RECT 0.576 14.352 3.604 14.448 ;
      RECT 0.576 15.120 3.604 15.216 ;
      RECT 0.576 15.888 3.604 15.984 ;
      RECT 0.576 16.656 3.604 16.752 ;
      RECT 0.576 17.424 3.604 17.520 ;
      RECT 0.576 18.192 3.604 18.288 ;
      RECT 0.576 18.960 3.604 19.056 ;
      RECT 0.576 19.728 3.604 19.824 ;
      RECT 0.576 20.496 3.604 20.592 ;
      RECT 0.576 21.264 3.604 21.360 ;
      RECT 0.576 22.032 3.604 22.128 ;
      RECT 0.576 22.800 3.604 22.896 ;
      RECT 0.576 23.568 3.604 23.664 ;
      RECT 0.576 24.336 3.604 24.432 ;
      RECT 0.576 25.104 3.604 25.200 ;
      RECT 0.576 25.872 3.604 25.968 ;
      RECT 0.576 26.640 3.604 26.736 ;
      RECT 0.576 27.408 3.604 27.504 ;
      RECT 0.576 28.176 3.604 28.272 ;
      RECT 0.576 28.944 3.604 29.040 ;
      RECT 0.576 29.712 3.604 29.808 ;
      RECT 0.576 30.480 3.604 30.576 ;
      RECT 0.576 31.248 3.604 31.344 ;
      RECT 0.576 32.016 3.604 32.112 ;
      RECT 0.576 32.784 3.604 32.880 ;
      RECT 0.576 33.552 3.604 33.648 ;
      RECT 0.576 34.320 3.604 34.416 ;
      RECT 0.576 35.088 3.604 35.184 ;
      RECT 0.576 35.856 3.604 35.952 ;
      RECT 0.576 36.624 3.604 36.720 ;
      RECT 0.576 37.392 3.604 37.488 ;
      RECT 0.576 38.160 3.604 38.256 ;
      RECT 0.576 38.928 3.604 39.024 ;
      RECT 0.576 39.696 3.604 39.792 ;
      RECT 0.576 40.464 3.604 40.560 ;
      RECT 0.576 41.232 3.604 41.328 ;
      RECT 0.576 42.000 3.604 42.096 ;
      RECT 0.576 42.768 3.604 42.864 ;
      RECT 0.576 43.536 3.604 43.632 ;
      RECT 0.576 44.304 3.604 44.400 ;
      RECT 0.576 45.072 3.604 45.168 ;
      RECT 0.576 45.840 3.604 45.936 ;
      RECT 0.576 46.608 3.604 46.704 ;
      RECT 0.576 47.376 3.604 47.472 ;
      RECT 0.576 48.144 3.604 48.240 ;
      RECT 0.576 48.912 3.604 49.008 ;
      RECT 0.576 49.680 3.604 49.776 ;
      RECT 0.576 50.448 3.604 50.544 ;
      RECT 0.576 51.216 3.604 51.312 ;
      RECT 0.576 51.984 3.604 52.080 ;
      RECT 0.576 52.752 3.604 52.848 ;
      RECT 0.576 53.520 3.604 53.616 ;
      RECT 0.576 54.288 3.604 54.384 ;
      RECT 0.576 55.056 3.604 55.152 ;
      RECT 0.576 55.824 3.604 55.920 ;
      RECT 0.576 56.592 3.604 56.688 ;
      RECT 0.576 57.360 3.604 57.456 ;
      RECT 0.576 58.128 3.604 58.224 ;
      RECT 0.576 58.896 3.604 58.992 ;
      RECT 0.576 59.664 3.604 59.760 ;
      RECT 0.576 60.432 3.604 60.528 ;
      RECT 0.576 61.200 3.604 61.296 ;
      RECT 0.576 61.968 3.604 62.064 ;
      RECT 0.576 62.736 3.604 62.832 ;
      RECT 0.576 63.504 3.604 63.600 ;
      RECT 0.576 64.272 3.604 64.368 ;
      RECT 0.576 65.040 3.604 65.136 ;
      RECT 0.576 65.808 3.604 65.904 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.576 0.912 3.604 1.008 ;
      RECT 0.576 1.680 3.604 1.776 ;
      RECT 0.576 2.448 3.604 2.544 ;
      RECT 0.576 3.216 3.604 3.312 ;
      RECT 0.576 3.984 3.604 4.080 ;
      RECT 0.576 4.752 3.604 4.848 ;
      RECT 0.576 5.520 3.604 5.616 ;
      RECT 0.576 6.288 3.604 6.384 ;
      RECT 0.576 7.056 3.604 7.152 ;
      RECT 0.576 7.824 3.604 7.920 ;
      RECT 0.576 8.592 3.604 8.688 ;
      RECT 0.576 9.360 3.604 9.456 ;
      RECT 0.576 10.128 3.604 10.224 ;
      RECT 0.576 10.896 3.604 10.992 ;
      RECT 0.576 11.664 3.604 11.760 ;
      RECT 0.576 12.432 3.604 12.528 ;
      RECT 0.576 13.200 3.604 13.296 ;
      RECT 0.576 13.968 3.604 14.064 ;
      RECT 0.576 14.736 3.604 14.832 ;
      RECT 0.576 15.504 3.604 15.600 ;
      RECT 0.576 16.272 3.604 16.368 ;
      RECT 0.576 17.040 3.604 17.136 ;
      RECT 0.576 17.808 3.604 17.904 ;
      RECT 0.576 18.576 3.604 18.672 ;
      RECT 0.576 19.344 3.604 19.440 ;
      RECT 0.576 20.112 3.604 20.208 ;
      RECT 0.576 20.880 3.604 20.976 ;
      RECT 0.576 21.648 3.604 21.744 ;
      RECT 0.576 22.416 3.604 22.512 ;
      RECT 0.576 23.184 3.604 23.280 ;
      RECT 0.576 23.952 3.604 24.048 ;
      RECT 0.576 24.720 3.604 24.816 ;
      RECT 0.576 25.488 3.604 25.584 ;
      RECT 0.576 26.256 3.604 26.352 ;
      RECT 0.576 27.024 3.604 27.120 ;
      RECT 0.576 27.792 3.604 27.888 ;
      RECT 0.576 28.560 3.604 28.656 ;
      RECT 0.576 29.328 3.604 29.424 ;
      RECT 0.576 30.096 3.604 30.192 ;
      RECT 0.576 30.864 3.604 30.960 ;
      RECT 0.576 31.632 3.604 31.728 ;
      RECT 0.576 32.400 3.604 32.496 ;
      RECT 0.576 33.168 3.604 33.264 ;
      RECT 0.576 33.936 3.604 34.032 ;
      RECT 0.576 34.704 3.604 34.800 ;
      RECT 0.576 35.472 3.604 35.568 ;
      RECT 0.576 36.240 3.604 36.336 ;
      RECT 0.576 37.008 3.604 37.104 ;
      RECT 0.576 37.776 3.604 37.872 ;
      RECT 0.576 38.544 3.604 38.640 ;
      RECT 0.576 39.312 3.604 39.408 ;
      RECT 0.576 40.080 3.604 40.176 ;
      RECT 0.576 40.848 3.604 40.944 ;
      RECT 0.576 41.616 3.604 41.712 ;
      RECT 0.576 42.384 3.604 42.480 ;
      RECT 0.576 43.152 3.604 43.248 ;
      RECT 0.576 43.920 3.604 44.016 ;
      RECT 0.576 44.688 3.604 44.784 ;
      RECT 0.576 45.456 3.604 45.552 ;
      RECT 0.576 46.224 3.604 46.320 ;
      RECT 0.576 46.992 3.604 47.088 ;
      RECT 0.576 47.760 3.604 47.856 ;
      RECT 0.576 48.528 3.604 48.624 ;
      RECT 0.576 49.296 3.604 49.392 ;
      RECT 0.576 50.064 3.604 50.160 ;
      RECT 0.576 50.832 3.604 50.928 ;
      RECT 0.576 51.600 3.604 51.696 ;
      RECT 0.576 52.368 3.604 52.464 ;
      RECT 0.576 53.136 3.604 53.232 ;
      RECT 0.576 53.904 3.604 54.000 ;
      RECT 0.576 54.672 3.604 54.768 ;
      RECT 0.576 55.440 3.604 55.536 ;
      RECT 0.576 56.208 3.604 56.304 ;
      RECT 0.576 56.976 3.604 57.072 ;
      RECT 0.576 57.744 3.604 57.840 ;
      RECT 0.576 58.512 3.604 58.608 ;
      RECT 0.576 59.280 3.604 59.376 ;
      RECT 0.576 60.048 3.604 60.144 ;
      RECT 0.576 60.816 3.604 60.912 ;
      RECT 0.576 61.584 3.604 61.680 ;
      RECT 0.576 62.352 3.604 62.448 ;
      RECT 0.576 63.120 3.604 63.216 ;
      RECT 0.576 63.888 3.604 63.984 ;
      RECT 0.576 64.656 3.604 64.752 ;
      RECT 0.576 65.424 3.604 65.520 ;
      RECT 0.576 66.192 3.604 66.288 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 4.180 67.200 ;
    LAYER M2 ;
    RECT 0 0 4.180 67.200 ;
    LAYER M3 ;
    RECT 0 0 4.180 67.200 ;
    LAYER M4 ;
    RECT 0.024 0 0.576 67.200 ;
    RECT 3.604 0 4.180 67.200 ;
    RECT 0.576 0.000 3.604 0.528 ;
    RECT 0.576 0.624 3.604 0.912 ;
    RECT 0.576 1.008 3.604 1.296 ;
    RECT 0.576 1.392 3.604 1.680 ;
    RECT 0.576 1.776 3.604 2.064 ;
    RECT 0.576 2.160 3.604 2.448 ;
    RECT 0.576 2.544 3.604 2.832 ;
    RECT 0.576 2.928 3.604 3.216 ;
    RECT 0.576 3.312 3.604 3.600 ;
    RECT 0.576 3.696 3.604 3.984 ;
    RECT 0.576 4.080 3.604 4.368 ;
    RECT 0.576 4.464 3.604 4.752 ;
    RECT 0.576 4.848 3.604 5.136 ;
    RECT 0.576 5.232 3.604 5.520 ;
    RECT 0.576 5.616 3.604 5.904 ;
    RECT 0.576 6.000 3.604 6.288 ;
    RECT 0.576 6.384 3.604 6.672 ;
    RECT 0.576 6.768 3.604 7.056 ;
    RECT 0.576 7.152 3.604 7.440 ;
    RECT 0.576 7.536 3.604 7.824 ;
    RECT 0.576 7.920 3.604 8.208 ;
    RECT 0.576 8.304 3.604 8.592 ;
    RECT 0.576 8.688 3.604 8.976 ;
    RECT 0.576 9.072 3.604 9.360 ;
    RECT 0.576 9.456 3.604 9.744 ;
    RECT 0.576 9.840 3.604 10.128 ;
    RECT 0.576 10.224 3.604 10.512 ;
    RECT 0.576 10.608 3.604 10.896 ;
    RECT 0.576 10.992 3.604 11.280 ;
    RECT 0.576 11.376 3.604 11.664 ;
    RECT 0.576 11.760 3.604 12.048 ;
    RECT 0.576 12.144 3.604 12.432 ;
    RECT 0.576 12.528 3.604 12.816 ;
    RECT 0.576 12.912 3.604 13.200 ;
    RECT 0.576 13.296 3.604 13.584 ;
    RECT 0.576 13.680 3.604 13.968 ;
    RECT 0.576 14.064 3.604 14.352 ;
    RECT 0.576 14.448 3.604 14.736 ;
    RECT 0.576 14.832 3.604 15.120 ;
    RECT 0.576 15.216 3.604 15.504 ;
    RECT 0.576 15.600 3.604 15.888 ;
    RECT 0.576 15.984 3.604 16.272 ;
    RECT 0.576 16.368 3.604 16.656 ;
    RECT 0.576 16.752 3.604 17.040 ;
    RECT 0.576 17.136 3.604 17.424 ;
    RECT 0.576 17.520 3.604 17.808 ;
    RECT 0.576 17.904 3.604 18.192 ;
    RECT 0.576 18.288 3.604 18.576 ;
    RECT 0.576 18.672 3.604 18.960 ;
    RECT 0.576 19.056 3.604 19.344 ;
    RECT 0.576 19.440 3.604 19.728 ;
    RECT 0.576 19.824 3.604 20.112 ;
    RECT 0.576 20.208 3.604 20.496 ;
    RECT 0.576 20.592 3.604 20.880 ;
    RECT 0.576 20.976 3.604 21.264 ;
    RECT 0.576 21.360 3.604 21.648 ;
    RECT 0.576 21.744 3.604 22.032 ;
    RECT 0.576 22.128 3.604 22.416 ;
    RECT 0.576 22.512 3.604 22.800 ;
    RECT 0.576 22.896 3.604 23.184 ;
    RECT 0.576 23.280 3.604 23.568 ;
    RECT 0.576 23.664 3.604 23.952 ;
    RECT 0.576 24.048 3.604 24.336 ;
    RECT 0.576 24.432 3.604 24.720 ;
    RECT 0.576 24.816 3.604 25.104 ;
    RECT 0.576 25.200 3.604 25.488 ;
    RECT 0.576 25.584 3.604 25.872 ;
    RECT 0.576 25.968 3.604 26.256 ;
    RECT 0.576 26.352 3.604 26.640 ;
    RECT 0.576 26.736 3.604 27.024 ;
    RECT 0.576 27.120 3.604 27.408 ;
    RECT 0.576 27.504 3.604 27.792 ;
    RECT 0.576 27.888 3.604 28.176 ;
    RECT 0.576 28.272 3.604 28.560 ;
    RECT 0.576 28.656 3.604 28.944 ;
    RECT 0.576 29.040 3.604 29.328 ;
    RECT 0.576 29.424 3.604 29.712 ;
    RECT 0.576 29.808 3.604 30.096 ;
    RECT 0.576 30.192 3.604 30.480 ;
    RECT 0.576 30.576 3.604 30.864 ;
    RECT 0.576 30.960 3.604 31.248 ;
    RECT 0.576 31.344 3.604 31.632 ;
    RECT 0.576 31.728 3.604 32.016 ;
    RECT 0.576 32.112 3.604 32.400 ;
    RECT 0.576 32.496 3.604 32.784 ;
    RECT 0.576 32.880 3.604 33.168 ;
    RECT 0.576 33.264 3.604 33.552 ;
    RECT 0.576 33.648 3.604 33.936 ;
    RECT 0.576 34.032 3.604 34.320 ;
    RECT 0.576 34.416 3.604 34.704 ;
    RECT 0.576 34.800 3.604 35.088 ;
    RECT 0.576 35.184 3.604 35.472 ;
    RECT 0.576 35.568 3.604 35.856 ;
    RECT 0.576 35.952 3.604 36.240 ;
    RECT 0.576 36.336 3.604 36.624 ;
    RECT 0.576 36.720 3.604 37.008 ;
    RECT 0.576 37.104 3.604 37.392 ;
    RECT 0.576 37.488 3.604 37.776 ;
    RECT 0.576 37.872 3.604 38.160 ;
    RECT 0.576 38.256 3.604 38.544 ;
    RECT 0.576 38.640 3.604 38.928 ;
    RECT 0.576 39.024 3.604 39.312 ;
    RECT 0.576 39.408 3.604 39.696 ;
    RECT 0.576 39.792 3.604 40.080 ;
    RECT 0.576 40.176 3.604 40.464 ;
    RECT 0.576 40.560 3.604 40.848 ;
    RECT 0.576 40.944 3.604 41.232 ;
    RECT 0.576 41.328 3.604 41.616 ;
    RECT 0.576 41.712 3.604 42.000 ;
    RECT 0.576 42.096 3.604 42.384 ;
    RECT 0.576 42.480 3.604 42.768 ;
    RECT 0.576 42.864 3.604 43.152 ;
    RECT 0.576 43.248 3.604 43.536 ;
    RECT 0.576 43.632 3.604 43.920 ;
    RECT 0.576 44.016 3.604 44.304 ;
    RECT 0.576 44.400 3.604 44.688 ;
    RECT 0.576 44.784 3.604 45.072 ;
    RECT 0.576 45.168 3.604 45.456 ;
    RECT 0.576 45.552 3.604 45.840 ;
    RECT 0.576 45.936 3.604 46.224 ;
    RECT 0.576 46.320 3.604 46.608 ;
    RECT 0.576 46.704 3.604 46.992 ;
    RECT 0.576 47.088 3.604 47.376 ;
    RECT 0.576 47.472 3.604 47.760 ;
    RECT 0.576 47.856 3.604 48.144 ;
    RECT 0.576 48.240 3.604 48.528 ;
    RECT 0.576 48.624 3.604 48.912 ;
    RECT 0.576 49.008 3.604 49.296 ;
    RECT 0.576 49.392 3.604 49.680 ;
    RECT 0.576 49.776 3.604 50.064 ;
    RECT 0.576 50.160 3.604 50.448 ;
    RECT 0.576 50.544 3.604 50.832 ;
    RECT 0.576 50.928 3.604 51.216 ;
    RECT 0.576 51.312 3.604 51.600 ;
    RECT 0.576 51.696 3.604 51.984 ;
    RECT 0.576 52.080 3.604 52.368 ;
    RECT 0.576 52.464 3.604 52.752 ;
    RECT 0.576 52.848 3.604 53.136 ;
    RECT 0.576 53.232 3.604 53.520 ;
    RECT 0.576 53.616 3.604 53.904 ;
    RECT 0.576 54.000 3.604 54.288 ;
    RECT 0.576 54.384 3.604 54.672 ;
    RECT 0.576 54.768 3.604 55.056 ;
    RECT 0.576 55.152 3.604 55.440 ;
    RECT 0.576 55.536 3.604 55.824 ;
    RECT 0.576 55.920 3.604 56.208 ;
    RECT 0.576 56.304 3.604 56.592 ;
    RECT 0.576 56.688 3.604 56.976 ;
    RECT 0.576 57.072 3.604 57.360 ;
    RECT 0.576 57.456 3.604 57.744 ;
    RECT 0.576 57.840 3.604 58.128 ;
    RECT 0.576 58.224 3.604 58.512 ;
    RECT 0.576 58.608 3.604 58.896 ;
    RECT 0.576 58.992 3.604 59.280 ;
    RECT 0.576 59.376 3.604 59.664 ;
    RECT 0.576 59.760 3.604 60.048 ;
    RECT 0.576 60.144 3.604 60.432 ;
    RECT 0.576 60.528 3.604 60.816 ;
    RECT 0.576 60.912 3.604 61.200 ;
    RECT 0.576 61.296 3.604 61.584 ;
    RECT 0.576 61.680 3.604 61.968 ;
    RECT 0.576 62.064 3.604 62.352 ;
    RECT 0.576 62.448 3.604 62.736 ;
    RECT 0.576 62.832 3.604 63.120 ;
    RECT 0.576 63.216 3.604 63.504 ;
    RECT 0.576 63.600 3.604 63.888 ;
    RECT 0.576 63.984 3.604 64.272 ;
    RECT 0.576 64.368 3.604 64.656 ;
    RECT 0.576 64.752 3.604 65.040 ;
    RECT 0.576 65.136 3.604 65.424 ;
    RECT 0.576 65.520 3.604 65.808 ;
    RECT 0.576 65.904 3.604 66.192 ;
    RECT 0.576 66.288 3.604 67.200 ;
    RECT 0 0.000 0.024 0.576 ;
    RECT 0 0.600 0.024 1.440 ;
    RECT 0 1.464 0.024 2.304 ;
    RECT 0 2.328 0.024 3.168 ;
    RECT 0 3.192 0.024 4.032 ;
    RECT 0 4.056 0.024 4.896 ;
    RECT 0 4.920 0.024 5.760 ;
    RECT 0 5.784 0.024 6.624 ;
    RECT 0 6.648 0.024 7.488 ;
    RECT 0 7.512 0.024 8.352 ;
    RECT 0 8.376 0.024 9.216 ;
    RECT 0 9.240 0.024 10.080 ;
    RECT 0 10.104 0.024 10.944 ;
    RECT 0 10.968 0.024 11.808 ;
    RECT 0 11.832 0.024 12.672 ;
    RECT 0 12.696 0.024 13.536 ;
    RECT 0 13.560 0.024 14.400 ;
    RECT 0 14.424 0.024 15.264 ;
    RECT 0 15.288 0.024 16.128 ;
    RECT 0 16.152 0.024 16.992 ;
    RECT 0 17.016 0.024 17.856 ;
    RECT 0 17.880 0.024 18.720 ;
    RECT 0 18.744 0.024 19.584 ;
    RECT 0 19.608 0.024 20.448 ;
    RECT 0 20.472 0.024 21.312 ;
    RECT 0 21.336 0.024 22.176 ;
    RECT 0 22.200 0.024 23.040 ;
    RECT 0 23.064 0.024 23.904 ;
    RECT 0 23.928 0.024 24.768 ;
    RECT 0 24.792 0.024 25.632 ;
    RECT 0 25.656 0.024 26.496 ;
    RECT 0 26.520 0.024 27.360 ;
    RECT 0 27.384 0.024 27.648 ;
    RECT 0 27.672 0.024 28.512 ;
    RECT 0 28.536 0.024 29.376 ;
    RECT 0 29.400 0.024 30.240 ;
    RECT 0 30.264 0.024 31.104 ;
    RECT 0 31.128 0.024 31.968 ;
    RECT 0 31.992 0.024 32.832 ;
    RECT 0 32.856 0.024 33.696 ;
    RECT 0 33.720 0.024 34.560 ;
    RECT 0 34.584 0.024 35.424 ;
    RECT 0 35.448 0.024 36.288 ;
    RECT 0 36.312 0.024 37.152 ;
    RECT 0 37.176 0.024 38.016 ;
    RECT 0 38.040 0.024 38.880 ;
    RECT 0 38.904 0.024 39.744 ;
    RECT 0 39.768 0.024 40.608 ;
    RECT 0 40.632 0.024 41.472 ;
    RECT 0 41.496 0.024 42.336 ;
    RECT 0 42.360 0.024 43.200 ;
    RECT 0 43.224 0.024 44.064 ;
    RECT 0 44.088 0.024 44.928 ;
    RECT 0 44.952 0.024 45.792 ;
    RECT 0 45.816 0.024 46.656 ;
    RECT 0 46.680 0.024 47.520 ;
    RECT 0 47.544 0.024 48.384 ;
    RECT 0 48.408 0.024 49.248 ;
    RECT 0 49.272 0.024 50.112 ;
    RECT 0 50.136 0.024 50.976 ;
    RECT 0 51.000 0.024 51.840 ;
    RECT 0 51.864 0.024 52.704 ;
    RECT 0 52.728 0.024 53.568 ;
    RECT 0 53.592 0.024 54.432 ;
    RECT 0 54.456 0.024 54.720 ;
    RECT 0 54.744 0.024 55.584 ;
    RECT 0 55.608 0.024 56.448 ;
    RECT 0 56.472 0.024 57.312 ;
    RECT 0 57.336 0.024 58.176 ;
    RECT 0 58.200 0.024 59.040 ;
    RECT 0 59.064 0.024 59.904 ;
    RECT 0 59.928 0.024 60.768 ;
    RECT 0 60.792 0.024 61.632 ;
    RECT 0 61.656 0.024 62.496 ;
    RECT 0 62.520 0.024 63.360 ;
    RECT 0 63.384 0.024 64.224 ;
    RECT 0 64.248 0.024 65.088 ;
    RECT 0 65.112 0.024 65.952 ;
    RECT 0 65.976 0.024 66.816 ;
    RECT 0 66.840 0.024 67.680 ;
    RECT 0 67.704 0.024 68.544 ;
    RECT 0 68.568 0.024 69.408 ;
    RECT 0 69.432 0.024 70.272 ;
    RECT 0 70.296 0.024 71.136 ;
    RECT 0 71.160 0.024 72.000 ;
    RECT 0 72.024 0.024 72.864 ;
    RECT 0 72.888 0.024 73.728 ;
    RECT 0 73.752 0.024 74.592 ;
    RECT 0 74.616 0.024 75.456 ;
    RECT 0 75.480 0.024 76.320 ;
    RECT 0 76.344 0.024 77.184 ;
    RECT 0 77.208 0.024 78.048 ;
    RECT 0 78.072 0.024 78.912 ;
    RECT 0 78.936 0.024 79.776 ;
    RECT 0 79.800 0.024 80.640 ;
    RECT 0 80.664 0.024 81.504 ;
    RECT 0 81.528 0.024 81.792 ;
    RECT 0 81.816 0.024 82.656 ;
    RECT 0 82.680 0.024 83.520 ;
    RECT 0 83.544 0.024 84.384 ;
    RECT 0 84.408 0.024 85.248 ;
    RECT 0 85.272 0.024 86.112 ;
    RECT 0 86.136 0.024 86.976 ;
    RECT 0 87.000 0.024 87.840 ;
    RECT 0 87.864 0.024 88.128 ;
    RECT 0 88.152 0.024 88.992 ;
    RECT 0 89.016 0.024 89.856 ;
    RECT 0 89.880 0.024 67.200 ;
    LAYER OVERLAP ;
    RECT 0 0 4.180 67.200 ;
  END
END fakeram7_256x32

END LIBRARY
