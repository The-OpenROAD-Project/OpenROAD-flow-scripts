module MuxTest_width_16_inputs_1_outputs_16_pipeline_5( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [2:0]  io_operation_0, // @[:@6.4]
  input  [2:0]  io_operation_1, // @[:@6.4]
  input  [2:0]  io_operation_2, // @[:@6.4]
  input  [2:0]  io_operation_3, // @[:@6.4]
  input  [2:0]  io_operation_4, // @[:@6.4]
  input  [2:0]  io_operation_5, // @[:@6.4]
  input  [2:0]  io_operation_6, // @[:@6.4]
  input  [2:0]  io_operation_7, // @[:@6.4]
  input  [2:0]  io_operation_8, // @[:@6.4]
  input  [2:0]  io_operation_9, // @[:@6.4]
  input  [2:0]  io_operation_10, // @[:@6.4]
  input  [2:0]  io_operation_11, // @[:@6.4]
  input  [2:0]  io_operation_12, // @[:@6.4]
  input  [2:0]  io_operation_13, // @[:@6.4]
  input  [2:0]  io_operation_14, // @[:@6.4]
  input  [2:0]  io_operation_15, // @[:@6.4]
  input  [15:0] io_inputs_0, // @[:@6.4]
  output [15:0] io_outputs_0, // @[:@6.4]
  output [15:0] io_outputs_1, // @[:@6.4]
  output [15:0] io_outputs_2, // @[:@6.4]
  output [15:0] io_outputs_3, // @[:@6.4]
  output [15:0] io_outputs_4, // @[:@6.4]
  output [15:0] io_outputs_5, // @[:@6.4]
  output [15:0] io_outputs_6, // @[:@6.4]
  output [15:0] io_outputs_7, // @[:@6.4]
  output [15:0] io_outputs_8, // @[:@6.4]
  output [15:0] io_outputs_9, // @[:@6.4]
  output [15:0] io_outputs_10, // @[:@6.4]
  output [15:0] io_outputs_11, // @[:@6.4]
  output [15:0] io_outputs_12, // @[:@6.4]
  output [15:0] io_outputs_13, // @[:@6.4]
  output [15:0] io_outputs_14, // @[:@6.4]
  output [15:0] io_outputs_15 // @[:@6.4]
);
  wire [16:0] _T_724; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 32:53:@8.4]
  wire [15:0] _T_725; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 32:53:@9.4]
  wire [31:0] _T_727; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 33:58:@10.4]
  wire [15:0] _T_729; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 34:56:@11.4]
  wire  _T_730; // @[Mux.scala 46:19:@12.4]
  wire [15:0] _T_731; // @[Mux.scala 46:16:@13.4]
  wire  _T_732; // @[Mux.scala 46:19:@14.4]
  wire [31:0] _T_733; // @[Mux.scala 46:16:@15.4]
  wire  _T_734; // @[Mux.scala 46:19:@16.4]
  wire [31:0] _T_735; // @[Mux.scala 46:16:@17.4]
  wire  _T_736; // @[Mux.scala 46:19:@18.4]
  wire  _T_747; // @[Mux.scala 46:19:@24.4]
  wire [15:0] _T_748; // @[Mux.scala 46:16:@25.4]
  wire  _T_749; // @[Mux.scala 46:19:@26.4]
  wire [31:0] _T_750; // @[Mux.scala 46:16:@27.4]
  wire  _T_751; // @[Mux.scala 46:19:@28.4]
  wire [31:0] _T_752; // @[Mux.scala 46:16:@29.4]
  wire  _T_753; // @[Mux.scala 46:19:@30.4]
  wire  _T_764; // @[Mux.scala 46:19:@36.4]
  wire [15:0] _T_765; // @[Mux.scala 46:16:@37.4]
  wire  _T_766; // @[Mux.scala 46:19:@38.4]
  wire [31:0] _T_767; // @[Mux.scala 46:16:@39.4]
  wire  _T_768; // @[Mux.scala 46:19:@40.4]
  wire [31:0] _T_769; // @[Mux.scala 46:16:@41.4]
  wire  _T_770; // @[Mux.scala 46:19:@42.4]
  wire  _T_781; // @[Mux.scala 46:19:@48.4]
  wire [15:0] _T_782; // @[Mux.scala 46:16:@49.4]
  wire  _T_783; // @[Mux.scala 46:19:@50.4]
  wire [31:0] _T_784; // @[Mux.scala 46:16:@51.4]
  wire  _T_785; // @[Mux.scala 46:19:@52.4]
  wire [31:0] _T_786; // @[Mux.scala 46:16:@53.4]
  wire  _T_787; // @[Mux.scala 46:19:@54.4]
  wire  _T_798; // @[Mux.scala 46:19:@60.4]
  wire [15:0] _T_799; // @[Mux.scala 46:16:@61.4]
  wire  _T_800; // @[Mux.scala 46:19:@62.4]
  wire [31:0] _T_801; // @[Mux.scala 46:16:@63.4]
  wire  _T_802; // @[Mux.scala 46:19:@64.4]
  wire [31:0] _T_803; // @[Mux.scala 46:16:@65.4]
  wire  _T_804; // @[Mux.scala 46:19:@66.4]
  wire  _T_815; // @[Mux.scala 46:19:@72.4]
  wire [15:0] _T_816; // @[Mux.scala 46:16:@73.4]
  wire  _T_817; // @[Mux.scala 46:19:@74.4]
  wire [31:0] _T_818; // @[Mux.scala 46:16:@75.4]
  wire  _T_819; // @[Mux.scala 46:19:@76.4]
  wire [31:0] _T_820; // @[Mux.scala 46:16:@77.4]
  wire  _T_821; // @[Mux.scala 46:19:@78.4]
  wire  _T_832; // @[Mux.scala 46:19:@84.4]
  wire [15:0] _T_833; // @[Mux.scala 46:16:@85.4]
  wire  _T_834; // @[Mux.scala 46:19:@86.4]
  wire [31:0] _T_835; // @[Mux.scala 46:16:@87.4]
  wire  _T_836; // @[Mux.scala 46:19:@88.4]
  wire [31:0] _T_837; // @[Mux.scala 46:16:@89.4]
  wire  _T_838; // @[Mux.scala 46:19:@90.4]
  wire  _T_849; // @[Mux.scala 46:19:@96.4]
  wire [15:0] _T_850; // @[Mux.scala 46:16:@97.4]
  wire  _T_851; // @[Mux.scala 46:19:@98.4]
  wire [31:0] _T_852; // @[Mux.scala 46:16:@99.4]
  wire  _T_853; // @[Mux.scala 46:19:@100.4]
  wire [31:0] _T_854; // @[Mux.scala 46:16:@101.4]
  wire  _T_855; // @[Mux.scala 46:19:@102.4]
  wire  _T_866; // @[Mux.scala 46:19:@108.4]
  wire [15:0] _T_867; // @[Mux.scala 46:16:@109.4]
  wire  _T_868; // @[Mux.scala 46:19:@110.4]
  wire [31:0] _T_869; // @[Mux.scala 46:16:@111.4]
  wire  _T_870; // @[Mux.scala 46:19:@112.4]
  wire [31:0] _T_871; // @[Mux.scala 46:16:@113.4]
  wire  _T_872; // @[Mux.scala 46:19:@114.4]
  wire  _T_883; // @[Mux.scala 46:19:@120.4]
  wire [15:0] _T_884; // @[Mux.scala 46:16:@121.4]
  wire  _T_885; // @[Mux.scala 46:19:@122.4]
  wire [31:0] _T_886; // @[Mux.scala 46:16:@123.4]
  wire  _T_887; // @[Mux.scala 46:19:@124.4]
  wire [31:0] _T_888; // @[Mux.scala 46:16:@125.4]
  wire  _T_889; // @[Mux.scala 46:19:@126.4]
  wire  _T_900; // @[Mux.scala 46:19:@132.4]
  wire [15:0] _T_901; // @[Mux.scala 46:16:@133.4]
  wire  _T_902; // @[Mux.scala 46:19:@134.4]
  wire [31:0] _T_903; // @[Mux.scala 46:16:@135.4]
  wire  _T_904; // @[Mux.scala 46:19:@136.4]
  wire [31:0] _T_905; // @[Mux.scala 46:16:@137.4]
  wire  _T_906; // @[Mux.scala 46:19:@138.4]
  wire  _T_917; // @[Mux.scala 46:19:@144.4]
  wire [15:0] _T_918; // @[Mux.scala 46:16:@145.4]
  wire  _T_919; // @[Mux.scala 46:19:@146.4]
  wire [31:0] _T_920; // @[Mux.scala 46:16:@147.4]
  wire  _T_921; // @[Mux.scala 46:19:@148.4]
  wire [31:0] _T_922; // @[Mux.scala 46:16:@149.4]
  wire  _T_923; // @[Mux.scala 46:19:@150.4]
  wire  _T_934; // @[Mux.scala 46:19:@156.4]
  wire [15:0] _T_935; // @[Mux.scala 46:16:@157.4]
  wire  _T_936; // @[Mux.scala 46:19:@158.4]
  wire [31:0] _T_937; // @[Mux.scala 46:16:@159.4]
  wire  _T_938; // @[Mux.scala 46:19:@160.4]
  wire [31:0] _T_939; // @[Mux.scala 46:16:@161.4]
  wire  _T_940; // @[Mux.scala 46:19:@162.4]
  wire  _T_951; // @[Mux.scala 46:19:@168.4]
  wire [15:0] _T_952; // @[Mux.scala 46:16:@169.4]
  wire  _T_953; // @[Mux.scala 46:19:@170.4]
  wire [31:0] _T_954; // @[Mux.scala 46:16:@171.4]
  wire  _T_955; // @[Mux.scala 46:19:@172.4]
  wire [31:0] _T_956; // @[Mux.scala 46:16:@173.4]
  wire  _T_957; // @[Mux.scala 46:19:@174.4]
  wire  _T_968; // @[Mux.scala 46:19:@180.4]
  wire [15:0] _T_969; // @[Mux.scala 46:16:@181.4]
  wire  _T_970; // @[Mux.scala 46:19:@182.4]
  wire [31:0] _T_971; // @[Mux.scala 46:16:@183.4]
  wire  _T_972; // @[Mux.scala 46:19:@184.4]
  wire [31:0] _T_973; // @[Mux.scala 46:16:@185.4]
  wire  _T_974; // @[Mux.scala 46:19:@186.4]
  wire  _T_985; // @[Mux.scala 46:19:@192.4]
  wire [15:0] _T_986; // @[Mux.scala 46:16:@193.4]
  wire  _T_987; // @[Mux.scala 46:19:@194.4]
  wire [31:0] _T_988; // @[Mux.scala 46:16:@195.4]
  wire  _T_989; // @[Mux.scala 46:19:@196.4]
  wire [31:0] _T_990; // @[Mux.scala 46:16:@197.4]
  wire  _T_991; // @[Mux.scala 46:19:@198.4]
  reg [31:0] _T_995; // @[Reg.scala 11:16:@200.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_997; // @[Reg.scala 11:16:@204.4]
  reg [31:0] _RAND_1;
  reg [31:0] _T_999; // @[Reg.scala 11:16:@208.4]
  reg [31:0] _RAND_2;
  reg [31:0] _T_1001; // @[Reg.scala 11:16:@212.4]
  reg [31:0] _RAND_3;
  reg [31:0] _T_1003; // @[Reg.scala 11:16:@216.4]
  reg [31:0] _RAND_4;
  reg [31:0] _T_1006; // @[Reg.scala 11:16:@220.4]
  reg [31:0] _RAND_5;
  reg [31:0] _T_1008; // @[Reg.scala 11:16:@224.4]
  reg [31:0] _RAND_6;
  reg [31:0] _T_1010; // @[Reg.scala 11:16:@228.4]
  reg [31:0] _RAND_7;
  reg [31:0] _T_1012; // @[Reg.scala 11:16:@232.4]
  reg [31:0] _RAND_8;
  reg [31:0] _T_1014; // @[Reg.scala 11:16:@236.4]
  reg [31:0] _RAND_9;
  reg [31:0] _T_1017; // @[Reg.scala 11:16:@240.4]
  reg [31:0] _RAND_10;
  reg [31:0] _T_1019; // @[Reg.scala 11:16:@244.4]
  reg [31:0] _RAND_11;
  reg [31:0] _T_1021; // @[Reg.scala 11:16:@248.4]
  reg [31:0] _RAND_12;
  reg [31:0] _T_1023; // @[Reg.scala 11:16:@252.4]
  reg [31:0] _RAND_13;
  reg [31:0] _T_1025; // @[Reg.scala 11:16:@256.4]
  reg [31:0] _RAND_14;
  reg [31:0] _T_1028; // @[Reg.scala 11:16:@260.4]
  reg [31:0] _RAND_15;
  reg [31:0] _T_1030; // @[Reg.scala 11:16:@264.4]
  reg [31:0] _RAND_16;
  reg [31:0] _T_1032; // @[Reg.scala 11:16:@268.4]
  reg [31:0] _RAND_17;
  reg [31:0] _T_1034; // @[Reg.scala 11:16:@272.4]
  reg [31:0] _RAND_18;
  reg [31:0] _T_1036; // @[Reg.scala 11:16:@276.4]
  reg [31:0] _RAND_19;
  reg [31:0] _T_1039; // @[Reg.scala 11:16:@280.4]
  reg [31:0] _RAND_20;
  reg [31:0] _T_1041; // @[Reg.scala 11:16:@284.4]
  reg [31:0] _RAND_21;
  reg [31:0] _T_1043; // @[Reg.scala 11:16:@288.4]
  reg [31:0] _RAND_22;
  reg [31:0] _T_1045; // @[Reg.scala 11:16:@292.4]
  reg [31:0] _RAND_23;
  reg [31:0] _T_1047; // @[Reg.scala 11:16:@296.4]
  reg [31:0] _RAND_24;
  reg [31:0] _T_1050; // @[Reg.scala 11:16:@300.4]
  reg [31:0] _RAND_25;
  reg [31:0] _T_1052; // @[Reg.scala 11:16:@304.4]
  reg [31:0] _RAND_26;
  reg [31:0] _T_1054; // @[Reg.scala 11:16:@308.4]
  reg [31:0] _RAND_27;
  reg [31:0] _T_1056; // @[Reg.scala 11:16:@312.4]
  reg [31:0] _RAND_28;
  reg [31:0] _T_1058; // @[Reg.scala 11:16:@316.4]
  reg [31:0] _RAND_29;
  reg [31:0] _T_1061; // @[Reg.scala 11:16:@320.4]
  reg [31:0] _RAND_30;
  reg [31:0] _T_1063; // @[Reg.scala 11:16:@324.4]
  reg [31:0] _RAND_31;
  reg [31:0] _T_1065; // @[Reg.scala 11:16:@328.4]
  reg [31:0] _RAND_32;
  reg [31:0] _T_1067; // @[Reg.scala 11:16:@332.4]
  reg [31:0] _RAND_33;
  reg [31:0] _T_1069; // @[Reg.scala 11:16:@336.4]
  reg [31:0] _RAND_34;
  reg [31:0] _T_1072; // @[Reg.scala 11:16:@340.4]
  reg [31:0] _RAND_35;
  reg [31:0] _T_1074; // @[Reg.scala 11:16:@344.4]
  reg [31:0] _RAND_36;
  reg [31:0] _T_1076; // @[Reg.scala 11:16:@348.4]
  reg [31:0] _RAND_37;
  reg [31:0] _T_1078; // @[Reg.scala 11:16:@352.4]
  reg [31:0] _RAND_38;
  reg [31:0] _T_1080; // @[Reg.scala 11:16:@356.4]
  reg [31:0] _RAND_39;
  reg [31:0] _T_1083; // @[Reg.scala 11:16:@360.4]
  reg [31:0] _RAND_40;
  reg [31:0] _T_1085; // @[Reg.scala 11:16:@364.4]
  reg [31:0] _RAND_41;
  reg [31:0] _T_1087; // @[Reg.scala 11:16:@368.4]
  reg [31:0] _RAND_42;
  reg [31:0] _T_1089; // @[Reg.scala 11:16:@372.4]
  reg [31:0] _RAND_43;
  reg [31:0] _T_1091; // @[Reg.scala 11:16:@376.4]
  reg [31:0] _RAND_44;
  reg [31:0] _T_1094; // @[Reg.scala 11:16:@380.4]
  reg [31:0] _RAND_45;
  reg [31:0] _T_1096; // @[Reg.scala 11:16:@384.4]
  reg [31:0] _RAND_46;
  reg [31:0] _T_1098; // @[Reg.scala 11:16:@388.4]
  reg [31:0] _RAND_47;
  reg [31:0] _T_1100; // @[Reg.scala 11:16:@392.4]
  reg [31:0] _RAND_48;
  reg [31:0] _T_1102; // @[Reg.scala 11:16:@396.4]
  reg [31:0] _RAND_49;
  reg [31:0] _T_1105; // @[Reg.scala 11:16:@400.4]
  reg [31:0] _RAND_50;
  reg [31:0] _T_1107; // @[Reg.scala 11:16:@404.4]
  reg [31:0] _RAND_51;
  reg [31:0] _T_1109; // @[Reg.scala 11:16:@408.4]
  reg [31:0] _RAND_52;
  reg [31:0] _T_1111; // @[Reg.scala 11:16:@412.4]
  reg [31:0] _RAND_53;
  reg [31:0] _T_1113; // @[Reg.scala 11:16:@416.4]
  reg [31:0] _RAND_54;
  reg [31:0] _T_1116; // @[Reg.scala 11:16:@420.4]
  reg [31:0] _RAND_55;
  reg [31:0] _T_1118; // @[Reg.scala 11:16:@424.4]
  reg [31:0] _RAND_56;
  reg [31:0] _T_1120; // @[Reg.scala 11:16:@428.4]
  reg [31:0] _RAND_57;
  reg [31:0] _T_1122; // @[Reg.scala 11:16:@432.4]
  reg [31:0] _RAND_58;
  reg [31:0] _T_1124; // @[Reg.scala 11:16:@436.4]
  reg [31:0] _RAND_59;
  reg [31:0] _T_1127; // @[Reg.scala 11:16:@440.4]
  reg [31:0] _RAND_60;
  reg [31:0] _T_1129; // @[Reg.scala 11:16:@444.4]
  reg [31:0] _RAND_61;
  reg [31:0] _T_1131; // @[Reg.scala 11:16:@448.4]
  reg [31:0] _RAND_62;
  reg [31:0] _T_1133; // @[Reg.scala 11:16:@452.4]
  reg [31:0] _RAND_63;
  reg [31:0] _T_1135; // @[Reg.scala 11:16:@456.4]
  reg [31:0] _RAND_64;
  reg [31:0] _T_1138; // @[Reg.scala 11:16:@460.4]
  reg [31:0] _RAND_65;
  reg [31:0] _T_1140; // @[Reg.scala 11:16:@464.4]
  reg [31:0] _RAND_66;
  reg [31:0] _T_1142; // @[Reg.scala 11:16:@468.4]
  reg [31:0] _RAND_67;
  reg [31:0] _T_1144; // @[Reg.scala 11:16:@472.4]
  reg [31:0] _RAND_68;
  reg [31:0] _T_1146; // @[Reg.scala 11:16:@476.4]
  reg [31:0] _RAND_69;
  reg [31:0] _T_1149; // @[Reg.scala 11:16:@480.4]
  reg [31:0] _RAND_70;
  reg [31:0] _T_1151; // @[Reg.scala 11:16:@484.4]
  reg [31:0] _RAND_71;
  reg [31:0] _T_1153; // @[Reg.scala 11:16:@488.4]
  reg [31:0] _RAND_72;
  reg [31:0] _T_1155; // @[Reg.scala 11:16:@492.4]
  reg [31:0] _RAND_73;
  reg [31:0] _T_1157; // @[Reg.scala 11:16:@496.4]
  reg [31:0] _RAND_74;
  reg [31:0] _T_1160; // @[Reg.scala 11:16:@500.4]
  reg [31:0] _RAND_75;
  reg [31:0] _T_1162; // @[Reg.scala 11:16:@504.4]
  reg [31:0] _RAND_76;
  reg [31:0] _T_1164; // @[Reg.scala 11:16:@508.4]
  reg [31:0] _RAND_77;
  reg [31:0] _T_1166; // @[Reg.scala 11:16:@512.4]
  reg [31:0] _RAND_78;
  reg [31:0] _T_1168; // @[Reg.scala 11:16:@516.4]
  reg [31:0] _RAND_79;
  assign _T_724 = io_inputs_0 + io_inputs_0; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 32:53:@8.4]
  assign _T_725 = io_inputs_0 + io_inputs_0; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 32:53:@9.4]
  assign _T_727 = io_inputs_0 * io_inputs_0; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 33:58:@10.4]
  assign _T_729 = io_inputs_0 / io_inputs_0; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 34:56:@11.4]
  assign _T_730 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_731 = _T_730 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_732 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_733 = _T_732 ? _T_727 : {{16'd0}, _T_731}; // @[Mux.scala 46:16:@15.4]
  assign _T_734 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_735 = _T_734 ? {{16'd0}, _T_725} : _T_733; // @[Mux.scala 46:16:@17.4]
  assign _T_736 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _T_747 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_748 = _T_747 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_749 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_750 = _T_749 ? _T_727 : {{16'd0}, _T_748}; // @[Mux.scala 46:16:@27.4]
  assign _T_751 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_752 = _T_751 ? {{16'd0}, _T_725} : _T_750; // @[Mux.scala 46:16:@29.4]
  assign _T_753 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _T_764 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_765 = _T_764 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_766 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_767 = _T_766 ? _T_727 : {{16'd0}, _T_765}; // @[Mux.scala 46:16:@39.4]
  assign _T_768 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_769 = _T_768 ? {{16'd0}, _T_725} : _T_767; // @[Mux.scala 46:16:@41.4]
  assign _T_770 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _T_781 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_782 = _T_781 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_783 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_784 = _T_783 ? _T_727 : {{16'd0}, _T_782}; // @[Mux.scala 46:16:@51.4]
  assign _T_785 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_786 = _T_785 ? {{16'd0}, _T_725} : _T_784; // @[Mux.scala 46:16:@53.4]
  assign _T_787 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _T_798 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_799 = _T_798 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_800 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_801 = _T_800 ? _T_727 : {{16'd0}, _T_799}; // @[Mux.scala 46:16:@63.4]
  assign _T_802 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_803 = _T_802 ? {{16'd0}, _T_725} : _T_801; // @[Mux.scala 46:16:@65.4]
  assign _T_804 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _T_815 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_816 = _T_815 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_817 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_818 = _T_817 ? _T_727 : {{16'd0}, _T_816}; // @[Mux.scala 46:16:@75.4]
  assign _T_819 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_820 = _T_819 ? {{16'd0}, _T_725} : _T_818; // @[Mux.scala 46:16:@77.4]
  assign _T_821 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _T_832 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_833 = _T_832 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_834 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_835 = _T_834 ? _T_727 : {{16'd0}, _T_833}; // @[Mux.scala 46:16:@87.4]
  assign _T_836 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_837 = _T_836 ? {{16'd0}, _T_725} : _T_835; // @[Mux.scala 46:16:@89.4]
  assign _T_838 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _T_849 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_850 = _T_849 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_851 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_852 = _T_851 ? _T_727 : {{16'd0}, _T_850}; // @[Mux.scala 46:16:@99.4]
  assign _T_853 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_854 = _T_853 ? {{16'd0}, _T_725} : _T_852; // @[Mux.scala 46:16:@101.4]
  assign _T_855 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign _T_866 = 3'h3 == io_operation_8; // @[Mux.scala 46:19:@108.4]
  assign _T_867 = _T_866 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@109.4]
  assign _T_868 = 3'h2 == io_operation_8; // @[Mux.scala 46:19:@110.4]
  assign _T_869 = _T_868 ? _T_727 : {{16'd0}, _T_867}; // @[Mux.scala 46:16:@111.4]
  assign _T_870 = 3'h1 == io_operation_8; // @[Mux.scala 46:19:@112.4]
  assign _T_871 = _T_870 ? {{16'd0}, _T_725} : _T_869; // @[Mux.scala 46:16:@113.4]
  assign _T_872 = 3'h0 == io_operation_8; // @[Mux.scala 46:19:@114.4]
  assign _T_883 = 3'h3 == io_operation_9; // @[Mux.scala 46:19:@120.4]
  assign _T_884 = _T_883 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@121.4]
  assign _T_885 = 3'h2 == io_operation_9; // @[Mux.scala 46:19:@122.4]
  assign _T_886 = _T_885 ? _T_727 : {{16'd0}, _T_884}; // @[Mux.scala 46:16:@123.4]
  assign _T_887 = 3'h1 == io_operation_9; // @[Mux.scala 46:19:@124.4]
  assign _T_888 = _T_887 ? {{16'd0}, _T_725} : _T_886; // @[Mux.scala 46:16:@125.4]
  assign _T_889 = 3'h0 == io_operation_9; // @[Mux.scala 46:19:@126.4]
  assign _T_900 = 3'h3 == io_operation_10; // @[Mux.scala 46:19:@132.4]
  assign _T_901 = _T_900 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@133.4]
  assign _T_902 = 3'h2 == io_operation_10; // @[Mux.scala 46:19:@134.4]
  assign _T_903 = _T_902 ? _T_727 : {{16'd0}, _T_901}; // @[Mux.scala 46:16:@135.4]
  assign _T_904 = 3'h1 == io_operation_10; // @[Mux.scala 46:19:@136.4]
  assign _T_905 = _T_904 ? {{16'd0}, _T_725} : _T_903; // @[Mux.scala 46:16:@137.4]
  assign _T_906 = 3'h0 == io_operation_10; // @[Mux.scala 46:19:@138.4]
  assign _T_917 = 3'h3 == io_operation_11; // @[Mux.scala 46:19:@144.4]
  assign _T_918 = _T_917 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@145.4]
  assign _T_919 = 3'h2 == io_operation_11; // @[Mux.scala 46:19:@146.4]
  assign _T_920 = _T_919 ? _T_727 : {{16'd0}, _T_918}; // @[Mux.scala 46:16:@147.4]
  assign _T_921 = 3'h1 == io_operation_11; // @[Mux.scala 46:19:@148.4]
  assign _T_922 = _T_921 ? {{16'd0}, _T_725} : _T_920; // @[Mux.scala 46:16:@149.4]
  assign _T_923 = 3'h0 == io_operation_11; // @[Mux.scala 46:19:@150.4]
  assign _T_934 = 3'h3 == io_operation_12; // @[Mux.scala 46:19:@156.4]
  assign _T_935 = _T_934 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@157.4]
  assign _T_936 = 3'h2 == io_operation_12; // @[Mux.scala 46:19:@158.4]
  assign _T_937 = _T_936 ? _T_727 : {{16'd0}, _T_935}; // @[Mux.scala 46:16:@159.4]
  assign _T_938 = 3'h1 == io_operation_12; // @[Mux.scala 46:19:@160.4]
  assign _T_939 = _T_938 ? {{16'd0}, _T_725} : _T_937; // @[Mux.scala 46:16:@161.4]
  assign _T_940 = 3'h0 == io_operation_12; // @[Mux.scala 46:19:@162.4]
  assign _T_951 = 3'h3 == io_operation_13; // @[Mux.scala 46:19:@168.4]
  assign _T_952 = _T_951 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@169.4]
  assign _T_953 = 3'h2 == io_operation_13; // @[Mux.scala 46:19:@170.4]
  assign _T_954 = _T_953 ? _T_727 : {{16'd0}, _T_952}; // @[Mux.scala 46:16:@171.4]
  assign _T_955 = 3'h1 == io_operation_13; // @[Mux.scala 46:19:@172.4]
  assign _T_956 = _T_955 ? {{16'd0}, _T_725} : _T_954; // @[Mux.scala 46:16:@173.4]
  assign _T_957 = 3'h0 == io_operation_13; // @[Mux.scala 46:19:@174.4]
  assign _T_968 = 3'h3 == io_operation_14; // @[Mux.scala 46:19:@180.4]
  assign _T_969 = _T_968 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@181.4]
  assign _T_970 = 3'h2 == io_operation_14; // @[Mux.scala 46:19:@182.4]
  assign _T_971 = _T_970 ? _T_727 : {{16'd0}, _T_969}; // @[Mux.scala 46:16:@183.4]
  assign _T_972 = 3'h1 == io_operation_14; // @[Mux.scala 46:19:@184.4]
  assign _T_973 = _T_972 ? {{16'd0}, _T_725} : _T_971; // @[Mux.scala 46:16:@185.4]
  assign _T_974 = 3'h0 == io_operation_14; // @[Mux.scala 46:19:@186.4]
  assign _T_985 = 3'h3 == io_operation_15; // @[Mux.scala 46:19:@192.4]
  assign _T_986 = _T_985 ? _T_729 : 16'h0; // @[Mux.scala 46:16:@193.4]
  assign _T_987 = 3'h2 == io_operation_15; // @[Mux.scala 46:19:@194.4]
  assign _T_988 = _T_987 ? _T_727 : {{16'd0}, _T_986}; // @[Mux.scala 46:16:@195.4]
  assign _T_989 = 3'h1 == io_operation_15; // @[Mux.scala 46:19:@196.4]
  assign _T_990 = _T_989 ? {{16'd0}, _T_725} : _T_988; // @[Mux.scala 46:16:@197.4]
  assign _T_991 = 3'h0 == io_operation_15; // @[Mux.scala 46:19:@198.4]
  assign io_outputs_0 = _T_1003[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@520.4]
  assign io_outputs_1 = _T_1014[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@521.4]
  assign io_outputs_2 = _T_1025[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@522.4]
  assign io_outputs_3 = _T_1036[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@523.4]
  assign io_outputs_4 = _T_1047[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@524.4]
  assign io_outputs_5 = _T_1058[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@525.4]
  assign io_outputs_6 = _T_1069[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@526.4]
  assign io_outputs_7 = _T_1080[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@527.4]
  assign io_outputs_8 = _T_1091[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@528.4]
  assign io_outputs_9 = _T_1102[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@529.4]
  assign io_outputs_10 = _T_1113[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@530.4]
  assign io_outputs_11 = _T_1124[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@531.4]
  assign io_outputs_12 = _T_1135[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@532.4]
  assign io_outputs_13 = _T_1146[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@533.4]
  assign io_outputs_14 = _T_1157[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@534.4]
  assign io_outputs_15 = _T_1168[15:0]; // @[MuxTest_width_16_inputs_1_outputs_16_pipeline_5s.scala 23:14:@535.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_995 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_997 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_999 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_1001 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_1003 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_1006 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1008 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1010 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_1012 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_1014 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_1017 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_1019 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_1021 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_1023 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_1025 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_1028 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1030 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_1032 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_1034 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_1036 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_1039 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_1041 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_1043 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_1045 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_1047 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_1050 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_1052 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_1054 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_1056 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_1058 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_1061 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_1063 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_1065 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_1067 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_1069 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_1072 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_1074 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_1076 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_1078 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_1080 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_1083 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_1085 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_1087 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_1089 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_1091 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_1094 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_1096 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_1098 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_1100 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_1102 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_1105 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1107 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_1109 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_1111 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_1113 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_1116 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_1118 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_1120 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_1122 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_1124 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_1127 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_1129 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_1131 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_1133 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_1135 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_1138 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_1140 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_1142 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_1144 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_1146 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_1149 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_1151 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1153 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1155 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1157 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1160 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_1162 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1164 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_1166 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_1168 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_736) begin
      _T_995 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_995 <= _T_735;
    end
    _T_997 <= _T_995;
    _T_999 <= _T_997;
    _T_1001 <= _T_999;
    _T_1003 <= _T_1001;
    if (_T_753) begin
      _T_1006 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1006 <= _T_752;
    end
    _T_1008 <= _T_1006;
    _T_1010 <= _T_1008;
    _T_1012 <= _T_1010;
    _T_1014 <= _T_1012;
    if (_T_770) begin
      _T_1017 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1017 <= _T_769;
    end
    _T_1019 <= _T_1017;
    _T_1021 <= _T_1019;
    _T_1023 <= _T_1021;
    _T_1025 <= _T_1023;
    if (_T_787) begin
      _T_1028 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1028 <= _T_786;
    end
    _T_1030 <= _T_1028;
    _T_1032 <= _T_1030;
    _T_1034 <= _T_1032;
    _T_1036 <= _T_1034;
    if (_T_804) begin
      _T_1039 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1039 <= _T_803;
    end
    _T_1041 <= _T_1039;
    _T_1043 <= _T_1041;
    _T_1045 <= _T_1043;
    _T_1047 <= _T_1045;
    if (_T_821) begin
      _T_1050 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1050 <= _T_820;
    end
    _T_1052 <= _T_1050;
    _T_1054 <= _T_1052;
    _T_1056 <= _T_1054;
    _T_1058 <= _T_1056;
    if (_T_838) begin
      _T_1061 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1061 <= _T_837;
    end
    _T_1063 <= _T_1061;
    _T_1065 <= _T_1063;
    _T_1067 <= _T_1065;
    _T_1069 <= _T_1067;
    if (_T_855) begin
      _T_1072 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1072 <= _T_854;
    end
    _T_1074 <= _T_1072;
    _T_1076 <= _T_1074;
    _T_1078 <= _T_1076;
    _T_1080 <= _T_1078;
    if (_T_872) begin
      _T_1083 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1083 <= _T_871;
    end
    _T_1085 <= _T_1083;
    _T_1087 <= _T_1085;
    _T_1089 <= _T_1087;
    _T_1091 <= _T_1089;
    if (_T_889) begin
      _T_1094 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1094 <= _T_888;
    end
    _T_1096 <= _T_1094;
    _T_1098 <= _T_1096;
    _T_1100 <= _T_1098;
    _T_1102 <= _T_1100;
    if (_T_906) begin
      _T_1105 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1105 <= _T_905;
    end
    _T_1107 <= _T_1105;
    _T_1109 <= _T_1107;
    _T_1111 <= _T_1109;
    _T_1113 <= _T_1111;
    if (_T_923) begin
      _T_1116 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1116 <= _T_922;
    end
    _T_1118 <= _T_1116;
    _T_1120 <= _T_1118;
    _T_1122 <= _T_1120;
    _T_1124 <= _T_1122;
    if (_T_940) begin
      _T_1127 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1127 <= _T_939;
    end
    _T_1129 <= _T_1127;
    _T_1131 <= _T_1129;
    _T_1133 <= _T_1131;
    _T_1135 <= _T_1133;
    if (_T_957) begin
      _T_1138 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1138 <= _T_956;
    end
    _T_1140 <= _T_1138;
    _T_1142 <= _T_1140;
    _T_1144 <= _T_1142;
    _T_1146 <= _T_1144;
    if (_T_974) begin
      _T_1149 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1149 <= _T_973;
    end
    _T_1151 <= _T_1149;
    _T_1153 <= _T_1151;
    _T_1155 <= _T_1153;
    _T_1157 <= _T_1155;
    if (_T_991) begin
      _T_1160 <= {{16'd0}, io_inputs_0};
    end else begin
      _T_1160 <= _T_990;
    end
    _T_1162 <= _T_1160;
    _T_1164 <= _T_1162;
    _T_1166 <= _T_1164;
    _T_1168 <= _T_1166;
  end
endmodule
