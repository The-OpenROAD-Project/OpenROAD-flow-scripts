VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram7_2048x39
  FOREIGN fakeram7_2048x39 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 5.130 BY 532.000 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.048 0.024 0.072 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.808 0.024 5.832 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.568 0.024 11.592 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 17.328 0.024 17.352 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 23.088 0.024 23.112 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 28.848 0.024 28.872 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 34.608 0.024 34.632 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 40.368 0.024 40.392 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 46.128 0.024 46.152 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 51.888 0.024 51.912 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 57.648 0.024 57.672 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 63.408 0.024 63.432 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 69.168 0.024 69.192 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 74.928 0.024 74.952 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 80.688 0.024 80.712 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 86.448 0.024 86.472 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 92.208 0.024 92.232 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 97.968 0.024 97.992 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 103.728 0.024 103.752 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 109.488 0.024 109.512 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 115.248 0.024 115.272 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 121.008 0.024 121.032 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 126.768 0.024 126.792 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 132.528 0.024 132.552 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 138.288 0.024 138.312 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 144.048 0.024 144.072 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 149.808 0.024 149.832 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 155.568 0.024 155.592 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 161.328 0.024 161.352 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 167.088 0.024 167.112 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 172.848 0.024 172.872 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 178.608 0.024 178.632 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 184.368 0.024 184.392 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 190.128 0.024 190.152 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 195.888 0.024 195.912 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 201.648 0.024 201.672 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 207.408 0.024 207.432 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 213.168 0.024 213.192 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 218.928 0.024 218.952 ;
    END
  END rd_out[38]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 219.408 0.024 219.432 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 225.168 0.024 225.192 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 230.928 0.024 230.952 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 236.688 0.024 236.712 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 242.448 0.024 242.472 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 248.208 0.024 248.232 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 253.968 0.024 253.992 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 259.728 0.024 259.752 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 265.488 0.024 265.512 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 271.248 0.024 271.272 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 277.008 0.024 277.032 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 282.768 0.024 282.792 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 288.528 0.024 288.552 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 294.288 0.024 294.312 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 300.048 0.024 300.072 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 305.808 0.024 305.832 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 311.568 0.024 311.592 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 317.328 0.024 317.352 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 323.088 0.024 323.112 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 328.848 0.024 328.872 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 334.608 0.024 334.632 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 340.368 0.024 340.392 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 346.128 0.024 346.152 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 351.888 0.024 351.912 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 357.648 0.024 357.672 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 363.408 0.024 363.432 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 369.168 0.024 369.192 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 374.928 0.024 374.952 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 380.688 0.024 380.712 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 386.448 0.024 386.472 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 392.208 0.024 392.232 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 397.968 0.024 397.992 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 403.728 0.024 403.752 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 409.488 0.024 409.512 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 415.248 0.024 415.272 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 421.008 0.024 421.032 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 426.768 0.024 426.792 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 432.528 0.024 432.552 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 438.288 0.024 438.312 ;
    END
  END wd_in[38]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 438.768 0.024 438.792 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 444.528 0.024 444.552 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 450.288 0.024 450.312 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 456.048 0.024 456.072 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 461.808 0.024 461.832 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 467.568 0.024 467.592 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 473.328 0.024 473.352 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 479.088 0.024 479.112 ;
    END
  END addr_in[7]
  PIN addr_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 484.848 0.024 484.872 ;
    END
  END addr_in[8]
  PIN addr_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 490.608 0.024 490.632 ;
    END
  END addr_in[9]
  PIN addr_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 496.368 0.024 496.392 ;
    END
  END addr_in[10]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 496.848 0.024 496.872 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 502.608 0.024 502.632 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 508.368 0.024 508.392 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.000 5.082 0.096 ;
      RECT 0.048 0.768 5.082 0.864 ;
      RECT 0.048 1.536 5.082 1.632 ;
      RECT 0.048 2.304 5.082 2.400 ;
      RECT 0.048 3.072 5.082 3.168 ;
      RECT 0.048 3.840 5.082 3.936 ;
      RECT 0.048 4.608 5.082 4.704 ;
      RECT 0.048 5.376 5.082 5.472 ;
      RECT 0.048 6.144 5.082 6.240 ;
      RECT 0.048 6.912 5.082 7.008 ;
      RECT 0.048 7.680 5.082 7.776 ;
      RECT 0.048 8.448 5.082 8.544 ;
      RECT 0.048 9.216 5.082 9.312 ;
      RECT 0.048 9.984 5.082 10.080 ;
      RECT 0.048 10.752 5.082 10.848 ;
      RECT 0.048 11.520 5.082 11.616 ;
      RECT 0.048 12.288 5.082 12.384 ;
      RECT 0.048 13.056 5.082 13.152 ;
      RECT 0.048 13.824 5.082 13.920 ;
      RECT 0.048 14.592 5.082 14.688 ;
      RECT 0.048 15.360 5.082 15.456 ;
      RECT 0.048 16.128 5.082 16.224 ;
      RECT 0.048 16.896 5.082 16.992 ;
      RECT 0.048 17.664 5.082 17.760 ;
      RECT 0.048 18.432 5.082 18.528 ;
      RECT 0.048 19.200 5.082 19.296 ;
      RECT 0.048 19.968 5.082 20.064 ;
      RECT 0.048 20.736 5.082 20.832 ;
      RECT 0.048 21.504 5.082 21.600 ;
      RECT 0.048 22.272 5.082 22.368 ;
      RECT 0.048 23.040 5.082 23.136 ;
      RECT 0.048 23.808 5.082 23.904 ;
      RECT 0.048 24.576 5.082 24.672 ;
      RECT 0.048 25.344 5.082 25.440 ;
      RECT 0.048 26.112 5.082 26.208 ;
      RECT 0.048 26.880 5.082 26.976 ;
      RECT 0.048 27.648 5.082 27.744 ;
      RECT 0.048 28.416 5.082 28.512 ;
      RECT 0.048 29.184 5.082 29.280 ;
      RECT 0.048 29.952 5.082 30.048 ;
      RECT 0.048 30.720 5.082 30.816 ;
      RECT 0.048 31.488 5.082 31.584 ;
      RECT 0.048 32.256 5.082 32.352 ;
      RECT 0.048 33.024 5.082 33.120 ;
      RECT 0.048 33.792 5.082 33.888 ;
      RECT 0.048 34.560 5.082 34.656 ;
      RECT 0.048 35.328 5.082 35.424 ;
      RECT 0.048 36.096 5.082 36.192 ;
      RECT 0.048 36.864 5.082 36.960 ;
      RECT 0.048 37.632 5.082 37.728 ;
      RECT 0.048 38.400 5.082 38.496 ;
      RECT 0.048 39.168 5.082 39.264 ;
      RECT 0.048 39.936 5.082 40.032 ;
      RECT 0.048 40.704 5.082 40.800 ;
      RECT 0.048 41.472 5.082 41.568 ;
      RECT 0.048 42.240 5.082 42.336 ;
      RECT 0.048 43.008 5.082 43.104 ;
      RECT 0.048 43.776 5.082 43.872 ;
      RECT 0.048 44.544 5.082 44.640 ;
      RECT 0.048 45.312 5.082 45.408 ;
      RECT 0.048 46.080 5.082 46.176 ;
      RECT 0.048 46.848 5.082 46.944 ;
      RECT 0.048 47.616 5.082 47.712 ;
      RECT 0.048 48.384 5.082 48.480 ;
      RECT 0.048 49.152 5.082 49.248 ;
      RECT 0.048 49.920 5.082 50.016 ;
      RECT 0.048 50.688 5.082 50.784 ;
      RECT 0.048 51.456 5.082 51.552 ;
      RECT 0.048 52.224 5.082 52.320 ;
      RECT 0.048 52.992 5.082 53.088 ;
      RECT 0.048 53.760 5.082 53.856 ;
      RECT 0.048 54.528 5.082 54.624 ;
      RECT 0.048 55.296 5.082 55.392 ;
      RECT 0.048 56.064 5.082 56.160 ;
      RECT 0.048 56.832 5.082 56.928 ;
      RECT 0.048 57.600 5.082 57.696 ;
      RECT 0.048 58.368 5.082 58.464 ;
      RECT 0.048 59.136 5.082 59.232 ;
      RECT 0.048 59.904 5.082 60.000 ;
      RECT 0.048 60.672 5.082 60.768 ;
      RECT 0.048 61.440 5.082 61.536 ;
      RECT 0.048 62.208 5.082 62.304 ;
      RECT 0.048 62.976 5.082 63.072 ;
      RECT 0.048 63.744 5.082 63.840 ;
      RECT 0.048 64.512 5.082 64.608 ;
      RECT 0.048 65.280 5.082 65.376 ;
      RECT 0.048 66.048 5.082 66.144 ;
      RECT 0.048 66.816 5.082 66.912 ;
      RECT 0.048 67.584 5.082 67.680 ;
      RECT 0.048 68.352 5.082 68.448 ;
      RECT 0.048 69.120 5.082 69.216 ;
      RECT 0.048 69.888 5.082 69.984 ;
      RECT 0.048 70.656 5.082 70.752 ;
      RECT 0.048 71.424 5.082 71.520 ;
      RECT 0.048 72.192 5.082 72.288 ;
      RECT 0.048 72.960 5.082 73.056 ;
      RECT 0.048 73.728 5.082 73.824 ;
      RECT 0.048 74.496 5.082 74.592 ;
      RECT 0.048 75.264 5.082 75.360 ;
      RECT 0.048 76.032 5.082 76.128 ;
      RECT 0.048 76.800 5.082 76.896 ;
      RECT 0.048 77.568 5.082 77.664 ;
      RECT 0.048 78.336 5.082 78.432 ;
      RECT 0.048 79.104 5.082 79.200 ;
      RECT 0.048 79.872 5.082 79.968 ;
      RECT 0.048 80.640 5.082 80.736 ;
      RECT 0.048 81.408 5.082 81.504 ;
      RECT 0.048 82.176 5.082 82.272 ;
      RECT 0.048 82.944 5.082 83.040 ;
      RECT 0.048 83.712 5.082 83.808 ;
      RECT 0.048 84.480 5.082 84.576 ;
      RECT 0.048 85.248 5.082 85.344 ;
      RECT 0.048 86.016 5.082 86.112 ;
      RECT 0.048 86.784 5.082 86.880 ;
      RECT 0.048 87.552 5.082 87.648 ;
      RECT 0.048 88.320 5.082 88.416 ;
      RECT 0.048 89.088 5.082 89.184 ;
      RECT 0.048 89.856 5.082 89.952 ;
      RECT 0.048 90.624 5.082 90.720 ;
      RECT 0.048 91.392 5.082 91.488 ;
      RECT 0.048 92.160 5.082 92.256 ;
      RECT 0.048 92.928 5.082 93.024 ;
      RECT 0.048 93.696 5.082 93.792 ;
      RECT 0.048 94.464 5.082 94.560 ;
      RECT 0.048 95.232 5.082 95.328 ;
      RECT 0.048 96.000 5.082 96.096 ;
      RECT 0.048 96.768 5.082 96.864 ;
      RECT 0.048 97.536 5.082 97.632 ;
      RECT 0.048 98.304 5.082 98.400 ;
      RECT 0.048 99.072 5.082 99.168 ;
      RECT 0.048 99.840 5.082 99.936 ;
      RECT 0.048 100.608 5.082 100.704 ;
      RECT 0.048 101.376 5.082 101.472 ;
      RECT 0.048 102.144 5.082 102.240 ;
      RECT 0.048 102.912 5.082 103.008 ;
      RECT 0.048 103.680 5.082 103.776 ;
      RECT 0.048 104.448 5.082 104.544 ;
      RECT 0.048 105.216 5.082 105.312 ;
      RECT 0.048 105.984 5.082 106.080 ;
      RECT 0.048 106.752 5.082 106.848 ;
      RECT 0.048 107.520 5.082 107.616 ;
      RECT 0.048 108.288 5.082 108.384 ;
      RECT 0.048 109.056 5.082 109.152 ;
      RECT 0.048 109.824 5.082 109.920 ;
      RECT 0.048 110.592 5.082 110.688 ;
      RECT 0.048 111.360 5.082 111.456 ;
      RECT 0.048 112.128 5.082 112.224 ;
      RECT 0.048 112.896 5.082 112.992 ;
      RECT 0.048 113.664 5.082 113.760 ;
      RECT 0.048 114.432 5.082 114.528 ;
      RECT 0.048 115.200 5.082 115.296 ;
      RECT 0.048 115.968 5.082 116.064 ;
      RECT 0.048 116.736 5.082 116.832 ;
      RECT 0.048 117.504 5.082 117.600 ;
      RECT 0.048 118.272 5.082 118.368 ;
      RECT 0.048 119.040 5.082 119.136 ;
      RECT 0.048 119.808 5.082 119.904 ;
      RECT 0.048 120.576 5.082 120.672 ;
      RECT 0.048 121.344 5.082 121.440 ;
      RECT 0.048 122.112 5.082 122.208 ;
      RECT 0.048 122.880 5.082 122.976 ;
      RECT 0.048 123.648 5.082 123.744 ;
      RECT 0.048 124.416 5.082 124.512 ;
      RECT 0.048 125.184 5.082 125.280 ;
      RECT 0.048 125.952 5.082 126.048 ;
      RECT 0.048 126.720 5.082 126.816 ;
      RECT 0.048 127.488 5.082 127.584 ;
      RECT 0.048 128.256 5.082 128.352 ;
      RECT 0.048 129.024 5.082 129.120 ;
      RECT 0.048 129.792 5.082 129.888 ;
      RECT 0.048 130.560 5.082 130.656 ;
      RECT 0.048 131.328 5.082 131.424 ;
      RECT 0.048 132.096 5.082 132.192 ;
      RECT 0.048 132.864 5.082 132.960 ;
      RECT 0.048 133.632 5.082 133.728 ;
      RECT 0.048 134.400 5.082 134.496 ;
      RECT 0.048 135.168 5.082 135.264 ;
      RECT 0.048 135.936 5.082 136.032 ;
      RECT 0.048 136.704 5.082 136.800 ;
      RECT 0.048 137.472 5.082 137.568 ;
      RECT 0.048 138.240 5.082 138.336 ;
      RECT 0.048 139.008 5.082 139.104 ;
      RECT 0.048 139.776 5.082 139.872 ;
      RECT 0.048 140.544 5.082 140.640 ;
      RECT 0.048 141.312 5.082 141.408 ;
      RECT 0.048 142.080 5.082 142.176 ;
      RECT 0.048 142.848 5.082 142.944 ;
      RECT 0.048 143.616 5.082 143.712 ;
      RECT 0.048 144.384 5.082 144.480 ;
      RECT 0.048 145.152 5.082 145.248 ;
      RECT 0.048 145.920 5.082 146.016 ;
      RECT 0.048 146.688 5.082 146.784 ;
      RECT 0.048 147.456 5.082 147.552 ;
      RECT 0.048 148.224 5.082 148.320 ;
      RECT 0.048 148.992 5.082 149.088 ;
      RECT 0.048 149.760 5.082 149.856 ;
      RECT 0.048 150.528 5.082 150.624 ;
      RECT 0.048 151.296 5.082 151.392 ;
      RECT 0.048 152.064 5.082 152.160 ;
      RECT 0.048 152.832 5.082 152.928 ;
      RECT 0.048 153.600 5.082 153.696 ;
      RECT 0.048 154.368 5.082 154.464 ;
      RECT 0.048 155.136 5.082 155.232 ;
      RECT 0.048 155.904 5.082 156.000 ;
      RECT 0.048 156.672 5.082 156.768 ;
      RECT 0.048 157.440 5.082 157.536 ;
      RECT 0.048 158.208 5.082 158.304 ;
      RECT 0.048 158.976 5.082 159.072 ;
      RECT 0.048 159.744 5.082 159.840 ;
      RECT 0.048 160.512 5.082 160.608 ;
      RECT 0.048 161.280 5.082 161.376 ;
      RECT 0.048 162.048 5.082 162.144 ;
      RECT 0.048 162.816 5.082 162.912 ;
      RECT 0.048 163.584 5.082 163.680 ;
      RECT 0.048 164.352 5.082 164.448 ;
      RECT 0.048 165.120 5.082 165.216 ;
      RECT 0.048 165.888 5.082 165.984 ;
      RECT 0.048 166.656 5.082 166.752 ;
      RECT 0.048 167.424 5.082 167.520 ;
      RECT 0.048 168.192 5.082 168.288 ;
      RECT 0.048 168.960 5.082 169.056 ;
      RECT 0.048 169.728 5.082 169.824 ;
      RECT 0.048 170.496 5.082 170.592 ;
      RECT 0.048 171.264 5.082 171.360 ;
      RECT 0.048 172.032 5.082 172.128 ;
      RECT 0.048 172.800 5.082 172.896 ;
      RECT 0.048 173.568 5.082 173.664 ;
      RECT 0.048 174.336 5.082 174.432 ;
      RECT 0.048 175.104 5.082 175.200 ;
      RECT 0.048 175.872 5.082 175.968 ;
      RECT 0.048 176.640 5.082 176.736 ;
      RECT 0.048 177.408 5.082 177.504 ;
      RECT 0.048 178.176 5.082 178.272 ;
      RECT 0.048 178.944 5.082 179.040 ;
      RECT 0.048 179.712 5.082 179.808 ;
      RECT 0.048 180.480 5.082 180.576 ;
      RECT 0.048 181.248 5.082 181.344 ;
      RECT 0.048 182.016 5.082 182.112 ;
      RECT 0.048 182.784 5.082 182.880 ;
      RECT 0.048 183.552 5.082 183.648 ;
      RECT 0.048 184.320 5.082 184.416 ;
      RECT 0.048 185.088 5.082 185.184 ;
      RECT 0.048 185.856 5.082 185.952 ;
      RECT 0.048 186.624 5.082 186.720 ;
      RECT 0.048 187.392 5.082 187.488 ;
      RECT 0.048 188.160 5.082 188.256 ;
      RECT 0.048 188.928 5.082 189.024 ;
      RECT 0.048 189.696 5.082 189.792 ;
      RECT 0.048 190.464 5.082 190.560 ;
      RECT 0.048 191.232 5.082 191.328 ;
      RECT 0.048 192.000 5.082 192.096 ;
      RECT 0.048 192.768 5.082 192.864 ;
      RECT 0.048 193.536 5.082 193.632 ;
      RECT 0.048 194.304 5.082 194.400 ;
      RECT 0.048 195.072 5.082 195.168 ;
      RECT 0.048 195.840 5.082 195.936 ;
      RECT 0.048 196.608 5.082 196.704 ;
      RECT 0.048 197.376 5.082 197.472 ;
      RECT 0.048 198.144 5.082 198.240 ;
      RECT 0.048 198.912 5.082 199.008 ;
      RECT 0.048 199.680 5.082 199.776 ;
      RECT 0.048 200.448 5.082 200.544 ;
      RECT 0.048 201.216 5.082 201.312 ;
      RECT 0.048 201.984 5.082 202.080 ;
      RECT 0.048 202.752 5.082 202.848 ;
      RECT 0.048 203.520 5.082 203.616 ;
      RECT 0.048 204.288 5.082 204.384 ;
      RECT 0.048 205.056 5.082 205.152 ;
      RECT 0.048 205.824 5.082 205.920 ;
      RECT 0.048 206.592 5.082 206.688 ;
      RECT 0.048 207.360 5.082 207.456 ;
      RECT 0.048 208.128 5.082 208.224 ;
      RECT 0.048 208.896 5.082 208.992 ;
      RECT 0.048 209.664 5.082 209.760 ;
      RECT 0.048 210.432 5.082 210.528 ;
      RECT 0.048 211.200 5.082 211.296 ;
      RECT 0.048 211.968 5.082 212.064 ;
      RECT 0.048 212.736 5.082 212.832 ;
      RECT 0.048 213.504 5.082 213.600 ;
      RECT 0.048 214.272 5.082 214.368 ;
      RECT 0.048 215.040 5.082 215.136 ;
      RECT 0.048 215.808 5.082 215.904 ;
      RECT 0.048 216.576 5.082 216.672 ;
      RECT 0.048 217.344 5.082 217.440 ;
      RECT 0.048 218.112 5.082 218.208 ;
      RECT 0.048 218.880 5.082 218.976 ;
      RECT 0.048 219.648 5.082 219.744 ;
      RECT 0.048 220.416 5.082 220.512 ;
      RECT 0.048 221.184 5.082 221.280 ;
      RECT 0.048 221.952 5.082 222.048 ;
      RECT 0.048 222.720 5.082 222.816 ;
      RECT 0.048 223.488 5.082 223.584 ;
      RECT 0.048 224.256 5.082 224.352 ;
      RECT 0.048 225.024 5.082 225.120 ;
      RECT 0.048 225.792 5.082 225.888 ;
      RECT 0.048 226.560 5.082 226.656 ;
      RECT 0.048 227.328 5.082 227.424 ;
      RECT 0.048 228.096 5.082 228.192 ;
      RECT 0.048 228.864 5.082 228.960 ;
      RECT 0.048 229.632 5.082 229.728 ;
      RECT 0.048 230.400 5.082 230.496 ;
      RECT 0.048 231.168 5.082 231.264 ;
      RECT 0.048 231.936 5.082 232.032 ;
      RECT 0.048 232.704 5.082 232.800 ;
      RECT 0.048 233.472 5.082 233.568 ;
      RECT 0.048 234.240 5.082 234.336 ;
      RECT 0.048 235.008 5.082 235.104 ;
      RECT 0.048 235.776 5.082 235.872 ;
      RECT 0.048 236.544 5.082 236.640 ;
      RECT 0.048 237.312 5.082 237.408 ;
      RECT 0.048 238.080 5.082 238.176 ;
      RECT 0.048 238.848 5.082 238.944 ;
      RECT 0.048 239.616 5.082 239.712 ;
      RECT 0.048 240.384 5.082 240.480 ;
      RECT 0.048 241.152 5.082 241.248 ;
      RECT 0.048 241.920 5.082 242.016 ;
      RECT 0.048 242.688 5.082 242.784 ;
      RECT 0.048 243.456 5.082 243.552 ;
      RECT 0.048 244.224 5.082 244.320 ;
      RECT 0.048 244.992 5.082 245.088 ;
      RECT 0.048 245.760 5.082 245.856 ;
      RECT 0.048 246.528 5.082 246.624 ;
      RECT 0.048 247.296 5.082 247.392 ;
      RECT 0.048 248.064 5.082 248.160 ;
      RECT 0.048 248.832 5.082 248.928 ;
      RECT 0.048 249.600 5.082 249.696 ;
      RECT 0.048 250.368 5.082 250.464 ;
      RECT 0.048 251.136 5.082 251.232 ;
      RECT 0.048 251.904 5.082 252.000 ;
      RECT 0.048 252.672 5.082 252.768 ;
      RECT 0.048 253.440 5.082 253.536 ;
      RECT 0.048 254.208 5.082 254.304 ;
      RECT 0.048 254.976 5.082 255.072 ;
      RECT 0.048 255.744 5.082 255.840 ;
      RECT 0.048 256.512 5.082 256.608 ;
      RECT 0.048 257.280 5.082 257.376 ;
      RECT 0.048 258.048 5.082 258.144 ;
      RECT 0.048 258.816 5.082 258.912 ;
      RECT 0.048 259.584 5.082 259.680 ;
      RECT 0.048 260.352 5.082 260.448 ;
      RECT 0.048 261.120 5.082 261.216 ;
      RECT 0.048 261.888 5.082 261.984 ;
      RECT 0.048 262.656 5.082 262.752 ;
      RECT 0.048 263.424 5.082 263.520 ;
      RECT 0.048 264.192 5.082 264.288 ;
      RECT 0.048 264.960 5.082 265.056 ;
      RECT 0.048 265.728 5.082 265.824 ;
      RECT 0.048 266.496 5.082 266.592 ;
      RECT 0.048 267.264 5.082 267.360 ;
      RECT 0.048 268.032 5.082 268.128 ;
      RECT 0.048 268.800 5.082 268.896 ;
      RECT 0.048 269.568 5.082 269.664 ;
      RECT 0.048 270.336 5.082 270.432 ;
      RECT 0.048 271.104 5.082 271.200 ;
      RECT 0.048 271.872 5.082 271.968 ;
      RECT 0.048 272.640 5.082 272.736 ;
      RECT 0.048 273.408 5.082 273.504 ;
      RECT 0.048 274.176 5.082 274.272 ;
      RECT 0.048 274.944 5.082 275.040 ;
      RECT 0.048 275.712 5.082 275.808 ;
      RECT 0.048 276.480 5.082 276.576 ;
      RECT 0.048 277.248 5.082 277.344 ;
      RECT 0.048 278.016 5.082 278.112 ;
      RECT 0.048 278.784 5.082 278.880 ;
      RECT 0.048 279.552 5.082 279.648 ;
      RECT 0.048 280.320 5.082 280.416 ;
      RECT 0.048 281.088 5.082 281.184 ;
      RECT 0.048 281.856 5.082 281.952 ;
      RECT 0.048 282.624 5.082 282.720 ;
      RECT 0.048 283.392 5.082 283.488 ;
      RECT 0.048 284.160 5.082 284.256 ;
      RECT 0.048 284.928 5.082 285.024 ;
      RECT 0.048 285.696 5.082 285.792 ;
      RECT 0.048 286.464 5.082 286.560 ;
      RECT 0.048 287.232 5.082 287.328 ;
      RECT 0.048 288.000 5.082 288.096 ;
      RECT 0.048 288.768 5.082 288.864 ;
      RECT 0.048 289.536 5.082 289.632 ;
      RECT 0.048 290.304 5.082 290.400 ;
      RECT 0.048 291.072 5.082 291.168 ;
      RECT 0.048 291.840 5.082 291.936 ;
      RECT 0.048 292.608 5.082 292.704 ;
      RECT 0.048 293.376 5.082 293.472 ;
      RECT 0.048 294.144 5.082 294.240 ;
      RECT 0.048 294.912 5.082 295.008 ;
      RECT 0.048 295.680 5.082 295.776 ;
      RECT 0.048 296.448 5.082 296.544 ;
      RECT 0.048 297.216 5.082 297.312 ;
      RECT 0.048 297.984 5.082 298.080 ;
      RECT 0.048 298.752 5.082 298.848 ;
      RECT 0.048 299.520 5.082 299.616 ;
      RECT 0.048 300.288 5.082 300.384 ;
      RECT 0.048 301.056 5.082 301.152 ;
      RECT 0.048 301.824 5.082 301.920 ;
      RECT 0.048 302.592 5.082 302.688 ;
      RECT 0.048 303.360 5.082 303.456 ;
      RECT 0.048 304.128 5.082 304.224 ;
      RECT 0.048 304.896 5.082 304.992 ;
      RECT 0.048 305.664 5.082 305.760 ;
      RECT 0.048 306.432 5.082 306.528 ;
      RECT 0.048 307.200 5.082 307.296 ;
      RECT 0.048 307.968 5.082 308.064 ;
      RECT 0.048 308.736 5.082 308.832 ;
      RECT 0.048 309.504 5.082 309.600 ;
      RECT 0.048 310.272 5.082 310.368 ;
      RECT 0.048 311.040 5.082 311.136 ;
      RECT 0.048 311.808 5.082 311.904 ;
      RECT 0.048 312.576 5.082 312.672 ;
      RECT 0.048 313.344 5.082 313.440 ;
      RECT 0.048 314.112 5.082 314.208 ;
      RECT 0.048 314.880 5.082 314.976 ;
      RECT 0.048 315.648 5.082 315.744 ;
      RECT 0.048 316.416 5.082 316.512 ;
      RECT 0.048 317.184 5.082 317.280 ;
      RECT 0.048 317.952 5.082 318.048 ;
      RECT 0.048 318.720 5.082 318.816 ;
      RECT 0.048 319.488 5.082 319.584 ;
      RECT 0.048 320.256 5.082 320.352 ;
      RECT 0.048 321.024 5.082 321.120 ;
      RECT 0.048 321.792 5.082 321.888 ;
      RECT 0.048 322.560 5.082 322.656 ;
      RECT 0.048 323.328 5.082 323.424 ;
      RECT 0.048 324.096 5.082 324.192 ;
      RECT 0.048 324.864 5.082 324.960 ;
      RECT 0.048 325.632 5.082 325.728 ;
      RECT 0.048 326.400 5.082 326.496 ;
      RECT 0.048 327.168 5.082 327.264 ;
      RECT 0.048 327.936 5.082 328.032 ;
      RECT 0.048 328.704 5.082 328.800 ;
      RECT 0.048 329.472 5.082 329.568 ;
      RECT 0.048 330.240 5.082 330.336 ;
      RECT 0.048 331.008 5.082 331.104 ;
      RECT 0.048 331.776 5.082 331.872 ;
      RECT 0.048 332.544 5.082 332.640 ;
      RECT 0.048 333.312 5.082 333.408 ;
      RECT 0.048 334.080 5.082 334.176 ;
      RECT 0.048 334.848 5.082 334.944 ;
      RECT 0.048 335.616 5.082 335.712 ;
      RECT 0.048 336.384 5.082 336.480 ;
      RECT 0.048 337.152 5.082 337.248 ;
      RECT 0.048 337.920 5.082 338.016 ;
      RECT 0.048 338.688 5.082 338.784 ;
      RECT 0.048 339.456 5.082 339.552 ;
      RECT 0.048 340.224 5.082 340.320 ;
      RECT 0.048 340.992 5.082 341.088 ;
      RECT 0.048 341.760 5.082 341.856 ;
      RECT 0.048 342.528 5.082 342.624 ;
      RECT 0.048 343.296 5.082 343.392 ;
      RECT 0.048 344.064 5.082 344.160 ;
      RECT 0.048 344.832 5.082 344.928 ;
      RECT 0.048 345.600 5.082 345.696 ;
      RECT 0.048 346.368 5.082 346.464 ;
      RECT 0.048 347.136 5.082 347.232 ;
      RECT 0.048 347.904 5.082 348.000 ;
      RECT 0.048 348.672 5.082 348.768 ;
      RECT 0.048 349.440 5.082 349.536 ;
      RECT 0.048 350.208 5.082 350.304 ;
      RECT 0.048 350.976 5.082 351.072 ;
      RECT 0.048 351.744 5.082 351.840 ;
      RECT 0.048 352.512 5.082 352.608 ;
      RECT 0.048 353.280 5.082 353.376 ;
      RECT 0.048 354.048 5.082 354.144 ;
      RECT 0.048 354.816 5.082 354.912 ;
      RECT 0.048 355.584 5.082 355.680 ;
      RECT 0.048 356.352 5.082 356.448 ;
      RECT 0.048 357.120 5.082 357.216 ;
      RECT 0.048 357.888 5.082 357.984 ;
      RECT 0.048 358.656 5.082 358.752 ;
      RECT 0.048 359.424 5.082 359.520 ;
      RECT 0.048 360.192 5.082 360.288 ;
      RECT 0.048 360.960 5.082 361.056 ;
      RECT 0.048 361.728 5.082 361.824 ;
      RECT 0.048 362.496 5.082 362.592 ;
      RECT 0.048 363.264 5.082 363.360 ;
      RECT 0.048 364.032 5.082 364.128 ;
      RECT 0.048 364.800 5.082 364.896 ;
      RECT 0.048 365.568 5.082 365.664 ;
      RECT 0.048 366.336 5.082 366.432 ;
      RECT 0.048 367.104 5.082 367.200 ;
      RECT 0.048 367.872 5.082 367.968 ;
      RECT 0.048 368.640 5.082 368.736 ;
      RECT 0.048 369.408 5.082 369.504 ;
      RECT 0.048 370.176 5.082 370.272 ;
      RECT 0.048 370.944 5.082 371.040 ;
      RECT 0.048 371.712 5.082 371.808 ;
      RECT 0.048 372.480 5.082 372.576 ;
      RECT 0.048 373.248 5.082 373.344 ;
      RECT 0.048 374.016 5.082 374.112 ;
      RECT 0.048 374.784 5.082 374.880 ;
      RECT 0.048 375.552 5.082 375.648 ;
      RECT 0.048 376.320 5.082 376.416 ;
      RECT 0.048 377.088 5.082 377.184 ;
      RECT 0.048 377.856 5.082 377.952 ;
      RECT 0.048 378.624 5.082 378.720 ;
      RECT 0.048 379.392 5.082 379.488 ;
      RECT 0.048 380.160 5.082 380.256 ;
      RECT 0.048 380.928 5.082 381.024 ;
      RECT 0.048 381.696 5.082 381.792 ;
      RECT 0.048 382.464 5.082 382.560 ;
      RECT 0.048 383.232 5.082 383.328 ;
      RECT 0.048 384.000 5.082 384.096 ;
      RECT 0.048 384.768 5.082 384.864 ;
      RECT 0.048 385.536 5.082 385.632 ;
      RECT 0.048 386.304 5.082 386.400 ;
      RECT 0.048 387.072 5.082 387.168 ;
      RECT 0.048 387.840 5.082 387.936 ;
      RECT 0.048 388.608 5.082 388.704 ;
      RECT 0.048 389.376 5.082 389.472 ;
      RECT 0.048 390.144 5.082 390.240 ;
      RECT 0.048 390.912 5.082 391.008 ;
      RECT 0.048 391.680 5.082 391.776 ;
      RECT 0.048 392.448 5.082 392.544 ;
      RECT 0.048 393.216 5.082 393.312 ;
      RECT 0.048 393.984 5.082 394.080 ;
      RECT 0.048 394.752 5.082 394.848 ;
      RECT 0.048 395.520 5.082 395.616 ;
      RECT 0.048 396.288 5.082 396.384 ;
      RECT 0.048 397.056 5.082 397.152 ;
      RECT 0.048 397.824 5.082 397.920 ;
      RECT 0.048 398.592 5.082 398.688 ;
      RECT 0.048 399.360 5.082 399.456 ;
      RECT 0.048 400.128 5.082 400.224 ;
      RECT 0.048 400.896 5.082 400.992 ;
      RECT 0.048 401.664 5.082 401.760 ;
      RECT 0.048 402.432 5.082 402.528 ;
      RECT 0.048 403.200 5.082 403.296 ;
      RECT 0.048 403.968 5.082 404.064 ;
      RECT 0.048 404.736 5.082 404.832 ;
      RECT 0.048 405.504 5.082 405.600 ;
      RECT 0.048 406.272 5.082 406.368 ;
      RECT 0.048 407.040 5.082 407.136 ;
      RECT 0.048 407.808 5.082 407.904 ;
      RECT 0.048 408.576 5.082 408.672 ;
      RECT 0.048 409.344 5.082 409.440 ;
      RECT 0.048 410.112 5.082 410.208 ;
      RECT 0.048 410.880 5.082 410.976 ;
      RECT 0.048 411.648 5.082 411.744 ;
      RECT 0.048 412.416 5.082 412.512 ;
      RECT 0.048 413.184 5.082 413.280 ;
      RECT 0.048 413.952 5.082 414.048 ;
      RECT 0.048 414.720 5.082 414.816 ;
      RECT 0.048 415.488 5.082 415.584 ;
      RECT 0.048 416.256 5.082 416.352 ;
      RECT 0.048 417.024 5.082 417.120 ;
      RECT 0.048 417.792 5.082 417.888 ;
      RECT 0.048 418.560 5.082 418.656 ;
      RECT 0.048 419.328 5.082 419.424 ;
      RECT 0.048 420.096 5.082 420.192 ;
      RECT 0.048 420.864 5.082 420.960 ;
      RECT 0.048 421.632 5.082 421.728 ;
      RECT 0.048 422.400 5.082 422.496 ;
      RECT 0.048 423.168 5.082 423.264 ;
      RECT 0.048 423.936 5.082 424.032 ;
      RECT 0.048 424.704 5.082 424.800 ;
      RECT 0.048 425.472 5.082 425.568 ;
      RECT 0.048 426.240 5.082 426.336 ;
      RECT 0.048 427.008 5.082 427.104 ;
      RECT 0.048 427.776 5.082 427.872 ;
      RECT 0.048 428.544 5.082 428.640 ;
      RECT 0.048 429.312 5.082 429.408 ;
      RECT 0.048 430.080 5.082 430.176 ;
      RECT 0.048 430.848 5.082 430.944 ;
      RECT 0.048 431.616 5.082 431.712 ;
      RECT 0.048 432.384 5.082 432.480 ;
      RECT 0.048 433.152 5.082 433.248 ;
      RECT 0.048 433.920 5.082 434.016 ;
      RECT 0.048 434.688 5.082 434.784 ;
      RECT 0.048 435.456 5.082 435.552 ;
      RECT 0.048 436.224 5.082 436.320 ;
      RECT 0.048 436.992 5.082 437.088 ;
      RECT 0.048 437.760 5.082 437.856 ;
      RECT 0.048 438.528 5.082 438.624 ;
      RECT 0.048 439.296 5.082 439.392 ;
      RECT 0.048 440.064 5.082 440.160 ;
      RECT 0.048 440.832 5.082 440.928 ;
      RECT 0.048 441.600 5.082 441.696 ;
      RECT 0.048 442.368 5.082 442.464 ;
      RECT 0.048 443.136 5.082 443.232 ;
      RECT 0.048 443.904 5.082 444.000 ;
      RECT 0.048 444.672 5.082 444.768 ;
      RECT 0.048 445.440 5.082 445.536 ;
      RECT 0.048 446.208 5.082 446.304 ;
      RECT 0.048 446.976 5.082 447.072 ;
      RECT 0.048 447.744 5.082 447.840 ;
      RECT 0.048 448.512 5.082 448.608 ;
      RECT 0.048 449.280 5.082 449.376 ;
      RECT 0.048 450.048 5.082 450.144 ;
      RECT 0.048 450.816 5.082 450.912 ;
      RECT 0.048 451.584 5.082 451.680 ;
      RECT 0.048 452.352 5.082 452.448 ;
      RECT 0.048 453.120 5.082 453.216 ;
      RECT 0.048 453.888 5.082 453.984 ;
      RECT 0.048 454.656 5.082 454.752 ;
      RECT 0.048 455.424 5.082 455.520 ;
      RECT 0.048 456.192 5.082 456.288 ;
      RECT 0.048 456.960 5.082 457.056 ;
      RECT 0.048 457.728 5.082 457.824 ;
      RECT 0.048 458.496 5.082 458.592 ;
      RECT 0.048 459.264 5.082 459.360 ;
      RECT 0.048 460.032 5.082 460.128 ;
      RECT 0.048 460.800 5.082 460.896 ;
      RECT 0.048 461.568 5.082 461.664 ;
      RECT 0.048 462.336 5.082 462.432 ;
      RECT 0.048 463.104 5.082 463.200 ;
      RECT 0.048 463.872 5.082 463.968 ;
      RECT 0.048 464.640 5.082 464.736 ;
      RECT 0.048 465.408 5.082 465.504 ;
      RECT 0.048 466.176 5.082 466.272 ;
      RECT 0.048 466.944 5.082 467.040 ;
      RECT 0.048 467.712 5.082 467.808 ;
      RECT 0.048 468.480 5.082 468.576 ;
      RECT 0.048 469.248 5.082 469.344 ;
      RECT 0.048 470.016 5.082 470.112 ;
      RECT 0.048 470.784 5.082 470.880 ;
      RECT 0.048 471.552 5.082 471.648 ;
      RECT 0.048 472.320 5.082 472.416 ;
      RECT 0.048 473.088 5.082 473.184 ;
      RECT 0.048 473.856 5.082 473.952 ;
      RECT 0.048 474.624 5.082 474.720 ;
      RECT 0.048 475.392 5.082 475.488 ;
      RECT 0.048 476.160 5.082 476.256 ;
      RECT 0.048 476.928 5.082 477.024 ;
      RECT 0.048 477.696 5.082 477.792 ;
      RECT 0.048 478.464 5.082 478.560 ;
      RECT 0.048 479.232 5.082 479.328 ;
      RECT 0.048 480.000 5.082 480.096 ;
      RECT 0.048 480.768 5.082 480.864 ;
      RECT 0.048 481.536 5.082 481.632 ;
      RECT 0.048 482.304 5.082 482.400 ;
      RECT 0.048 483.072 5.082 483.168 ;
      RECT 0.048 483.840 5.082 483.936 ;
      RECT 0.048 484.608 5.082 484.704 ;
      RECT 0.048 485.376 5.082 485.472 ;
      RECT 0.048 486.144 5.082 486.240 ;
      RECT 0.048 486.912 5.082 487.008 ;
      RECT 0.048 487.680 5.082 487.776 ;
      RECT 0.048 488.448 5.082 488.544 ;
      RECT 0.048 489.216 5.082 489.312 ;
      RECT 0.048 489.984 5.082 490.080 ;
      RECT 0.048 490.752 5.082 490.848 ;
      RECT 0.048 491.520 5.082 491.616 ;
      RECT 0.048 492.288 5.082 492.384 ;
      RECT 0.048 493.056 5.082 493.152 ;
      RECT 0.048 493.824 5.082 493.920 ;
      RECT 0.048 494.592 5.082 494.688 ;
      RECT 0.048 495.360 5.082 495.456 ;
      RECT 0.048 496.128 5.082 496.224 ;
      RECT 0.048 496.896 5.082 496.992 ;
      RECT 0.048 497.664 5.082 497.760 ;
      RECT 0.048 498.432 5.082 498.528 ;
      RECT 0.048 499.200 5.082 499.296 ;
      RECT 0.048 499.968 5.082 500.064 ;
      RECT 0.048 500.736 5.082 500.832 ;
      RECT 0.048 501.504 5.082 501.600 ;
      RECT 0.048 502.272 5.082 502.368 ;
      RECT 0.048 503.040 5.082 503.136 ;
      RECT 0.048 503.808 5.082 503.904 ;
      RECT 0.048 504.576 5.082 504.672 ;
      RECT 0.048 505.344 5.082 505.440 ;
      RECT 0.048 506.112 5.082 506.208 ;
      RECT 0.048 506.880 5.082 506.976 ;
      RECT 0.048 507.648 5.082 507.744 ;
      RECT 0.048 508.416 5.082 508.512 ;
      RECT 0.048 509.184 5.082 509.280 ;
      RECT 0.048 509.952 5.082 510.048 ;
      RECT 0.048 510.720 5.082 510.816 ;
      RECT 0.048 511.488 5.082 511.584 ;
      RECT 0.048 512.256 5.082 512.352 ;
      RECT 0.048 513.024 5.082 513.120 ;
      RECT 0.048 513.792 5.082 513.888 ;
      RECT 0.048 514.560 5.082 514.656 ;
      RECT 0.048 515.328 5.082 515.424 ;
      RECT 0.048 516.096 5.082 516.192 ;
      RECT 0.048 516.864 5.082 516.960 ;
      RECT 0.048 517.632 5.082 517.728 ;
      RECT 0.048 518.400 5.082 518.496 ;
      RECT 0.048 519.168 5.082 519.264 ;
      RECT 0.048 519.936 5.082 520.032 ;
      RECT 0.048 520.704 5.082 520.800 ;
      RECT 0.048 521.472 5.082 521.568 ;
      RECT 0.048 522.240 5.082 522.336 ;
      RECT 0.048 523.008 5.082 523.104 ;
      RECT 0.048 523.776 5.082 523.872 ;
      RECT 0.048 524.544 5.082 524.640 ;
      RECT 0.048 525.312 5.082 525.408 ;
      RECT 0.048 526.080 5.082 526.176 ;
      RECT 0.048 526.848 5.082 526.944 ;
      RECT 0.048 527.616 5.082 527.712 ;
      RECT 0.048 528.384 5.082 528.480 ;
      RECT 0.048 529.152 5.082 529.248 ;
      RECT 0.048 529.920 5.082 530.016 ;
      RECT 0.048 530.688 5.082 530.784 ;
      RECT 0.048 531.456 5.082 531.552 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.384 5.082 0.480 ;
      RECT 0.048 1.152 5.082 1.248 ;
      RECT 0.048 1.920 5.082 2.016 ;
      RECT 0.048 2.688 5.082 2.784 ;
      RECT 0.048 3.456 5.082 3.552 ;
      RECT 0.048 4.224 5.082 4.320 ;
      RECT 0.048 4.992 5.082 5.088 ;
      RECT 0.048 5.760 5.082 5.856 ;
      RECT 0.048 6.528 5.082 6.624 ;
      RECT 0.048 7.296 5.082 7.392 ;
      RECT 0.048 8.064 5.082 8.160 ;
      RECT 0.048 8.832 5.082 8.928 ;
      RECT 0.048 9.600 5.082 9.696 ;
      RECT 0.048 10.368 5.082 10.464 ;
      RECT 0.048 11.136 5.082 11.232 ;
      RECT 0.048 11.904 5.082 12.000 ;
      RECT 0.048 12.672 5.082 12.768 ;
      RECT 0.048 13.440 5.082 13.536 ;
      RECT 0.048 14.208 5.082 14.304 ;
      RECT 0.048 14.976 5.082 15.072 ;
      RECT 0.048 15.744 5.082 15.840 ;
      RECT 0.048 16.512 5.082 16.608 ;
      RECT 0.048 17.280 5.082 17.376 ;
      RECT 0.048 18.048 5.082 18.144 ;
      RECT 0.048 18.816 5.082 18.912 ;
      RECT 0.048 19.584 5.082 19.680 ;
      RECT 0.048 20.352 5.082 20.448 ;
      RECT 0.048 21.120 5.082 21.216 ;
      RECT 0.048 21.888 5.082 21.984 ;
      RECT 0.048 22.656 5.082 22.752 ;
      RECT 0.048 23.424 5.082 23.520 ;
      RECT 0.048 24.192 5.082 24.288 ;
      RECT 0.048 24.960 5.082 25.056 ;
      RECT 0.048 25.728 5.082 25.824 ;
      RECT 0.048 26.496 5.082 26.592 ;
      RECT 0.048 27.264 5.082 27.360 ;
      RECT 0.048 28.032 5.082 28.128 ;
      RECT 0.048 28.800 5.082 28.896 ;
      RECT 0.048 29.568 5.082 29.664 ;
      RECT 0.048 30.336 5.082 30.432 ;
      RECT 0.048 31.104 5.082 31.200 ;
      RECT 0.048 31.872 5.082 31.968 ;
      RECT 0.048 32.640 5.082 32.736 ;
      RECT 0.048 33.408 5.082 33.504 ;
      RECT 0.048 34.176 5.082 34.272 ;
      RECT 0.048 34.944 5.082 35.040 ;
      RECT 0.048 35.712 5.082 35.808 ;
      RECT 0.048 36.480 5.082 36.576 ;
      RECT 0.048 37.248 5.082 37.344 ;
      RECT 0.048 38.016 5.082 38.112 ;
      RECT 0.048 38.784 5.082 38.880 ;
      RECT 0.048 39.552 5.082 39.648 ;
      RECT 0.048 40.320 5.082 40.416 ;
      RECT 0.048 41.088 5.082 41.184 ;
      RECT 0.048 41.856 5.082 41.952 ;
      RECT 0.048 42.624 5.082 42.720 ;
      RECT 0.048 43.392 5.082 43.488 ;
      RECT 0.048 44.160 5.082 44.256 ;
      RECT 0.048 44.928 5.082 45.024 ;
      RECT 0.048 45.696 5.082 45.792 ;
      RECT 0.048 46.464 5.082 46.560 ;
      RECT 0.048 47.232 5.082 47.328 ;
      RECT 0.048 48.000 5.082 48.096 ;
      RECT 0.048 48.768 5.082 48.864 ;
      RECT 0.048 49.536 5.082 49.632 ;
      RECT 0.048 50.304 5.082 50.400 ;
      RECT 0.048 51.072 5.082 51.168 ;
      RECT 0.048 51.840 5.082 51.936 ;
      RECT 0.048 52.608 5.082 52.704 ;
      RECT 0.048 53.376 5.082 53.472 ;
      RECT 0.048 54.144 5.082 54.240 ;
      RECT 0.048 54.912 5.082 55.008 ;
      RECT 0.048 55.680 5.082 55.776 ;
      RECT 0.048 56.448 5.082 56.544 ;
      RECT 0.048 57.216 5.082 57.312 ;
      RECT 0.048 57.984 5.082 58.080 ;
      RECT 0.048 58.752 5.082 58.848 ;
      RECT 0.048 59.520 5.082 59.616 ;
      RECT 0.048 60.288 5.082 60.384 ;
      RECT 0.048 61.056 5.082 61.152 ;
      RECT 0.048 61.824 5.082 61.920 ;
      RECT 0.048 62.592 5.082 62.688 ;
      RECT 0.048 63.360 5.082 63.456 ;
      RECT 0.048 64.128 5.082 64.224 ;
      RECT 0.048 64.896 5.082 64.992 ;
      RECT 0.048 65.664 5.082 65.760 ;
      RECT 0.048 66.432 5.082 66.528 ;
      RECT 0.048 67.200 5.082 67.296 ;
      RECT 0.048 67.968 5.082 68.064 ;
      RECT 0.048 68.736 5.082 68.832 ;
      RECT 0.048 69.504 5.082 69.600 ;
      RECT 0.048 70.272 5.082 70.368 ;
      RECT 0.048 71.040 5.082 71.136 ;
      RECT 0.048 71.808 5.082 71.904 ;
      RECT 0.048 72.576 5.082 72.672 ;
      RECT 0.048 73.344 5.082 73.440 ;
      RECT 0.048 74.112 5.082 74.208 ;
      RECT 0.048 74.880 5.082 74.976 ;
      RECT 0.048 75.648 5.082 75.744 ;
      RECT 0.048 76.416 5.082 76.512 ;
      RECT 0.048 77.184 5.082 77.280 ;
      RECT 0.048 77.952 5.082 78.048 ;
      RECT 0.048 78.720 5.082 78.816 ;
      RECT 0.048 79.488 5.082 79.584 ;
      RECT 0.048 80.256 5.082 80.352 ;
      RECT 0.048 81.024 5.082 81.120 ;
      RECT 0.048 81.792 5.082 81.888 ;
      RECT 0.048 82.560 5.082 82.656 ;
      RECT 0.048 83.328 5.082 83.424 ;
      RECT 0.048 84.096 5.082 84.192 ;
      RECT 0.048 84.864 5.082 84.960 ;
      RECT 0.048 85.632 5.082 85.728 ;
      RECT 0.048 86.400 5.082 86.496 ;
      RECT 0.048 87.168 5.082 87.264 ;
      RECT 0.048 87.936 5.082 88.032 ;
      RECT 0.048 88.704 5.082 88.800 ;
      RECT 0.048 89.472 5.082 89.568 ;
      RECT 0.048 90.240 5.082 90.336 ;
      RECT 0.048 91.008 5.082 91.104 ;
      RECT 0.048 91.776 5.082 91.872 ;
      RECT 0.048 92.544 5.082 92.640 ;
      RECT 0.048 93.312 5.082 93.408 ;
      RECT 0.048 94.080 5.082 94.176 ;
      RECT 0.048 94.848 5.082 94.944 ;
      RECT 0.048 95.616 5.082 95.712 ;
      RECT 0.048 96.384 5.082 96.480 ;
      RECT 0.048 97.152 5.082 97.248 ;
      RECT 0.048 97.920 5.082 98.016 ;
      RECT 0.048 98.688 5.082 98.784 ;
      RECT 0.048 99.456 5.082 99.552 ;
      RECT 0.048 100.224 5.082 100.320 ;
      RECT 0.048 100.992 5.082 101.088 ;
      RECT 0.048 101.760 5.082 101.856 ;
      RECT 0.048 102.528 5.082 102.624 ;
      RECT 0.048 103.296 5.082 103.392 ;
      RECT 0.048 104.064 5.082 104.160 ;
      RECT 0.048 104.832 5.082 104.928 ;
      RECT 0.048 105.600 5.082 105.696 ;
      RECT 0.048 106.368 5.082 106.464 ;
      RECT 0.048 107.136 5.082 107.232 ;
      RECT 0.048 107.904 5.082 108.000 ;
      RECT 0.048 108.672 5.082 108.768 ;
      RECT 0.048 109.440 5.082 109.536 ;
      RECT 0.048 110.208 5.082 110.304 ;
      RECT 0.048 110.976 5.082 111.072 ;
      RECT 0.048 111.744 5.082 111.840 ;
      RECT 0.048 112.512 5.082 112.608 ;
      RECT 0.048 113.280 5.082 113.376 ;
      RECT 0.048 114.048 5.082 114.144 ;
      RECT 0.048 114.816 5.082 114.912 ;
      RECT 0.048 115.584 5.082 115.680 ;
      RECT 0.048 116.352 5.082 116.448 ;
      RECT 0.048 117.120 5.082 117.216 ;
      RECT 0.048 117.888 5.082 117.984 ;
      RECT 0.048 118.656 5.082 118.752 ;
      RECT 0.048 119.424 5.082 119.520 ;
      RECT 0.048 120.192 5.082 120.288 ;
      RECT 0.048 120.960 5.082 121.056 ;
      RECT 0.048 121.728 5.082 121.824 ;
      RECT 0.048 122.496 5.082 122.592 ;
      RECT 0.048 123.264 5.082 123.360 ;
      RECT 0.048 124.032 5.082 124.128 ;
      RECT 0.048 124.800 5.082 124.896 ;
      RECT 0.048 125.568 5.082 125.664 ;
      RECT 0.048 126.336 5.082 126.432 ;
      RECT 0.048 127.104 5.082 127.200 ;
      RECT 0.048 127.872 5.082 127.968 ;
      RECT 0.048 128.640 5.082 128.736 ;
      RECT 0.048 129.408 5.082 129.504 ;
      RECT 0.048 130.176 5.082 130.272 ;
      RECT 0.048 130.944 5.082 131.040 ;
      RECT 0.048 131.712 5.082 131.808 ;
      RECT 0.048 132.480 5.082 132.576 ;
      RECT 0.048 133.248 5.082 133.344 ;
      RECT 0.048 134.016 5.082 134.112 ;
      RECT 0.048 134.784 5.082 134.880 ;
      RECT 0.048 135.552 5.082 135.648 ;
      RECT 0.048 136.320 5.082 136.416 ;
      RECT 0.048 137.088 5.082 137.184 ;
      RECT 0.048 137.856 5.082 137.952 ;
      RECT 0.048 138.624 5.082 138.720 ;
      RECT 0.048 139.392 5.082 139.488 ;
      RECT 0.048 140.160 5.082 140.256 ;
      RECT 0.048 140.928 5.082 141.024 ;
      RECT 0.048 141.696 5.082 141.792 ;
      RECT 0.048 142.464 5.082 142.560 ;
      RECT 0.048 143.232 5.082 143.328 ;
      RECT 0.048 144.000 5.082 144.096 ;
      RECT 0.048 144.768 5.082 144.864 ;
      RECT 0.048 145.536 5.082 145.632 ;
      RECT 0.048 146.304 5.082 146.400 ;
      RECT 0.048 147.072 5.082 147.168 ;
      RECT 0.048 147.840 5.082 147.936 ;
      RECT 0.048 148.608 5.082 148.704 ;
      RECT 0.048 149.376 5.082 149.472 ;
      RECT 0.048 150.144 5.082 150.240 ;
      RECT 0.048 150.912 5.082 151.008 ;
      RECT 0.048 151.680 5.082 151.776 ;
      RECT 0.048 152.448 5.082 152.544 ;
      RECT 0.048 153.216 5.082 153.312 ;
      RECT 0.048 153.984 5.082 154.080 ;
      RECT 0.048 154.752 5.082 154.848 ;
      RECT 0.048 155.520 5.082 155.616 ;
      RECT 0.048 156.288 5.082 156.384 ;
      RECT 0.048 157.056 5.082 157.152 ;
      RECT 0.048 157.824 5.082 157.920 ;
      RECT 0.048 158.592 5.082 158.688 ;
      RECT 0.048 159.360 5.082 159.456 ;
      RECT 0.048 160.128 5.082 160.224 ;
      RECT 0.048 160.896 5.082 160.992 ;
      RECT 0.048 161.664 5.082 161.760 ;
      RECT 0.048 162.432 5.082 162.528 ;
      RECT 0.048 163.200 5.082 163.296 ;
      RECT 0.048 163.968 5.082 164.064 ;
      RECT 0.048 164.736 5.082 164.832 ;
      RECT 0.048 165.504 5.082 165.600 ;
      RECT 0.048 166.272 5.082 166.368 ;
      RECT 0.048 167.040 5.082 167.136 ;
      RECT 0.048 167.808 5.082 167.904 ;
      RECT 0.048 168.576 5.082 168.672 ;
      RECT 0.048 169.344 5.082 169.440 ;
      RECT 0.048 170.112 5.082 170.208 ;
      RECT 0.048 170.880 5.082 170.976 ;
      RECT 0.048 171.648 5.082 171.744 ;
      RECT 0.048 172.416 5.082 172.512 ;
      RECT 0.048 173.184 5.082 173.280 ;
      RECT 0.048 173.952 5.082 174.048 ;
      RECT 0.048 174.720 5.082 174.816 ;
      RECT 0.048 175.488 5.082 175.584 ;
      RECT 0.048 176.256 5.082 176.352 ;
      RECT 0.048 177.024 5.082 177.120 ;
      RECT 0.048 177.792 5.082 177.888 ;
      RECT 0.048 178.560 5.082 178.656 ;
      RECT 0.048 179.328 5.082 179.424 ;
      RECT 0.048 180.096 5.082 180.192 ;
      RECT 0.048 180.864 5.082 180.960 ;
      RECT 0.048 181.632 5.082 181.728 ;
      RECT 0.048 182.400 5.082 182.496 ;
      RECT 0.048 183.168 5.082 183.264 ;
      RECT 0.048 183.936 5.082 184.032 ;
      RECT 0.048 184.704 5.082 184.800 ;
      RECT 0.048 185.472 5.082 185.568 ;
      RECT 0.048 186.240 5.082 186.336 ;
      RECT 0.048 187.008 5.082 187.104 ;
      RECT 0.048 187.776 5.082 187.872 ;
      RECT 0.048 188.544 5.082 188.640 ;
      RECT 0.048 189.312 5.082 189.408 ;
      RECT 0.048 190.080 5.082 190.176 ;
      RECT 0.048 190.848 5.082 190.944 ;
      RECT 0.048 191.616 5.082 191.712 ;
      RECT 0.048 192.384 5.082 192.480 ;
      RECT 0.048 193.152 5.082 193.248 ;
      RECT 0.048 193.920 5.082 194.016 ;
      RECT 0.048 194.688 5.082 194.784 ;
      RECT 0.048 195.456 5.082 195.552 ;
      RECT 0.048 196.224 5.082 196.320 ;
      RECT 0.048 196.992 5.082 197.088 ;
      RECT 0.048 197.760 5.082 197.856 ;
      RECT 0.048 198.528 5.082 198.624 ;
      RECT 0.048 199.296 5.082 199.392 ;
      RECT 0.048 200.064 5.082 200.160 ;
      RECT 0.048 200.832 5.082 200.928 ;
      RECT 0.048 201.600 5.082 201.696 ;
      RECT 0.048 202.368 5.082 202.464 ;
      RECT 0.048 203.136 5.082 203.232 ;
      RECT 0.048 203.904 5.082 204.000 ;
      RECT 0.048 204.672 5.082 204.768 ;
      RECT 0.048 205.440 5.082 205.536 ;
      RECT 0.048 206.208 5.082 206.304 ;
      RECT 0.048 206.976 5.082 207.072 ;
      RECT 0.048 207.744 5.082 207.840 ;
      RECT 0.048 208.512 5.082 208.608 ;
      RECT 0.048 209.280 5.082 209.376 ;
      RECT 0.048 210.048 5.082 210.144 ;
      RECT 0.048 210.816 5.082 210.912 ;
      RECT 0.048 211.584 5.082 211.680 ;
      RECT 0.048 212.352 5.082 212.448 ;
      RECT 0.048 213.120 5.082 213.216 ;
      RECT 0.048 213.888 5.082 213.984 ;
      RECT 0.048 214.656 5.082 214.752 ;
      RECT 0.048 215.424 5.082 215.520 ;
      RECT 0.048 216.192 5.082 216.288 ;
      RECT 0.048 216.960 5.082 217.056 ;
      RECT 0.048 217.728 5.082 217.824 ;
      RECT 0.048 218.496 5.082 218.592 ;
      RECT 0.048 219.264 5.082 219.360 ;
      RECT 0.048 220.032 5.082 220.128 ;
      RECT 0.048 220.800 5.082 220.896 ;
      RECT 0.048 221.568 5.082 221.664 ;
      RECT 0.048 222.336 5.082 222.432 ;
      RECT 0.048 223.104 5.082 223.200 ;
      RECT 0.048 223.872 5.082 223.968 ;
      RECT 0.048 224.640 5.082 224.736 ;
      RECT 0.048 225.408 5.082 225.504 ;
      RECT 0.048 226.176 5.082 226.272 ;
      RECT 0.048 226.944 5.082 227.040 ;
      RECT 0.048 227.712 5.082 227.808 ;
      RECT 0.048 228.480 5.082 228.576 ;
      RECT 0.048 229.248 5.082 229.344 ;
      RECT 0.048 230.016 5.082 230.112 ;
      RECT 0.048 230.784 5.082 230.880 ;
      RECT 0.048 231.552 5.082 231.648 ;
      RECT 0.048 232.320 5.082 232.416 ;
      RECT 0.048 233.088 5.082 233.184 ;
      RECT 0.048 233.856 5.082 233.952 ;
      RECT 0.048 234.624 5.082 234.720 ;
      RECT 0.048 235.392 5.082 235.488 ;
      RECT 0.048 236.160 5.082 236.256 ;
      RECT 0.048 236.928 5.082 237.024 ;
      RECT 0.048 237.696 5.082 237.792 ;
      RECT 0.048 238.464 5.082 238.560 ;
      RECT 0.048 239.232 5.082 239.328 ;
      RECT 0.048 240.000 5.082 240.096 ;
      RECT 0.048 240.768 5.082 240.864 ;
      RECT 0.048 241.536 5.082 241.632 ;
      RECT 0.048 242.304 5.082 242.400 ;
      RECT 0.048 243.072 5.082 243.168 ;
      RECT 0.048 243.840 5.082 243.936 ;
      RECT 0.048 244.608 5.082 244.704 ;
      RECT 0.048 245.376 5.082 245.472 ;
      RECT 0.048 246.144 5.082 246.240 ;
      RECT 0.048 246.912 5.082 247.008 ;
      RECT 0.048 247.680 5.082 247.776 ;
      RECT 0.048 248.448 5.082 248.544 ;
      RECT 0.048 249.216 5.082 249.312 ;
      RECT 0.048 249.984 5.082 250.080 ;
      RECT 0.048 250.752 5.082 250.848 ;
      RECT 0.048 251.520 5.082 251.616 ;
      RECT 0.048 252.288 5.082 252.384 ;
      RECT 0.048 253.056 5.082 253.152 ;
      RECT 0.048 253.824 5.082 253.920 ;
      RECT 0.048 254.592 5.082 254.688 ;
      RECT 0.048 255.360 5.082 255.456 ;
      RECT 0.048 256.128 5.082 256.224 ;
      RECT 0.048 256.896 5.082 256.992 ;
      RECT 0.048 257.664 5.082 257.760 ;
      RECT 0.048 258.432 5.082 258.528 ;
      RECT 0.048 259.200 5.082 259.296 ;
      RECT 0.048 259.968 5.082 260.064 ;
      RECT 0.048 260.736 5.082 260.832 ;
      RECT 0.048 261.504 5.082 261.600 ;
      RECT 0.048 262.272 5.082 262.368 ;
      RECT 0.048 263.040 5.082 263.136 ;
      RECT 0.048 263.808 5.082 263.904 ;
      RECT 0.048 264.576 5.082 264.672 ;
      RECT 0.048 265.344 5.082 265.440 ;
      RECT 0.048 266.112 5.082 266.208 ;
      RECT 0.048 266.880 5.082 266.976 ;
      RECT 0.048 267.648 5.082 267.744 ;
      RECT 0.048 268.416 5.082 268.512 ;
      RECT 0.048 269.184 5.082 269.280 ;
      RECT 0.048 269.952 5.082 270.048 ;
      RECT 0.048 270.720 5.082 270.816 ;
      RECT 0.048 271.488 5.082 271.584 ;
      RECT 0.048 272.256 5.082 272.352 ;
      RECT 0.048 273.024 5.082 273.120 ;
      RECT 0.048 273.792 5.082 273.888 ;
      RECT 0.048 274.560 5.082 274.656 ;
      RECT 0.048 275.328 5.082 275.424 ;
      RECT 0.048 276.096 5.082 276.192 ;
      RECT 0.048 276.864 5.082 276.960 ;
      RECT 0.048 277.632 5.082 277.728 ;
      RECT 0.048 278.400 5.082 278.496 ;
      RECT 0.048 279.168 5.082 279.264 ;
      RECT 0.048 279.936 5.082 280.032 ;
      RECT 0.048 280.704 5.082 280.800 ;
      RECT 0.048 281.472 5.082 281.568 ;
      RECT 0.048 282.240 5.082 282.336 ;
      RECT 0.048 283.008 5.082 283.104 ;
      RECT 0.048 283.776 5.082 283.872 ;
      RECT 0.048 284.544 5.082 284.640 ;
      RECT 0.048 285.312 5.082 285.408 ;
      RECT 0.048 286.080 5.082 286.176 ;
      RECT 0.048 286.848 5.082 286.944 ;
      RECT 0.048 287.616 5.082 287.712 ;
      RECT 0.048 288.384 5.082 288.480 ;
      RECT 0.048 289.152 5.082 289.248 ;
      RECT 0.048 289.920 5.082 290.016 ;
      RECT 0.048 290.688 5.082 290.784 ;
      RECT 0.048 291.456 5.082 291.552 ;
      RECT 0.048 292.224 5.082 292.320 ;
      RECT 0.048 292.992 5.082 293.088 ;
      RECT 0.048 293.760 5.082 293.856 ;
      RECT 0.048 294.528 5.082 294.624 ;
      RECT 0.048 295.296 5.082 295.392 ;
      RECT 0.048 296.064 5.082 296.160 ;
      RECT 0.048 296.832 5.082 296.928 ;
      RECT 0.048 297.600 5.082 297.696 ;
      RECT 0.048 298.368 5.082 298.464 ;
      RECT 0.048 299.136 5.082 299.232 ;
      RECT 0.048 299.904 5.082 300.000 ;
      RECT 0.048 300.672 5.082 300.768 ;
      RECT 0.048 301.440 5.082 301.536 ;
      RECT 0.048 302.208 5.082 302.304 ;
      RECT 0.048 302.976 5.082 303.072 ;
      RECT 0.048 303.744 5.082 303.840 ;
      RECT 0.048 304.512 5.082 304.608 ;
      RECT 0.048 305.280 5.082 305.376 ;
      RECT 0.048 306.048 5.082 306.144 ;
      RECT 0.048 306.816 5.082 306.912 ;
      RECT 0.048 307.584 5.082 307.680 ;
      RECT 0.048 308.352 5.082 308.448 ;
      RECT 0.048 309.120 5.082 309.216 ;
      RECT 0.048 309.888 5.082 309.984 ;
      RECT 0.048 310.656 5.082 310.752 ;
      RECT 0.048 311.424 5.082 311.520 ;
      RECT 0.048 312.192 5.082 312.288 ;
      RECT 0.048 312.960 5.082 313.056 ;
      RECT 0.048 313.728 5.082 313.824 ;
      RECT 0.048 314.496 5.082 314.592 ;
      RECT 0.048 315.264 5.082 315.360 ;
      RECT 0.048 316.032 5.082 316.128 ;
      RECT 0.048 316.800 5.082 316.896 ;
      RECT 0.048 317.568 5.082 317.664 ;
      RECT 0.048 318.336 5.082 318.432 ;
      RECT 0.048 319.104 5.082 319.200 ;
      RECT 0.048 319.872 5.082 319.968 ;
      RECT 0.048 320.640 5.082 320.736 ;
      RECT 0.048 321.408 5.082 321.504 ;
      RECT 0.048 322.176 5.082 322.272 ;
      RECT 0.048 322.944 5.082 323.040 ;
      RECT 0.048 323.712 5.082 323.808 ;
      RECT 0.048 324.480 5.082 324.576 ;
      RECT 0.048 325.248 5.082 325.344 ;
      RECT 0.048 326.016 5.082 326.112 ;
      RECT 0.048 326.784 5.082 326.880 ;
      RECT 0.048 327.552 5.082 327.648 ;
      RECT 0.048 328.320 5.082 328.416 ;
      RECT 0.048 329.088 5.082 329.184 ;
      RECT 0.048 329.856 5.082 329.952 ;
      RECT 0.048 330.624 5.082 330.720 ;
      RECT 0.048 331.392 5.082 331.488 ;
      RECT 0.048 332.160 5.082 332.256 ;
      RECT 0.048 332.928 5.082 333.024 ;
      RECT 0.048 333.696 5.082 333.792 ;
      RECT 0.048 334.464 5.082 334.560 ;
      RECT 0.048 335.232 5.082 335.328 ;
      RECT 0.048 336.000 5.082 336.096 ;
      RECT 0.048 336.768 5.082 336.864 ;
      RECT 0.048 337.536 5.082 337.632 ;
      RECT 0.048 338.304 5.082 338.400 ;
      RECT 0.048 339.072 5.082 339.168 ;
      RECT 0.048 339.840 5.082 339.936 ;
      RECT 0.048 340.608 5.082 340.704 ;
      RECT 0.048 341.376 5.082 341.472 ;
      RECT 0.048 342.144 5.082 342.240 ;
      RECT 0.048 342.912 5.082 343.008 ;
      RECT 0.048 343.680 5.082 343.776 ;
      RECT 0.048 344.448 5.082 344.544 ;
      RECT 0.048 345.216 5.082 345.312 ;
      RECT 0.048 345.984 5.082 346.080 ;
      RECT 0.048 346.752 5.082 346.848 ;
      RECT 0.048 347.520 5.082 347.616 ;
      RECT 0.048 348.288 5.082 348.384 ;
      RECT 0.048 349.056 5.082 349.152 ;
      RECT 0.048 349.824 5.082 349.920 ;
      RECT 0.048 350.592 5.082 350.688 ;
      RECT 0.048 351.360 5.082 351.456 ;
      RECT 0.048 352.128 5.082 352.224 ;
      RECT 0.048 352.896 5.082 352.992 ;
      RECT 0.048 353.664 5.082 353.760 ;
      RECT 0.048 354.432 5.082 354.528 ;
      RECT 0.048 355.200 5.082 355.296 ;
      RECT 0.048 355.968 5.082 356.064 ;
      RECT 0.048 356.736 5.082 356.832 ;
      RECT 0.048 357.504 5.082 357.600 ;
      RECT 0.048 358.272 5.082 358.368 ;
      RECT 0.048 359.040 5.082 359.136 ;
      RECT 0.048 359.808 5.082 359.904 ;
      RECT 0.048 360.576 5.082 360.672 ;
      RECT 0.048 361.344 5.082 361.440 ;
      RECT 0.048 362.112 5.082 362.208 ;
      RECT 0.048 362.880 5.082 362.976 ;
      RECT 0.048 363.648 5.082 363.744 ;
      RECT 0.048 364.416 5.082 364.512 ;
      RECT 0.048 365.184 5.082 365.280 ;
      RECT 0.048 365.952 5.082 366.048 ;
      RECT 0.048 366.720 5.082 366.816 ;
      RECT 0.048 367.488 5.082 367.584 ;
      RECT 0.048 368.256 5.082 368.352 ;
      RECT 0.048 369.024 5.082 369.120 ;
      RECT 0.048 369.792 5.082 369.888 ;
      RECT 0.048 370.560 5.082 370.656 ;
      RECT 0.048 371.328 5.082 371.424 ;
      RECT 0.048 372.096 5.082 372.192 ;
      RECT 0.048 372.864 5.082 372.960 ;
      RECT 0.048 373.632 5.082 373.728 ;
      RECT 0.048 374.400 5.082 374.496 ;
      RECT 0.048 375.168 5.082 375.264 ;
      RECT 0.048 375.936 5.082 376.032 ;
      RECT 0.048 376.704 5.082 376.800 ;
      RECT 0.048 377.472 5.082 377.568 ;
      RECT 0.048 378.240 5.082 378.336 ;
      RECT 0.048 379.008 5.082 379.104 ;
      RECT 0.048 379.776 5.082 379.872 ;
      RECT 0.048 380.544 5.082 380.640 ;
      RECT 0.048 381.312 5.082 381.408 ;
      RECT 0.048 382.080 5.082 382.176 ;
      RECT 0.048 382.848 5.082 382.944 ;
      RECT 0.048 383.616 5.082 383.712 ;
      RECT 0.048 384.384 5.082 384.480 ;
      RECT 0.048 385.152 5.082 385.248 ;
      RECT 0.048 385.920 5.082 386.016 ;
      RECT 0.048 386.688 5.082 386.784 ;
      RECT 0.048 387.456 5.082 387.552 ;
      RECT 0.048 388.224 5.082 388.320 ;
      RECT 0.048 388.992 5.082 389.088 ;
      RECT 0.048 389.760 5.082 389.856 ;
      RECT 0.048 390.528 5.082 390.624 ;
      RECT 0.048 391.296 5.082 391.392 ;
      RECT 0.048 392.064 5.082 392.160 ;
      RECT 0.048 392.832 5.082 392.928 ;
      RECT 0.048 393.600 5.082 393.696 ;
      RECT 0.048 394.368 5.082 394.464 ;
      RECT 0.048 395.136 5.082 395.232 ;
      RECT 0.048 395.904 5.082 396.000 ;
      RECT 0.048 396.672 5.082 396.768 ;
      RECT 0.048 397.440 5.082 397.536 ;
      RECT 0.048 398.208 5.082 398.304 ;
      RECT 0.048 398.976 5.082 399.072 ;
      RECT 0.048 399.744 5.082 399.840 ;
      RECT 0.048 400.512 5.082 400.608 ;
      RECT 0.048 401.280 5.082 401.376 ;
      RECT 0.048 402.048 5.082 402.144 ;
      RECT 0.048 402.816 5.082 402.912 ;
      RECT 0.048 403.584 5.082 403.680 ;
      RECT 0.048 404.352 5.082 404.448 ;
      RECT 0.048 405.120 5.082 405.216 ;
      RECT 0.048 405.888 5.082 405.984 ;
      RECT 0.048 406.656 5.082 406.752 ;
      RECT 0.048 407.424 5.082 407.520 ;
      RECT 0.048 408.192 5.082 408.288 ;
      RECT 0.048 408.960 5.082 409.056 ;
      RECT 0.048 409.728 5.082 409.824 ;
      RECT 0.048 410.496 5.082 410.592 ;
      RECT 0.048 411.264 5.082 411.360 ;
      RECT 0.048 412.032 5.082 412.128 ;
      RECT 0.048 412.800 5.082 412.896 ;
      RECT 0.048 413.568 5.082 413.664 ;
      RECT 0.048 414.336 5.082 414.432 ;
      RECT 0.048 415.104 5.082 415.200 ;
      RECT 0.048 415.872 5.082 415.968 ;
      RECT 0.048 416.640 5.082 416.736 ;
      RECT 0.048 417.408 5.082 417.504 ;
      RECT 0.048 418.176 5.082 418.272 ;
      RECT 0.048 418.944 5.082 419.040 ;
      RECT 0.048 419.712 5.082 419.808 ;
      RECT 0.048 420.480 5.082 420.576 ;
      RECT 0.048 421.248 5.082 421.344 ;
      RECT 0.048 422.016 5.082 422.112 ;
      RECT 0.048 422.784 5.082 422.880 ;
      RECT 0.048 423.552 5.082 423.648 ;
      RECT 0.048 424.320 5.082 424.416 ;
      RECT 0.048 425.088 5.082 425.184 ;
      RECT 0.048 425.856 5.082 425.952 ;
      RECT 0.048 426.624 5.082 426.720 ;
      RECT 0.048 427.392 5.082 427.488 ;
      RECT 0.048 428.160 5.082 428.256 ;
      RECT 0.048 428.928 5.082 429.024 ;
      RECT 0.048 429.696 5.082 429.792 ;
      RECT 0.048 430.464 5.082 430.560 ;
      RECT 0.048 431.232 5.082 431.328 ;
      RECT 0.048 432.000 5.082 432.096 ;
      RECT 0.048 432.768 5.082 432.864 ;
      RECT 0.048 433.536 5.082 433.632 ;
      RECT 0.048 434.304 5.082 434.400 ;
      RECT 0.048 435.072 5.082 435.168 ;
      RECT 0.048 435.840 5.082 435.936 ;
      RECT 0.048 436.608 5.082 436.704 ;
      RECT 0.048 437.376 5.082 437.472 ;
      RECT 0.048 438.144 5.082 438.240 ;
      RECT 0.048 438.912 5.082 439.008 ;
      RECT 0.048 439.680 5.082 439.776 ;
      RECT 0.048 440.448 5.082 440.544 ;
      RECT 0.048 441.216 5.082 441.312 ;
      RECT 0.048 441.984 5.082 442.080 ;
      RECT 0.048 442.752 5.082 442.848 ;
      RECT 0.048 443.520 5.082 443.616 ;
      RECT 0.048 444.288 5.082 444.384 ;
      RECT 0.048 445.056 5.082 445.152 ;
      RECT 0.048 445.824 5.082 445.920 ;
      RECT 0.048 446.592 5.082 446.688 ;
      RECT 0.048 447.360 5.082 447.456 ;
      RECT 0.048 448.128 5.082 448.224 ;
      RECT 0.048 448.896 5.082 448.992 ;
      RECT 0.048 449.664 5.082 449.760 ;
      RECT 0.048 450.432 5.082 450.528 ;
      RECT 0.048 451.200 5.082 451.296 ;
      RECT 0.048 451.968 5.082 452.064 ;
      RECT 0.048 452.736 5.082 452.832 ;
      RECT 0.048 453.504 5.082 453.600 ;
      RECT 0.048 454.272 5.082 454.368 ;
      RECT 0.048 455.040 5.082 455.136 ;
      RECT 0.048 455.808 5.082 455.904 ;
      RECT 0.048 456.576 5.082 456.672 ;
      RECT 0.048 457.344 5.082 457.440 ;
      RECT 0.048 458.112 5.082 458.208 ;
      RECT 0.048 458.880 5.082 458.976 ;
      RECT 0.048 459.648 5.082 459.744 ;
      RECT 0.048 460.416 5.082 460.512 ;
      RECT 0.048 461.184 5.082 461.280 ;
      RECT 0.048 461.952 5.082 462.048 ;
      RECT 0.048 462.720 5.082 462.816 ;
      RECT 0.048 463.488 5.082 463.584 ;
      RECT 0.048 464.256 5.082 464.352 ;
      RECT 0.048 465.024 5.082 465.120 ;
      RECT 0.048 465.792 5.082 465.888 ;
      RECT 0.048 466.560 5.082 466.656 ;
      RECT 0.048 467.328 5.082 467.424 ;
      RECT 0.048 468.096 5.082 468.192 ;
      RECT 0.048 468.864 5.082 468.960 ;
      RECT 0.048 469.632 5.082 469.728 ;
      RECT 0.048 470.400 5.082 470.496 ;
      RECT 0.048 471.168 5.082 471.264 ;
      RECT 0.048 471.936 5.082 472.032 ;
      RECT 0.048 472.704 5.082 472.800 ;
      RECT 0.048 473.472 5.082 473.568 ;
      RECT 0.048 474.240 5.082 474.336 ;
      RECT 0.048 475.008 5.082 475.104 ;
      RECT 0.048 475.776 5.082 475.872 ;
      RECT 0.048 476.544 5.082 476.640 ;
      RECT 0.048 477.312 5.082 477.408 ;
      RECT 0.048 478.080 5.082 478.176 ;
      RECT 0.048 478.848 5.082 478.944 ;
      RECT 0.048 479.616 5.082 479.712 ;
      RECT 0.048 480.384 5.082 480.480 ;
      RECT 0.048 481.152 5.082 481.248 ;
      RECT 0.048 481.920 5.082 482.016 ;
      RECT 0.048 482.688 5.082 482.784 ;
      RECT 0.048 483.456 5.082 483.552 ;
      RECT 0.048 484.224 5.082 484.320 ;
      RECT 0.048 484.992 5.082 485.088 ;
      RECT 0.048 485.760 5.082 485.856 ;
      RECT 0.048 486.528 5.082 486.624 ;
      RECT 0.048 487.296 5.082 487.392 ;
      RECT 0.048 488.064 5.082 488.160 ;
      RECT 0.048 488.832 5.082 488.928 ;
      RECT 0.048 489.600 5.082 489.696 ;
      RECT 0.048 490.368 5.082 490.464 ;
      RECT 0.048 491.136 5.082 491.232 ;
      RECT 0.048 491.904 5.082 492.000 ;
      RECT 0.048 492.672 5.082 492.768 ;
      RECT 0.048 493.440 5.082 493.536 ;
      RECT 0.048 494.208 5.082 494.304 ;
      RECT 0.048 494.976 5.082 495.072 ;
      RECT 0.048 495.744 5.082 495.840 ;
      RECT 0.048 496.512 5.082 496.608 ;
      RECT 0.048 497.280 5.082 497.376 ;
      RECT 0.048 498.048 5.082 498.144 ;
      RECT 0.048 498.816 5.082 498.912 ;
      RECT 0.048 499.584 5.082 499.680 ;
      RECT 0.048 500.352 5.082 500.448 ;
      RECT 0.048 501.120 5.082 501.216 ;
      RECT 0.048 501.888 5.082 501.984 ;
      RECT 0.048 502.656 5.082 502.752 ;
      RECT 0.048 503.424 5.082 503.520 ;
      RECT 0.048 504.192 5.082 504.288 ;
      RECT 0.048 504.960 5.082 505.056 ;
      RECT 0.048 505.728 5.082 505.824 ;
      RECT 0.048 506.496 5.082 506.592 ;
      RECT 0.048 507.264 5.082 507.360 ;
      RECT 0.048 508.032 5.082 508.128 ;
      RECT 0.048 508.800 5.082 508.896 ;
      RECT 0.048 509.568 5.082 509.664 ;
      RECT 0.048 510.336 5.082 510.432 ;
      RECT 0.048 511.104 5.082 511.200 ;
      RECT 0.048 511.872 5.082 511.968 ;
      RECT 0.048 512.640 5.082 512.736 ;
      RECT 0.048 513.408 5.082 513.504 ;
      RECT 0.048 514.176 5.082 514.272 ;
      RECT 0.048 514.944 5.082 515.040 ;
      RECT 0.048 515.712 5.082 515.808 ;
      RECT 0.048 516.480 5.082 516.576 ;
      RECT 0.048 517.248 5.082 517.344 ;
      RECT 0.048 518.016 5.082 518.112 ;
      RECT 0.048 518.784 5.082 518.880 ;
      RECT 0.048 519.552 5.082 519.648 ;
      RECT 0.048 520.320 5.082 520.416 ;
      RECT 0.048 521.088 5.082 521.184 ;
      RECT 0.048 521.856 5.082 521.952 ;
      RECT 0.048 522.624 5.082 522.720 ;
      RECT 0.048 523.392 5.082 523.488 ;
      RECT 0.048 524.160 5.082 524.256 ;
      RECT 0.048 524.928 5.082 525.024 ;
      RECT 0.048 525.696 5.082 525.792 ;
      RECT 0.048 526.464 5.082 526.560 ;
      RECT 0.048 527.232 5.082 527.328 ;
      RECT 0.048 528.000 5.082 528.096 ;
      RECT 0.048 528.768 5.082 528.864 ;
      RECT 0.048 529.536 5.082 529.632 ;
      RECT 0.048 530.304 5.082 530.400 ;
      RECT 0.048 531.072 5.082 531.168 ;
      RECT 0.048 531.840 5.082 531.936 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 5.130 532.000 ;
    LAYER M2 ;
    RECT 0 0 5.130 532.000 ;
    LAYER M3 ;
    RECT 0 0 5.130 532.000 ;
    LAYER M4 ;
    RECT 0.1 0 5.030 532.000 ;
  END
END fakeram7_2048x39

END LIBRARY
