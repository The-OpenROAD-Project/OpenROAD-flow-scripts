../../nangate45/lef/fakeram45_256x16.lef