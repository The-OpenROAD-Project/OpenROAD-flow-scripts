VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 2000 ;
END UNITS
MACRO or1200_spram4
  FOREIGN or1200_spram4 0 0 ;
  CLASS BLOCK ;
  SIZE 293.635 BY 410.29 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  2.94 402.7 283.34 404.1 ;
        RECT  2.94 362.7 283.34 364.1 ;
        RECT  2.94 322.7 283.34 324.1 ;
        RECT  2.94 282.7 283.34 284.1 ;
        RECT  2.94 242.7 283.34 244.1 ;
        RECT  2.94 202.7 283.34 204.1 ;
        RECT  2.94 162.7 283.34 164.1 ;
        RECT  2.94 122.7 283.34 124.1 ;
        RECT  2.94 82.7 283.34 84.1 ;
        RECT  2.94 42.7 283.34 44.1 ;
        RECT  2.94 2.7 283.34 4.1 ;
      LAYER metal4 ;
        RECT  283.04 1.33 283.24 407.47 ;
        RECT  227.04 1.33 227.24 407.47 ;
        RECT  171.04 1.33 171.24 407.47 ;
        RECT  115.04 1.33 115.24 407.47 ;
        RECT  59.04 1.33 59.24 407.47 ;
        RECT  3.04 1.33 3.24 407.47 ;
      LAYER metal1 ;
        RECT  1.14 407.35 292.6 407.45 ;
        RECT  1.14 404.55 292.6 404.65 ;
        RECT  1.14 401.75 292.6 401.85 ;
        RECT  1.14 398.95 292.6 399.05 ;
        RECT  1.14 396.15 292.6 396.25 ;
        RECT  1.14 393.35 292.6 393.45 ;
        RECT  1.14 390.55 292.6 390.65 ;
        RECT  1.14 387.75 292.6 387.85 ;
        RECT  1.14 384.95 292.6 385.05 ;
        RECT  1.14 382.15 292.6 382.25 ;
        RECT  1.14 379.35 292.6 379.45 ;
        RECT  1.14 376.55 292.6 376.65 ;
        RECT  1.14 373.75 292.6 373.85 ;
        RECT  1.14 370.95 292.6 371.05 ;
        RECT  1.14 368.15 292.6 368.25 ;
        RECT  1.14 365.35 292.6 365.45 ;
        RECT  1.14 362.55 292.6 362.65 ;
        RECT  1.14 359.75 292.6 359.85 ;
        RECT  1.14 356.95 292.6 357.05 ;
        RECT  1.14 354.15 292.6 354.25 ;
        RECT  1.14 351.35 292.6 351.45 ;
        RECT  1.14 348.55 292.6 348.65 ;
        RECT  1.14 345.75 292.6 345.85 ;
        RECT  1.14 342.95 292.6 343.05 ;
        RECT  1.14 340.15 292.6 340.25 ;
        RECT  1.14 337.35 292.6 337.45 ;
        RECT  1.14 334.55 292.6 334.65 ;
        RECT  1.14 331.75 292.6 331.85 ;
        RECT  1.14 328.95 292.6 329.05 ;
        RECT  1.14 326.15 292.6 326.25 ;
        RECT  1.14 323.35 292.6 323.45 ;
        RECT  1.14 320.55 292.6 320.65 ;
        RECT  1.14 317.75 292.6 317.85 ;
        RECT  1.14 314.95 292.6 315.05 ;
        RECT  1.14 312.15 292.6 312.25 ;
        RECT  1.14 309.35 292.6 309.45 ;
        RECT  1.14 306.55 292.6 306.65 ;
        RECT  1.14 303.75 292.6 303.85 ;
        RECT  1.14 300.95 292.6 301.05 ;
        RECT  1.14 298.15 292.6 298.25 ;
        RECT  1.14 295.35 292.6 295.45 ;
        RECT  1.14 292.55 292.6 292.65 ;
        RECT  1.14 289.75 292.6 289.85 ;
        RECT  1.14 286.95 292.6 287.05 ;
        RECT  1.14 284.15 292.6 284.25 ;
        RECT  1.14 281.35 292.6 281.45 ;
        RECT  1.14 278.55 292.6 278.65 ;
        RECT  1.14 275.75 292.6 275.85 ;
        RECT  1.14 272.95 292.6 273.05 ;
        RECT  1.14 270.15 292.6 270.25 ;
        RECT  1.14 267.35 292.6 267.45 ;
        RECT  1.14 264.55 292.6 264.65 ;
        RECT  1.14 261.75 292.6 261.85 ;
        RECT  1.14 258.95 292.6 259.05 ;
        RECT  1.14 256.15 292.6 256.25 ;
        RECT  1.14 253.35 292.6 253.45 ;
        RECT  1.14 250.55 292.6 250.65 ;
        RECT  1.14 247.75 292.6 247.85 ;
        RECT  1.14 244.95 292.6 245.05 ;
        RECT  1.14 242.15 292.6 242.25 ;
        RECT  1.14 239.35 292.6 239.45 ;
        RECT  1.14 236.55 292.6 236.65 ;
        RECT  1.14 233.75 292.6 233.85 ;
        RECT  1.14 230.95 292.6 231.05 ;
        RECT  1.14 228.15 292.6 228.25 ;
        RECT  1.14 225.35 292.6 225.45 ;
        RECT  1.14 222.55 292.6 222.65 ;
        RECT  1.14 219.75 292.6 219.85 ;
        RECT  1.14 216.95 292.6 217.05 ;
        RECT  1.14 214.15 292.6 214.25 ;
        RECT  1.14 211.35 292.6 211.45 ;
        RECT  1.14 208.55 292.6 208.65 ;
        RECT  1.14 205.75 292.6 205.85 ;
        RECT  1.14 202.95 292.6 203.05 ;
        RECT  1.14 200.15 292.6 200.25 ;
        RECT  1.14 197.35 292.6 197.45 ;
        RECT  1.14 194.55 292.6 194.65 ;
        RECT  1.14 191.75 292.6 191.85 ;
        RECT  1.14 188.95 292.6 189.05 ;
        RECT  1.14 186.15 292.6 186.25 ;
        RECT  1.14 183.35 292.6 183.45 ;
        RECT  1.14 180.55 292.6 180.65 ;
        RECT  1.14 177.75 292.6 177.85 ;
        RECT  1.14 174.95 292.6 175.05 ;
        RECT  1.14 172.15 292.6 172.25 ;
        RECT  1.14 169.35 292.6 169.45 ;
        RECT  1.14 166.55 292.6 166.65 ;
        RECT  1.14 163.75 292.6 163.85 ;
        RECT  1.14 160.95 292.6 161.05 ;
        RECT  1.14 158.15 292.6 158.25 ;
        RECT  1.14 155.35 292.6 155.45 ;
        RECT  1.14 152.55 292.6 152.65 ;
        RECT  1.14 149.75 292.6 149.85 ;
        RECT  1.14 146.95 292.6 147.05 ;
        RECT  1.14 144.15 292.6 144.25 ;
        RECT  1.14 141.35 292.6 141.45 ;
        RECT  1.14 138.55 292.6 138.65 ;
        RECT  1.14 135.75 292.6 135.85 ;
        RECT  1.14 132.95 292.6 133.05 ;
        RECT  1.14 130.15 292.6 130.25 ;
        RECT  1.14 127.35 292.6 127.45 ;
        RECT  1.14 124.55 292.6 124.65 ;
        RECT  1.14 121.75 292.6 121.85 ;
        RECT  1.14 118.95 292.6 119.05 ;
        RECT  1.14 116.15 292.6 116.25 ;
        RECT  1.14 113.35 292.6 113.45 ;
        RECT  1.14 110.55 292.6 110.65 ;
        RECT  1.14 107.75 292.6 107.85 ;
        RECT  1.14 104.95 292.6 105.05 ;
        RECT  1.14 102.15 292.6 102.25 ;
        RECT  1.14 99.35 292.6 99.45 ;
        RECT  1.14 96.55 292.6 96.65 ;
        RECT  1.14 93.75 292.6 93.85 ;
        RECT  1.14 90.95 292.6 91.05 ;
        RECT  1.14 88.15 292.6 88.25 ;
        RECT  1.14 85.35 292.6 85.45 ;
        RECT  1.14 82.55 292.6 82.65 ;
        RECT  1.14 79.75 292.6 79.85 ;
        RECT  1.14 76.95 292.6 77.05 ;
        RECT  1.14 74.15 292.6 74.25 ;
        RECT  1.14 71.35 292.6 71.45 ;
        RECT  1.14 68.55 292.6 68.65 ;
        RECT  1.14 65.75 292.6 65.85 ;
        RECT  1.14 62.95 292.6 63.05 ;
        RECT  1.14 60.15 292.6 60.25 ;
        RECT  1.14 57.35 292.6 57.45 ;
        RECT  1.14 54.55 292.6 54.65 ;
        RECT  1.14 51.75 292.6 51.85 ;
        RECT  1.14 48.95 292.6 49.05 ;
        RECT  1.14 46.15 292.6 46.25 ;
        RECT  1.14 43.35 292.6 43.45 ;
        RECT  1.14 40.55 292.6 40.65 ;
        RECT  1.14 37.75 292.6 37.85 ;
        RECT  1.14 34.95 292.6 35.05 ;
        RECT  1.14 32.15 292.6 32.25 ;
        RECT  1.14 29.35 292.6 29.45 ;
        RECT  1.14 26.55 292.6 26.65 ;
        RECT  1.14 23.75 292.6 23.85 ;
        RECT  1.14 20.95 292.6 21.05 ;
        RECT  1.14 18.15 292.6 18.25 ;
        RECT  1.14 15.35 292.6 15.45 ;
        RECT  1.14 12.55 292.6 12.65 ;
        RECT  1.14 9.75 292.6 9.85 ;
        RECT  1.14 6.95 292.6 7.05 ;
        RECT  1.14 4.15 292.6 4.25 ;
        RECT  1.14 1.35 292.6 1.45 ;
      VIA 283.14 403.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 403.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 403.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 363.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 363.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 363.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 283.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 283.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 403.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 403.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 403.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 363.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 363.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 363.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 227.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 227.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 227.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 403.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 403.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 403.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 363.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 363.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 363.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 171.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 171.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 171.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 403.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 403.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 403.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 363.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 363.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 363.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 115.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 115.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 115.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 403.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 403.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 403.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 363.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 363.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 363.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 59.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 59.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 59.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 403.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 403.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 403.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 363.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 363.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 363.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 323.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 323.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 323.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 283.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 283.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 283.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 243.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 243.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 243.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 203.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 203.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 203.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 163.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 163.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 163.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 123.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 123.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 123.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 83.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 83.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 83.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 43.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 43.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 43.4 via4_5_400_2800_5_1_600_600 ;
      VIA 3.14 3.4 via6_7_400_2800_4_1_600_600 ;
      VIA 3.14 3.4 via5_6_400_2800_5_1_600_600 ;
      VIA 3.14 3.4 via4_5_400_2800_5_1_600_600 ;
      VIA 283.14 407.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 407.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 407.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 404.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 404.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 404.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 401.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 401.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 401.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 399 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 399 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 399 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 396.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 396.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 396.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 393.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 393.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 393.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 390.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 390.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 390.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 387.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 387.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 387.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 385 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 385 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 385 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 382.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 382.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 382.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 379.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 379.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 379.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 376.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 376.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 376.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 373.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 373.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 373.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 371 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 371 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 371 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 368.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 368.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 368.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 365.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 365.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 365.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 362.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 362.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 362.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 359.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 359.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 359.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 357 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 357 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 357 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 354.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 354.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 354.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 351.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 351.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 351.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 348.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 348.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 348.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 345.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 345.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 345.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 343 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 343 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 343 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 340.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 340.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 340.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 283.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 283.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 283.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 407.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 407.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 407.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 404.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 404.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 404.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 401.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 401.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 401.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 399 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 399 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 399 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 396.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 396.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 396.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 393.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 393.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 393.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 390.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 390.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 390.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 387.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 387.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 387.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 385 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 385 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 385 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 382.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 382.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 382.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 379.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 379.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 379.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 376.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 376.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 376.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 373.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 373.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 373.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 371 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 371 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 371 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 368.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 368.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 368.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 365.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 365.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 365.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 362.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 362.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 362.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 359.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 359.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 359.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 357 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 357 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 357 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 354.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 354.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 354.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 351.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 351.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 351.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 348.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 348.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 348.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 345.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 345.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 345.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 343 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 343 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 343 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 340.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 340.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 340.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 227.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 227.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 227.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 407.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 407.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 407.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 404.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 404.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 404.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 401.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 401.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 401.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 399 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 399 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 399 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 396.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 396.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 396.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 393.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 393.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 393.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 390.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 390.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 390.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 387.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 387.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 387.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 385 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 385 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 385 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 382.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 382.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 382.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 379.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 379.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 379.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 376.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 376.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 376.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 373.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 373.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 373.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 371 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 371 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 371 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 368.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 368.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 368.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 365.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 365.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 365.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 362.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 362.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 362.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 359.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 359.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 359.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 357 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 357 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 357 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 354.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 354.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 354.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 351.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 351.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 351.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 348.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 348.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 348.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 345.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 345.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 345.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 343 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 343 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 343 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 340.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 340.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 340.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 171.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 171.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 171.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 407.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 407.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 407.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 404.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 404.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 404.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 401.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 401.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 401.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 399 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 399 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 399 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 396.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 396.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 396.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 393.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 393.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 393.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 390.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 390.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 390.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 387.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 387.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 387.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 385 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 385 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 385 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 382.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 382.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 382.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 379.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 379.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 379.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 376.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 376.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 376.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 373.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 373.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 373.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 371 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 371 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 371 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 368.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 368.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 368.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 365.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 365.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 365.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 362.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 362.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 362.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 359.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 359.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 359.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 357 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 357 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 357 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 354.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 354.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 354.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 351.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 351.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 351.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 348.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 348.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 348.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 345.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 345.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 345.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 343 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 343 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 343 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 340.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 340.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 340.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 115.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 115.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 115.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 407.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 407.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 407.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 404.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 404.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 404.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 401.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 401.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 401.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 399 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 399 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 399 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 396.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 396.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 396.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 393.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 393.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 393.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 390.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 390.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 390.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 387.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 387.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 387.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 385 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 385 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 385 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 382.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 382.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 382.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 379.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 379.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 379.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 376.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 376.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 376.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 373.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 373.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 373.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 371 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 371 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 371 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 368.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 368.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 368.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 365.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 365.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 365.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 362.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 362.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 362.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 359.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 359.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 359.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 357 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 357 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 357 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 354.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 354.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 354.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 351.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 351.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 351.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 348.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 348.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 348.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 345.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 345.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 345.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 343 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 343 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 343 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 340.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 340.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 340.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 59.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 59.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 59.14 1.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 407.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 407.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 407.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 404.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 404.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 404.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 401.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 401.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 401.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 399 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 399 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 399 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 396.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 396.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 396.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 393.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 393.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 393.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 390.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 390.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 390.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 387.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 387.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 387.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 385 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 385 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 385 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 382.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 382.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 382.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 379.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 379.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 379.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 376.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 376.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 376.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 373.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 373.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 373.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 371 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 371 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 371 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 368.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 368.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 368.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 365.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 365.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 365.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 362.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 362.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 362.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 359.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 359.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 359.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 357 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 357 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 357 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 354.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 354.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 354.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 351.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 351.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 351.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 348.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 348.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 348.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 345.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 345.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 345.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 343 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 343 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 343 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 340.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 340.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 340.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 337.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 337.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 337.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 334.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 334.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 334.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 331.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 331.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 331.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 329 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 329 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 329 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 326.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 326.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 326.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 323.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 323.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 323.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 320.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 320.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 320.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 317.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 317.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 317.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 315 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 315 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 315 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 312.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 312.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 312.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 309.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 309.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 309.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 306.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 306.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 306.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 303.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 303.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 303.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 301 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 301 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 301 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 298.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 298.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 298.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 295.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 295.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 295.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 292.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 292.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 292.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 289.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 289.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 289.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 287 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 287 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 287 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 284.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 284.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 284.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 281.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 281.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 281.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 278.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 278.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 278.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 275.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 275.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 275.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 273 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 273 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 273 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 270.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 270.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 270.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 267.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 267.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 267.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 264.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 264.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 264.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 261.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 261.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 261.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 259 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 259 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 259 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 256.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 256.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 256.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 253.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 253.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 253.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 250.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 250.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 250.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 247.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 247.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 247.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 245 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 245 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 245 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 242.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 242.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 242.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 239.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 239.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 239.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 236.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 236.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 236.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 233.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 233.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 233.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 231 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 231 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 231 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 228.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 228.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 228.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 225.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 225.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 225.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 222.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 222.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 222.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 219.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 219.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 219.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 217 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 217 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 217 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 214.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 214.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 214.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 211.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 211.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 211.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 208.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 208.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 208.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 205.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 205.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 205.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 203 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 203 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 203 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 200.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 200.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 200.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 197.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 197.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 197.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 194.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 194.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 194.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 191.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 191.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 191.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 189 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 189 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 189 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 186.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 186.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 186.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 183.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 183.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 183.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 180.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 180.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 180.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 177.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 177.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 177.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 175 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 175 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 175 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 172.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 172.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 172.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 169.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 169.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 169.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 166.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 166.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 166.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 163.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 163.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 163.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 161 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 161 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 161 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 158.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 158.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 158.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 155.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 155.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 155.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 152.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 152.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 152.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 149.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 149.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 149.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 147 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 147 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 147 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 144.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 144.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 144.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 141.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 141.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 141.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 138.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 138.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 138.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 135.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 135.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 135.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 133 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 133 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 133 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 130.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 130.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 130.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 127.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 127.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 127.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 124.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 124.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 124.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 121.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 121.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 121.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 119 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 119 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 119 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 116.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 116.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 116.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 113.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 113.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 113.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 110.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 110.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 110.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 107.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 107.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 107.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 105 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 105 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 105 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 102.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 102.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 102.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 99.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 99.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 99.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 96.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 96.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 96.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 93.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 93.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 93.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 91 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 91 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 91 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 88.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 88.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 88.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 85.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 85.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 85.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 82.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 82.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 82.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 79.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 79.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 79.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 77 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 77 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 77 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 74.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 74.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 74.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 71.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 71.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 71.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 68.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 68.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 68.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 65.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 65.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 65.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 63 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 63 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 63 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 60.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 60.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 60.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 57.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 57.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 57.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 54.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 54.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 54.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 51.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 51.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 51.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 49 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 49 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 49 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 46.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 46.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 46.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 43.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 43.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 43.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 40.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 40.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 40.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 37.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 37.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 37.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 35 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 35 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 35 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 32.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 32.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 32.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 29.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 29.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 29.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 26.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 26.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 26.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 23.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 23.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 23.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 21 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 21 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 21 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 18.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 18.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 18.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 15.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 15.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 15.4 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 12.6 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 12.6 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 12.6 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 9.8 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 9.8 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 9.8 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 7 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 7 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 7 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 4.2 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 4.2 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 4.2 via1_2_400_200_1_1_300_300 ;
      VIA 3.14 1.4 via3_4_400_200_1_1_320_320 ;
      VIA 3.14 1.4 via2_3_400_200_1_1_320_320 ;
      VIA 3.14 1.4 via1_2_400_200_1_1_300_300 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER metal7 ;
        RECT  30.94 382.7 255.34 384.1 ;
        RECT  30.94 342.7 255.34 344.1 ;
        RECT  30.94 302.7 255.34 304.1 ;
        RECT  30.94 262.7 255.34 264.1 ;
        RECT  30.94 222.7 255.34 224.1 ;
        RECT  30.94 182.7 255.34 184.1 ;
        RECT  30.94 142.7 255.34 144.1 ;
        RECT  30.94 102.7 255.34 104.1 ;
        RECT  30.94 62.7 255.34 64.1 ;
        RECT  30.94 22.7 255.34 24.1 ;
      LAYER metal4 ;
        RECT  255.04 2.73 255.24 408.87 ;
        RECT  199.04 2.73 199.24 408.87 ;
        RECT  143.04 2.73 143.24 408.87 ;
        RECT  87.04 2.73 87.24 408.87 ;
        RECT  31.04 2.73 31.24 408.87 ;
      LAYER metal1 ;
        RECT  1.14 408.75 292.6 408.85 ;
        RECT  1.14 405.95 292.6 406.05 ;
        RECT  1.14 403.15 292.6 403.25 ;
        RECT  1.14 400.35 292.6 400.45 ;
        RECT  1.14 397.55 292.6 397.65 ;
        RECT  1.14 394.75 292.6 394.85 ;
        RECT  1.14 391.95 292.6 392.05 ;
        RECT  1.14 389.15 292.6 389.25 ;
        RECT  1.14 386.35 292.6 386.45 ;
        RECT  1.14 383.55 292.6 383.65 ;
        RECT  1.14 380.75 292.6 380.85 ;
        RECT  1.14 377.95 292.6 378.05 ;
        RECT  1.14 375.15 292.6 375.25 ;
        RECT  1.14 372.35 292.6 372.45 ;
        RECT  1.14 369.55 292.6 369.65 ;
        RECT  1.14 366.75 292.6 366.85 ;
        RECT  1.14 363.95 292.6 364.05 ;
        RECT  1.14 361.15 292.6 361.25 ;
        RECT  1.14 358.35 292.6 358.45 ;
        RECT  1.14 355.55 292.6 355.65 ;
        RECT  1.14 352.75 292.6 352.85 ;
        RECT  1.14 349.95 292.6 350.05 ;
        RECT  1.14 347.15 292.6 347.25 ;
        RECT  1.14 344.35 292.6 344.45 ;
        RECT  1.14 341.55 292.6 341.65 ;
        RECT  1.14 338.75 292.6 338.85 ;
        RECT  1.14 335.95 292.6 336.05 ;
        RECT  1.14 333.15 292.6 333.25 ;
        RECT  1.14 330.35 292.6 330.45 ;
        RECT  1.14 327.55 292.6 327.65 ;
        RECT  1.14 324.75 292.6 324.85 ;
        RECT  1.14 321.95 292.6 322.05 ;
        RECT  1.14 319.15 292.6 319.25 ;
        RECT  1.14 316.35 292.6 316.45 ;
        RECT  1.14 313.55 292.6 313.65 ;
        RECT  1.14 310.75 292.6 310.85 ;
        RECT  1.14 307.95 292.6 308.05 ;
        RECT  1.14 305.15 292.6 305.25 ;
        RECT  1.14 302.35 292.6 302.45 ;
        RECT  1.14 299.55 292.6 299.65 ;
        RECT  1.14 296.75 292.6 296.85 ;
        RECT  1.14 293.95 292.6 294.05 ;
        RECT  1.14 291.15 292.6 291.25 ;
        RECT  1.14 288.35 292.6 288.45 ;
        RECT  1.14 285.55 292.6 285.65 ;
        RECT  1.14 282.75 292.6 282.85 ;
        RECT  1.14 279.95 292.6 280.05 ;
        RECT  1.14 277.15 292.6 277.25 ;
        RECT  1.14 274.35 292.6 274.45 ;
        RECT  1.14 271.55 292.6 271.65 ;
        RECT  1.14 268.75 292.6 268.85 ;
        RECT  1.14 265.95 292.6 266.05 ;
        RECT  1.14 263.15 292.6 263.25 ;
        RECT  1.14 260.35 292.6 260.45 ;
        RECT  1.14 257.55 292.6 257.65 ;
        RECT  1.14 254.75 292.6 254.85 ;
        RECT  1.14 251.95 292.6 252.05 ;
        RECT  1.14 249.15 292.6 249.25 ;
        RECT  1.14 246.35 292.6 246.45 ;
        RECT  1.14 243.55 292.6 243.65 ;
        RECT  1.14 240.75 292.6 240.85 ;
        RECT  1.14 237.95 292.6 238.05 ;
        RECT  1.14 235.15 292.6 235.25 ;
        RECT  1.14 232.35 292.6 232.45 ;
        RECT  1.14 229.55 292.6 229.65 ;
        RECT  1.14 226.75 292.6 226.85 ;
        RECT  1.14 223.95 292.6 224.05 ;
        RECT  1.14 221.15 292.6 221.25 ;
        RECT  1.14 218.35 292.6 218.45 ;
        RECT  1.14 215.55 292.6 215.65 ;
        RECT  1.14 212.75 292.6 212.85 ;
        RECT  1.14 209.95 292.6 210.05 ;
        RECT  1.14 207.15 292.6 207.25 ;
        RECT  1.14 204.35 292.6 204.45 ;
        RECT  1.14 201.55 292.6 201.65 ;
        RECT  1.14 198.75 292.6 198.85 ;
        RECT  1.14 195.95 292.6 196.05 ;
        RECT  1.14 193.15 292.6 193.25 ;
        RECT  1.14 190.35 292.6 190.45 ;
        RECT  1.14 187.55 292.6 187.65 ;
        RECT  1.14 184.75 292.6 184.85 ;
        RECT  1.14 181.95 292.6 182.05 ;
        RECT  1.14 179.15 292.6 179.25 ;
        RECT  1.14 176.35 292.6 176.45 ;
        RECT  1.14 173.55 292.6 173.65 ;
        RECT  1.14 170.75 292.6 170.85 ;
        RECT  1.14 167.95 292.6 168.05 ;
        RECT  1.14 165.15 292.6 165.25 ;
        RECT  1.14 162.35 292.6 162.45 ;
        RECT  1.14 159.55 292.6 159.65 ;
        RECT  1.14 156.75 292.6 156.85 ;
        RECT  1.14 153.95 292.6 154.05 ;
        RECT  1.14 151.15 292.6 151.25 ;
        RECT  1.14 148.35 292.6 148.45 ;
        RECT  1.14 145.55 292.6 145.65 ;
        RECT  1.14 142.75 292.6 142.85 ;
        RECT  1.14 139.95 292.6 140.05 ;
        RECT  1.14 137.15 292.6 137.25 ;
        RECT  1.14 134.35 292.6 134.45 ;
        RECT  1.14 131.55 292.6 131.65 ;
        RECT  1.14 128.75 292.6 128.85 ;
        RECT  1.14 125.95 292.6 126.05 ;
        RECT  1.14 123.15 292.6 123.25 ;
        RECT  1.14 120.35 292.6 120.45 ;
        RECT  1.14 117.55 292.6 117.65 ;
        RECT  1.14 114.75 292.6 114.85 ;
        RECT  1.14 111.95 292.6 112.05 ;
        RECT  1.14 109.15 292.6 109.25 ;
        RECT  1.14 106.35 292.6 106.45 ;
        RECT  1.14 103.55 292.6 103.65 ;
        RECT  1.14 100.75 292.6 100.85 ;
        RECT  1.14 97.95 292.6 98.05 ;
        RECT  1.14 95.15 292.6 95.25 ;
        RECT  1.14 92.35 292.6 92.45 ;
        RECT  1.14 89.55 292.6 89.65 ;
        RECT  1.14 86.75 292.6 86.85 ;
        RECT  1.14 83.95 292.6 84.05 ;
        RECT  1.14 81.15 292.6 81.25 ;
        RECT  1.14 78.35 292.6 78.45 ;
        RECT  1.14 75.55 292.6 75.65 ;
        RECT  1.14 72.75 292.6 72.85 ;
        RECT  1.14 69.95 292.6 70.05 ;
        RECT  1.14 67.15 292.6 67.25 ;
        RECT  1.14 64.35 292.6 64.45 ;
        RECT  1.14 61.55 292.6 61.65 ;
        RECT  1.14 58.75 292.6 58.85 ;
        RECT  1.14 55.95 292.6 56.05 ;
        RECT  1.14 53.15 292.6 53.25 ;
        RECT  1.14 50.35 292.6 50.45 ;
        RECT  1.14 47.55 292.6 47.65 ;
        RECT  1.14 44.75 292.6 44.85 ;
        RECT  1.14 41.95 292.6 42.05 ;
        RECT  1.14 39.15 292.6 39.25 ;
        RECT  1.14 36.35 292.6 36.45 ;
        RECT  1.14 33.55 292.6 33.65 ;
        RECT  1.14 30.75 292.6 30.85 ;
        RECT  1.14 27.95 292.6 28.05 ;
        RECT  1.14 25.15 292.6 25.25 ;
        RECT  1.14 22.35 292.6 22.45 ;
        RECT  1.14 19.55 292.6 19.65 ;
        RECT  1.14 16.75 292.6 16.85 ;
        RECT  1.14 13.95 292.6 14.05 ;
        RECT  1.14 11.15 292.6 11.25 ;
        RECT  1.14 8.35 292.6 8.45 ;
        RECT  1.14 5.55 292.6 5.65 ;
        RECT  1.14 2.75 292.6 2.85 ;
      VIA 255.14 383.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 383.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 383.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 343.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 343.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 343.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 255.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 255.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 383.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 383.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 383.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 343.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 343.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 343.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 199.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 199.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 199.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 383.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 383.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 383.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 343.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 343.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 343.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 143.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 143.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 143.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 383.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 383.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 383.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 343.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 343.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 343.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 87.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 87.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 87.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 383.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 383.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 383.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 343.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 343.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 343.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 303.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 303.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 303.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 263.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 263.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 263.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 223.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 223.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 223.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 183.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 183.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 183.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 143.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 143.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 143.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 103.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 103.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 103.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 63.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 63.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 63.4 via4_5_400_2800_5_1_600_600 ;
      VIA 31.14 23.4 via6_7_400_2800_4_1_600_600 ;
      VIA 31.14 23.4 via5_6_400_2800_5_1_600_600 ;
      VIA 31.14 23.4 via4_5_400_2800_5_1_600_600 ;
      VIA 255.14 408.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 408.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 408.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 406 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 406 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 406 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 403.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 403.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 403.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 400.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 400.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 400.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 397.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 397.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 397.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 394.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 394.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 394.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 392 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 392 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 392 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 389.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 389.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 389.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 386.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 386.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 386.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 383.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 383.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 383.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 380.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 380.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 380.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 378 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 378 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 378 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 375.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 375.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 375.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 372.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 372.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 372.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 369.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 369.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 369.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 366.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 366.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 366.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 364 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 364 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 364 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 361.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 361.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 361.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 358.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 358.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 358.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 355.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 355.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 355.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 352.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 352.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 352.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 350 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 350 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 350 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 347.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 347.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 347.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 344.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 344.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 344.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 341.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 341.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 341.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 255.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 255.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 255.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 408.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 408.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 408.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 406 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 406 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 406 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 403.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 403.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 403.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 400.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 400.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 400.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 397.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 397.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 397.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 394.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 394.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 394.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 392 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 392 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 392 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 389.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 389.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 389.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 386.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 386.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 386.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 383.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 383.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 383.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 380.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 380.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 380.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 378 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 378 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 378 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 375.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 375.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 375.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 372.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 372.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 372.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 369.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 369.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 369.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 366.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 366.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 366.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 364 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 364 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 364 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 361.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 361.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 361.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 358.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 358.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 358.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 355.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 355.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 355.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 352.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 352.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 352.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 350 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 350 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 350 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 347.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 347.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 347.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 344.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 344.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 344.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 341.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 341.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 341.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 199.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 199.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 199.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 408.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 408.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 408.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 406 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 406 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 406 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 403.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 403.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 403.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 400.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 400.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 400.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 397.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 397.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 397.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 394.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 394.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 394.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 392 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 392 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 392 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 389.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 389.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 389.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 386.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 386.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 386.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 383.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 383.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 383.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 380.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 380.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 380.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 378 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 378 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 378 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 375.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 375.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 375.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 372.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 372.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 372.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 369.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 369.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 369.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 366.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 366.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 366.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 364 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 364 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 364 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 361.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 361.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 361.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 358.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 358.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 358.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 355.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 355.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 355.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 352.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 352.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 352.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 350 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 350 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 350 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 347.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 347.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 347.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 344.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 344.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 344.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 341.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 341.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 341.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 143.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 143.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 143.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 408.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 408.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 408.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 406 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 406 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 406 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 403.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 403.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 403.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 400.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 400.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 400.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 397.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 397.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 397.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 394.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 394.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 394.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 392 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 392 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 392 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 389.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 389.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 389.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 386.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 386.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 386.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 383.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 383.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 383.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 380.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 380.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 380.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 378 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 378 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 378 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 375.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 375.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 375.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 372.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 372.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 372.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 369.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 369.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 369.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 366.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 366.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 366.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 364 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 364 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 364 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 361.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 361.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 361.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 358.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 358.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 358.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 355.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 355.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 355.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 352.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 352.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 352.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 350 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 350 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 350 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 347.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 347.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 347.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 344.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 344.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 344.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 341.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 341.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 341.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 87.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 87.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 87.14 2.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 408.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 408.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 408.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 406 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 406 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 406 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 403.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 403.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 403.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 400.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 400.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 400.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 397.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 397.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 397.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 394.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 394.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 394.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 392 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 392 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 392 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 389.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 389.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 389.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 386.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 386.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 386.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 383.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 383.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 383.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 380.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 380.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 380.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 378 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 378 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 378 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 375.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 375.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 375.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 372.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 372.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 372.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 369.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 369.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 369.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 366.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 366.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 366.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 364 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 364 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 364 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 361.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 361.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 361.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 358.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 358.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 358.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 355.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 355.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 355.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 352.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 352.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 352.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 350 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 350 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 350 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 347.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 347.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 347.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 344.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 344.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 344.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 341.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 341.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 341.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 338.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 338.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 338.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 336 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 336 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 336 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 333.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 333.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 333.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 330.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 330.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 330.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 327.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 327.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 327.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 324.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 324.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 324.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 322 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 322 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 322 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 319.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 319.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 319.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 316.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 316.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 316.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 313.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 313.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 313.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 310.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 310.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 310.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 308 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 308 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 308 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 305.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 305.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 305.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 302.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 302.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 302.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 299.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 299.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 299.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 296.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 296.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 296.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 294 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 294 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 294 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 291.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 291.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 291.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 288.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 288.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 288.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 285.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 285.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 285.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 282.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 282.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 282.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 280 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 280 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 280 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 277.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 277.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 277.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 274.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 274.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 274.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 271.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 271.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 271.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 268.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 268.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 268.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 266 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 266 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 266 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 263.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 263.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 263.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 260.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 260.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 260.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 257.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 257.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 257.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 254.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 254.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 254.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 252 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 252 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 252 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 249.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 249.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 249.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 246.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 246.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 246.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 243.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 243.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 243.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 240.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 240.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 240.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 238 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 238 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 238 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 235.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 235.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 235.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 232.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 232.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 232.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 229.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 229.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 229.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 226.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 226.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 226.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 224 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 224 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 224 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 221.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 221.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 221.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 218.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 218.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 218.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 215.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 215.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 215.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 212.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 212.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 212.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 210 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 210 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 210 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 207.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 207.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 207.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 204.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 204.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 204.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 201.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 201.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 201.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 198.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 198.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 198.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 196 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 196 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 196 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 193.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 193.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 193.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 190.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 190.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 190.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 187.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 187.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 187.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 184.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 184.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 184.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 182 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 182 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 182 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 179.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 179.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 179.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 176.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 176.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 176.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 173.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 173.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 173.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 170.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 170.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 170.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 168 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 168 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 168 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 165.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 165.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 165.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 162.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 162.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 162.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 159.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 159.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 159.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 156.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 156.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 156.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 154 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 154 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 154 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 151.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 151.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 151.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 148.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 148.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 148.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 145.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 145.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 145.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 142.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 142.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 142.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 140 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 140 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 140 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 137.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 137.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 137.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 134.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 134.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 134.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 131.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 131.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 131.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 128.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 128.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 128.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 126 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 126 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 126 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 123.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 123.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 123.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 120.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 120.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 120.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 117.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 117.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 117.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 114.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 114.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 114.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 112 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 112 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 112 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 109.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 109.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 109.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 106.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 106.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 106.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 103.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 103.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 103.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 100.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 100.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 100.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 98 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 98 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 98 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 95.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 95.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 95.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 92.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 92.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 92.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 89.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 89.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 89.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 86.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 86.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 86.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 84 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 84 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 84 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 81.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 81.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 81.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 78.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 78.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 78.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 75.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 75.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 75.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 72.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 72.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 72.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 70 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 70 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 70 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 67.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 67.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 67.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 64.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 64.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 64.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 61.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 61.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 61.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 58.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 58.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 58.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 56 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 56 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 56 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 53.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 53.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 53.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 50.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 50.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 50.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 47.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 47.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 47.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 44.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 44.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 44.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 42 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 42 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 42 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 39.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 39.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 39.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 36.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 36.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 36.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 33.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 33.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 33.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 30.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 30.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 30.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 28 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 28 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 28 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 25.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 25.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 25.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 22.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 22.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 22.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 19.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 19.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 19.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 16.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 16.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 16.8 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 14 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 14 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 14 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 11.2 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 11.2 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 11.2 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 8.4 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 8.4 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 8.4 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 5.6 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 5.6 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 5.6 via1_2_400_200_1_1_300_300 ;
      VIA 31.14 2.8 via3_4_400_200_1_1_320_320 ;
      VIA 31.14 2.8 via2_3_400_200_1_1_320_320 ;
      VIA 31.14 2.8 via1_2_400_200_1_1_300_300 ;
    END
  END VDD
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 260.4 0.14 260.54 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 97.44 293.635 97.58 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 253.68 293.635 253.82 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  78.425 0 78.565 0.14 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 201.6 293.635 201.74 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  215.065 410.15 215.205 410.29 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  286.185 0 286.325 0.14 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 104.16 0.14 104.3 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 156.24 0.14 156.38 ;
    END
  END addr[8]
  PIN ce
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 338.24 0.14 338.38 ;
    END
  END ce
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 123.76 293.635 123.9 ;
    END
  END clk
  PIN di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  162.985 410.15 163.125 410.29 ;
    END
  END di[0]
  PIN di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 208.32 0.14 208.46 ;
    END
  END di[10]
  PIN di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  208.345 0 208.485 0.14 ;
    END
  END di[11]
  PIN di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 149.52 293.635 149.66 ;
    END
  END di[12]
  PIN di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 305.76 293.635 305.9 ;
    END
  END di[13]
  PIN di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 364.56 0.14 364.7 ;
    END
  END di[14]
  PIN di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 234.08 0.14 234.22 ;
    END
  END di[15]
  PIN di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 383.6 293.635 383.74 ;
    END
  END di[16]
  PIN di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  260.425 0 260.565 0.14 ;
    END
  END di[17]
  PIN di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 19.6 293.635 19.74 ;
    END
  END di[18]
  PIN di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 286.16 0.14 286.3 ;
    END
  END di[19]
  PIN di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 71.68 293.635 71.82 ;
    END
  END di[1]
  PIN di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  85.145 410.15 85.285 410.29 ;
    END
  END di[20]
  PIN di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  241.385 410.15 241.525 410.29 ;
    END
  END di[2]
  PIN di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 52.08 0.14 52.22 ;
    END
  END di[3]
  PIN di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  137.225 410.15 137.365 410.29 ;
    END
  END di[4]
  PIN di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 78.4 0.14 78.54 ;
    END
  END di[5]
  PIN di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  292.905 410.15 293.045 410.29 ;
    END
  END di[6]
  PIN di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 331.52 293.635 331.66 ;
    END
  END di[7]
  PIN di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 390.32 0.14 390.46 ;
    END
  END di[8]
  PIN di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  189.305 410.15 189.445 410.29 ;
    END
  END di[9]
  PIN doq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  26.345 0 26.485 0.14 ;
    END
  END doq[0]
  PIN doq[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  0.585 0 0.725 0.14 ;
    END
  END doq[10]
  PIN doq[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  33.065 410.15 33.205 410.29 ;
    END
  END doq[11]
  PIN doq[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 357.84 293.635 357.98 ;
    END
  END doq[12]
  PIN doq[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  130.505 0 130.645 0.14 ;
    END
  END doq[13]
  PIN doq[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 279.44 293.635 279.58 ;
    END
  END doq[14]
  PIN doq[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 45.36 293.635 45.5 ;
    END
  END doq[15]
  PIN doq[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  110.905 410.15 111.045 410.29 ;
    END
  END doq[16]
  PIN doq[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 175.84 293.635 175.98 ;
    END
  END doq[17]
  PIN doq[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  52.105 0 52.245 0.14 ;
    END
  END doq[18]
  PIN doq[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  104.185 0 104.325 0.14 ;
    END
  END doq[19]
  PIN doq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  156.265 0 156.405 0.14 ;
    END
  END doq[1]
  PIN doq[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 26.32 0.14 26.46 ;
    END
  END doq[20]
  PIN doq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  182.585 0 182.725 0.14 ;
    END
  END doq[2]
  PIN doq[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 182.56 0.14 182.7 ;
    END
  END doq[3]
  PIN doq[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  267.145 410.15 267.285 410.29 ;
    END
  END doq[4]
  PIN doq[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  7.305 410.15 7.445 410.29 ;
    END
  END doq[5]
  PIN doq[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  58.825 410.15 58.965 410.29 ;
    END
  END doq[6]
  PIN doq[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT  234.665 0 234.805 0.14 ;
    END
  END doq[7]
  PIN doq[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 130.48 0.14 130.62 ;
    END
  END doq[8]
  PIN doq[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  0 312.48 0.14 312.62 ;
    END
  END doq[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT  293.495 227.36 293.635 227.5 ;
    END
  END we
  OBS
    LAYER metal1 ;
     RECT  0 0 293.635 410.29 ;
    LAYER metal2 ;
     RECT  0 0 293.635 410.29 ;
    LAYER metal3 ;
     RECT  0 0 293.635 410.29 ;
    LAYER metal4 ;
     RECT  0 0 293.635 410.29 ;
    LAYER metal5 ;
     RECT  0 0 293.635 410.29 ;
    LAYER metal6 ;
     RECT  0 0 293.635 410.29 ;
    LAYER metal7 ;
     RECT  0 0 293.635 410.29 ;
    LAYER metal8 ;
     RECT  0 0 293.635 410.29 ;
    LAYER metal9 ;
     RECT  0 0 293.635 410.29 ;
  END
END or1200_spram4
END LIBRARY
