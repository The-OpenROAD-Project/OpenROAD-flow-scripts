VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_64x7
  FOREIGN fakeram130_64x7 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 104.500 BY 900.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 27.550 0.900 28.450 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 55.550 0.900 56.450 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 83.550 0.900 84.450 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 111.550 0.900 112.450 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.550 0.900 140.450 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 167.550 0.900 168.450 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 195.550 0.900 196.450 ;
    END
  END w_mask_in[6]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 195.550 0.900 196.450 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 223.550 0.900 224.450 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 251.550 0.900 252.450 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 279.550 0.900 280.450 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 307.550 0.900 308.450 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 335.550 0.900 336.450 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 363.550 0.900 364.450 ;
    END
  END rd_out[6]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 363.550 0.900 364.450 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 391.550 0.900 392.450 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 419.550 0.900 420.450 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 447.550 0.900 448.450 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 475.550 0.900 476.450 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 503.550 0.900 504.450 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 531.550 0.900 532.450 ;
    END
  END wd_in[6]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 531.550 0.900 532.450 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 559.550 0.900 560.450 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 587.550 0.900 588.450 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 615.550 0.900 616.450 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 643.550 0.900 644.450 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 671.550 0.900 672.450 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 671.550 0.900 672.450 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 699.550 0.900 700.450 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 727.550 0.900 728.450 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 26.200 28.000 29.800 872.000 ;
      RECT 71.000 28.000 74.600 872.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 48.600 28.000 52.200 872.000 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 104.500 900.000 ;
    LAYER met2 ;
    RECT 0 0 104.500 900.000 ;
    LAYER met3 ;
    RECT 0.900 0 104.500 900.000 ;
    RECT 0 0.000 0.900 27.550 ;
    RECT 0 28.450 0.900 55.550 ;
    RECT 0 56.450 0.900 83.550 ;
    RECT 0 84.450 0.900 111.550 ;
    RECT 0 112.450 0.900 139.550 ;
    RECT 0 140.450 0.900 167.550 ;
    RECT 0 168.450 0.900 195.550 ;
    RECT 0 196.450 0.900 195.550 ;
    RECT 0 196.450 0.900 223.550 ;
    RECT 0 224.450 0.900 251.550 ;
    RECT 0 252.450 0.900 279.550 ;
    RECT 0 280.450 0.900 307.550 ;
    RECT 0 308.450 0.900 335.550 ;
    RECT 0 336.450 0.900 363.550 ;
    RECT 0 364.450 0.900 363.550 ;
    RECT 0 364.450 0.900 391.550 ;
    RECT 0 392.450 0.900 419.550 ;
    RECT 0 420.450 0.900 447.550 ;
    RECT 0 448.450 0.900 475.550 ;
    RECT 0 476.450 0.900 503.550 ;
    RECT 0 504.450 0.900 531.550 ;
    RECT 0 532.450 0.900 531.550 ;
    RECT 0 532.450 0.900 559.550 ;
    RECT 0 560.450 0.900 587.550 ;
    RECT 0 588.450 0.900 615.550 ;
    RECT 0 616.450 0.900 643.550 ;
    RECT 0 644.450 0.900 671.550 ;
    RECT 0 672.450 0.900 671.550 ;
    RECT 0 672.450 0.900 699.550 ;
    RECT 0 700.450 0.900 727.550 ;
    RECT 0 728.450 0.900 900.000 ;
    LAYER met4 ;
    RECT 0 0 104.500 28.000 ;
    RECT 0 872.000 104.500 900.000 ;
    RECT 0.000 28.000 26.200 872.000 ;
    RECT 29.800 28.000 48.600 872.000 ;
    RECT 52.200 28.000 71.000 872.000 ;
    RECT 74.600 28.000 104.500 872.000 ;
    LAYER OVERLAP ;
    RECT 0 0 104.500 900.000 ;
  END
END fakeram130_64x7

END LIBRARY
