module RegisterSRAM(
  input         clock,
  input  [6:0]  io_read_0_address,
                io_read_1_address,
                io_read_2_address,
                io_read_3_address,
                io_read_4_address,
                io_read_5_address,
                io_read_6_address,
                io_read_7_address,
  input         io_write_0_write,
  input  [6:0]  io_write_0_address,
  input  [63:0] io_write_0_value,
  input         io_write_0_byteMask_0,
                io_write_0_byteMask_1,
                io_write_0_byteMask_2,
                io_write_0_byteMask_3,
                io_write_0_byteMask_4,
                io_write_0_byteMask_5,
                io_write_0_byteMask_6,
                io_write_0_byteMask_7,
                io_write_1_write,
  input  [6:0]  io_write_1_address,
  input  [63:0] io_write_1_value,
  input         io_write_1_byteMask_0,
                io_write_1_byteMask_1,
                io_write_1_byteMask_2,
                io_write_1_byteMask_3,
                io_write_1_byteMask_4,
                io_write_1_byteMask_5,
                io_write_1_byteMask_6,
                io_write_1_byteMask_7,
                io_write_2_write,
  input  [6:0]  io_write_2_address,
  input  [63:0] io_write_2_value,
  input         io_write_2_byteMask_0,
                io_write_2_byteMask_1,
                io_write_2_byteMask_2,
                io_write_2_byteMask_3,
                io_write_2_byteMask_4,
                io_write_2_byteMask_5,
                io_write_2_byteMask_6,
                io_write_2_byteMask_7,
                io_write_3_write,
  input  [6:0]  io_write_3_address,
  input  [63:0] io_write_3_value,
  input         io_write_3_byteMask_0,
                io_write_3_byteMask_1,
                io_write_3_byteMask_2,
                io_write_3_byteMask_3,
                io_write_3_byteMask_4,
                io_write_3_byteMask_5,
                io_write_3_byteMask_6,
                io_write_3_byteMask_7,
  output [63:0] io_read_0_value,
                io_read_1_value,
                io_read_2_value,
                io_read_3_value,
                io_read_4_value,
                io_read_5_value,
                io_read_6_value,
                io_read_7_value
);

  ram_32x64 ram_ext (
    .R0_addr (io_read_7_address[4:0]),
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R1_addr (io_read_6_address[4:0]),
    .R1_en   (1'h1),
    .R1_clk  (clock),
    .R2_addr (io_read_5_address[4:0]),
    .R2_en   (1'h1),
    .R2_clk  (clock),
    .R3_addr (io_read_4_address[4:0]),
    .R3_en   (1'h1),
    .R3_clk  (clock),
    .R4_addr (io_read_3_address[4:0]),
    .R4_en   (1'h1),
    .R4_clk  (clock),
    .R5_addr (io_read_2_address[4:0]),
    .R5_en   (1'h1),
    .R5_clk  (clock),
    .R6_addr (io_read_1_address[4:0]),
    .R6_en   (1'h1),
    .R6_clk  (clock),
    .R7_addr (io_read_0_address[4:0]),
    .R7_en   (1'h1),
    .R7_clk  (clock),
    .W0_addr (io_write_3_address[4:0]),
    .W0_en   (io_write_3_write),
    .W0_clk  (clock),
    .W0_data (io_write_3_value),
    .W0_mask
      ({io_write_3_byteMask_7,
        io_write_3_byteMask_6,
        io_write_3_byteMask_5,
        io_write_3_byteMask_4,
        io_write_3_byteMask_3,
        io_write_3_byteMask_2,
        io_write_3_byteMask_1,
        io_write_3_byteMask_0}),
    .W1_addr (io_write_2_address[4:0]),
    .W1_en   (io_write_2_write),
    .W1_clk  (clock),
    .W1_data (io_write_2_value),
    .W1_mask
      ({io_write_2_byteMask_7,
        io_write_2_byteMask_6,
        io_write_2_byteMask_5,
        io_write_2_byteMask_4,
        io_write_2_byteMask_3,
        io_write_2_byteMask_2,
        io_write_2_byteMask_1,
        io_write_2_byteMask_0}),
    .W2_addr (io_write_1_address[4:0]),
    .W2_en   (io_write_1_write),
    .W2_clk  (clock),
    .W2_data (io_write_1_value),
    .W2_mask
      ({io_write_1_byteMask_7,
        io_write_1_byteMask_6,
        io_write_1_byteMask_5,
        io_write_1_byteMask_4,
        io_write_1_byteMask_3,
        io_write_1_byteMask_2,
        io_write_1_byteMask_1,
        io_write_1_byteMask_0}),
    .W3_addr (io_write_0_address[4:0]),
    .W3_en   (io_write_0_write),
    .W3_clk  (clock),
    .W3_data (io_write_0_value),
    .W3_mask
      ({io_write_0_byteMask_7,
        io_write_0_byteMask_6,
        io_write_0_byteMask_5,
        io_write_0_byteMask_4,
        io_write_0_byteMask_3,
        io_write_0_byteMask_2,
        io_write_0_byteMask_1,
        io_write_0_byteMask_0}),
    .R0_data (io_read_7_value),
    .R1_data (io_read_6_value),
    .R2_data (io_read_5_value),
    .R3_data (io_read_4_value),
    .R4_data (io_read_3_value),
    .R5_data (io_read_2_value),
    .R6_data (io_read_1_value),
    .R7_data (io_read_0_value)
  );
endmodule

