VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_64x7
  FOREIGN fakeram45_64x7 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 10.640 BY 36.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.065 0.070 2.135 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.115 0.070 3.185 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.215 0.070 5.285 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.265 0.070 6.335 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.315 0.070 7.385 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[6]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.415 0.070 9.485 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.465 0.070 10.535 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.515 0.070 11.585 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.615 0.070 13.685 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END rd_out[6]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.665 0.070 14.735 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.715 0.070 15.785 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.815 0.070 17.885 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.865 0.070 18.935 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.915 0.070 19.985 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END wd_in[6]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.015 0.070 22.085 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.065 0.070 23.135 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.115 0.070 24.185 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.215 0.070 26.285 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.215 0.070 26.285 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.265 0.070 27.335 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.315 0.070 28.385 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.960 2.100 2.240 34.300 ;
      RECT 5.320 2.100 5.600 34.300 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 3.640 2.100 3.920 34.300 ;
      RECT 7.000 2.100 7.280 34.300 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 10.640 36.400 ;
    LAYER metal2 ;
    RECT 0 0 10.640 36.400 ;
    LAYER metal3 ;
    RECT 0.070 0 10.640 36.400 ;
    RECT 0 0.000 0.070 2.065 ;
    RECT 0 2.135 0.070 3.115 ;
    RECT 0 3.185 0.070 4.165 ;
    RECT 0 4.235 0.070 5.215 ;
    RECT 0 5.285 0.070 6.265 ;
    RECT 0 6.335 0.070 7.315 ;
    RECT 0 7.385 0.070 8.365 ;
    RECT 0 8.435 0.070 8.365 ;
    RECT 0 8.435 0.070 9.415 ;
    RECT 0 9.485 0.070 10.465 ;
    RECT 0 10.535 0.070 11.515 ;
    RECT 0 11.585 0.070 12.565 ;
    RECT 0 12.635 0.070 13.615 ;
    RECT 0 13.685 0.070 14.665 ;
    RECT 0 14.735 0.070 14.665 ;
    RECT 0 14.735 0.070 15.715 ;
    RECT 0 15.785 0.070 16.765 ;
    RECT 0 16.835 0.070 17.815 ;
    RECT 0 17.885 0.070 18.865 ;
    RECT 0 18.935 0.070 19.915 ;
    RECT 0 19.985 0.070 20.965 ;
    RECT 0 21.035 0.070 20.965 ;
    RECT 0 21.035 0.070 22.015 ;
    RECT 0 22.085 0.070 23.065 ;
    RECT 0 23.135 0.070 24.115 ;
    RECT 0 24.185 0.070 25.165 ;
    RECT 0 25.235 0.070 26.215 ;
    RECT 0 26.285 0.070 26.215 ;
    RECT 0 26.285 0.070 27.265 ;
    RECT 0 27.335 0.070 28.315 ;
    RECT 0 28.385 0.070 36.400 ;
    LAYER metal4 ;
    RECT 0 0 10.640 2.100 ;
    RECT 0 34.300 10.640 36.400 ;
    RECT 0.000 2.100 1.960 34.300 ;
    RECT 2.240 2.100 3.640 34.300 ;
    RECT 3.920 2.100 5.320 34.300 ;
    RECT 5.600 2.100 7.000 34.300 ;
    RECT 7.280 2.100 10.640 34.300 ;
    LAYER OVERLAP ;
    RECT 0 0 10.640 36.400 ;
  END
END fakeram45_64x7

END LIBRARY
