module MuxTest_width_16_inputs_16_outputs_8_pipeline_0( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [3:0]  io_selects_0_0, // @[:@6.4]
  input  [3:0]  io_selects_0_1, // @[:@6.4]
  input  [3:0]  io_selects_1_0, // @[:@6.4]
  input  [3:0]  io_selects_1_1, // @[:@6.4]
  input  [3:0]  io_selects_2_0, // @[:@6.4]
  input  [3:0]  io_selects_2_1, // @[:@6.4]
  input  [3:0]  io_selects_3_0, // @[:@6.4]
  input  [3:0]  io_selects_3_1, // @[:@6.4]
  input  [3:0]  io_selects_4_0, // @[:@6.4]
  input  [3:0]  io_selects_4_1, // @[:@6.4]
  input  [3:0]  io_selects_5_0, // @[:@6.4]
  input  [3:0]  io_selects_5_1, // @[:@6.4]
  input  [3:0]  io_selects_6_0, // @[:@6.4]
  input  [3:0]  io_selects_6_1, // @[:@6.4]
  input  [3:0]  io_selects_7_0, // @[:@6.4]
  input  [3:0]  io_selects_7_1, // @[:@6.4]
  input  [2:0]  io_operation_0, // @[:@6.4]
  input  [2:0]  io_operation_1, // @[:@6.4]
  input  [2:0]  io_operation_2, // @[:@6.4]
  input  [2:0]  io_operation_3, // @[:@6.4]
  input  [2:0]  io_operation_4, // @[:@6.4]
  input  [2:0]  io_operation_5, // @[:@6.4]
  input  [2:0]  io_operation_6, // @[:@6.4]
  input  [2:0]  io_operation_7, // @[:@6.4]
  input  [15:0] io_inputs_0, // @[:@6.4]
  input  [15:0] io_inputs_1, // @[:@6.4]
  input  [15:0] io_inputs_2, // @[:@6.4]
  input  [15:0] io_inputs_3, // @[:@6.4]
  input  [15:0] io_inputs_4, // @[:@6.4]
  input  [15:0] io_inputs_5, // @[:@6.4]
  input  [15:0] io_inputs_6, // @[:@6.4]
  input  [15:0] io_inputs_7, // @[:@6.4]
  input  [15:0] io_inputs_8, // @[:@6.4]
  input  [15:0] io_inputs_9, // @[:@6.4]
  input  [15:0] io_inputs_10, // @[:@6.4]
  input  [15:0] io_inputs_11, // @[:@6.4]
  input  [15:0] io_inputs_12, // @[:@6.4]
  input  [15:0] io_inputs_13, // @[:@6.4]
  input  [15:0] io_inputs_14, // @[:@6.4]
  input  [15:0] io_inputs_15, // @[:@6.4]
  output [15:0] io_outputs_0, // @[:@6.4]
  output [15:0] io_outputs_1, // @[:@6.4]
  output [15:0] io_outputs_2, // @[:@6.4]
  output [15:0] io_outputs_3, // @[:@6.4]
  output [15:0] io_outputs_4, // @[:@6.4]
  output [15:0] io_outputs_5, // @[:@6.4]
  output [15:0] io_outputs_6, // @[:@6.4]
  output [15:0] io_outputs_7 // @[:@6.4]
);
  wire [15:0] _GEN_1; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_2; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_3; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_4; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_5; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_6; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_7; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_8; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_9; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_10; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_11; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_12; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_13; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_14; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_15; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_17; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_18; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_19; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_20; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_21; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_22; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_23; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_24; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_25; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_26; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_27; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_28; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_29; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_30; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _GEN_31; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [16:0] _T_418; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [15:0] _T_419; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@9.4]
  wire [31:0] _T_421; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@10.4]
  wire [15:0] _T_423; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@11.4]
  wire  _T_424; // @[Mux.scala 46:19:@12.4]
  wire [15:0] _T_425; // @[Mux.scala 46:16:@13.4]
  wire  _T_426; // @[Mux.scala 46:19:@14.4]
  wire [31:0] _T_427; // @[Mux.scala 46:16:@15.4]
  wire  _T_428; // @[Mux.scala 46:19:@16.4]
  wire [31:0] _T_429; // @[Mux.scala 46:16:@17.4]
  wire  _T_430; // @[Mux.scala 46:19:@18.4]
  wire [31:0] _T_431; // @[Mux.scala 46:16:@19.4]
  wire [15:0] _GEN_33; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_34; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_35; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_36; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_37; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_38; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_39; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_40; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_41; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_42; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_43; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_44; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_45; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_46; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_47; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_49; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_50; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_51; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_52; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_53; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_54; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_55; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_56; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_57; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_58; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_59; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_60; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_61; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_62; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _GEN_63; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [16:0] _T_435; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  wire [15:0] _T_436; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@21.4]
  wire [31:0] _T_438; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@22.4]
  wire [15:0] _T_440; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@23.4]
  wire  _T_441; // @[Mux.scala 46:19:@24.4]
  wire [15:0] _T_442; // @[Mux.scala 46:16:@25.4]
  wire  _T_443; // @[Mux.scala 46:19:@26.4]
  wire [31:0] _T_444; // @[Mux.scala 46:16:@27.4]
  wire  _T_445; // @[Mux.scala 46:19:@28.4]
  wire [31:0] _T_446; // @[Mux.scala 46:16:@29.4]
  wire  _T_447; // @[Mux.scala 46:19:@30.4]
  wire [31:0] _T_448; // @[Mux.scala 46:16:@31.4]
  wire [15:0] _GEN_65; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_66; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_67; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_68; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_69; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_70; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_71; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_72; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_73; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_74; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_75; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_76; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_77; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_78; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_79; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_81; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_82; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_83; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_84; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_85; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_86; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_87; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_88; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_89; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_90; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_91; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_92; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_93; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_94; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _GEN_95; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [16:0] _T_452; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  wire [15:0] _T_453; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@33.4]
  wire [31:0] _T_455; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@34.4]
  wire [15:0] _T_457; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@35.4]
  wire  _T_458; // @[Mux.scala 46:19:@36.4]
  wire [15:0] _T_459; // @[Mux.scala 46:16:@37.4]
  wire  _T_460; // @[Mux.scala 46:19:@38.4]
  wire [31:0] _T_461; // @[Mux.scala 46:16:@39.4]
  wire  _T_462; // @[Mux.scala 46:19:@40.4]
  wire [31:0] _T_463; // @[Mux.scala 46:16:@41.4]
  wire  _T_464; // @[Mux.scala 46:19:@42.4]
  wire [31:0] _T_465; // @[Mux.scala 46:16:@43.4]
  wire [15:0] _GEN_97; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_98; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_99; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_100; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_101; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_102; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_103; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_104; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_105; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_106; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_107; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_108; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_109; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_110; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_111; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_113; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_114; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_115; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_116; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_117; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_118; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_119; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_120; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_121; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_122; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_123; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_124; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_125; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_126; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _GEN_127; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [16:0] _T_469; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  wire [15:0] _T_470; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@45.4]
  wire [31:0] _T_472; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@46.4]
  wire [15:0] _T_474; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@47.4]
  wire  _T_475; // @[Mux.scala 46:19:@48.4]
  wire [15:0] _T_476; // @[Mux.scala 46:16:@49.4]
  wire  _T_477; // @[Mux.scala 46:19:@50.4]
  wire [31:0] _T_478; // @[Mux.scala 46:16:@51.4]
  wire  _T_479; // @[Mux.scala 46:19:@52.4]
  wire [31:0] _T_480; // @[Mux.scala 46:16:@53.4]
  wire  _T_481; // @[Mux.scala 46:19:@54.4]
  wire [31:0] _T_482; // @[Mux.scala 46:16:@55.4]
  wire [15:0] _GEN_129; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_130; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_131; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_132; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_133; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_134; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_135; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_136; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_137; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_138; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_139; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_140; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_141; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_142; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_143; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_145; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_146; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_147; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_148; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_149; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_150; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_151; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_152; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_153; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_154; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_155; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_156; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_157; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_158; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _GEN_159; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [16:0] _T_486; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  wire [15:0] _T_487; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@57.4]
  wire [31:0] _T_489; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@58.4]
  wire [15:0] _T_491; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@59.4]
  wire  _T_492; // @[Mux.scala 46:19:@60.4]
  wire [15:0] _T_493; // @[Mux.scala 46:16:@61.4]
  wire  _T_494; // @[Mux.scala 46:19:@62.4]
  wire [31:0] _T_495; // @[Mux.scala 46:16:@63.4]
  wire  _T_496; // @[Mux.scala 46:19:@64.4]
  wire [31:0] _T_497; // @[Mux.scala 46:16:@65.4]
  wire  _T_498; // @[Mux.scala 46:19:@66.4]
  wire [31:0] _T_499; // @[Mux.scala 46:16:@67.4]
  wire [15:0] _GEN_161; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_162; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_163; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_164; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_165; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_166; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_167; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_168; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_169; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_170; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_171; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_172; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_173; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_174; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_175; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_177; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_178; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_179; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_180; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_181; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_182; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_183; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_184; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_185; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_186; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_187; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_188; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_189; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_190; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _GEN_191; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [16:0] _T_503; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  wire [15:0] _T_504; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@69.4]
  wire [31:0] _T_506; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@70.4]
  wire [15:0] _T_508; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@71.4]
  wire  _T_509; // @[Mux.scala 46:19:@72.4]
  wire [15:0] _T_510; // @[Mux.scala 46:16:@73.4]
  wire  _T_511; // @[Mux.scala 46:19:@74.4]
  wire [31:0] _T_512; // @[Mux.scala 46:16:@75.4]
  wire  _T_513; // @[Mux.scala 46:19:@76.4]
  wire [31:0] _T_514; // @[Mux.scala 46:16:@77.4]
  wire  _T_515; // @[Mux.scala 46:19:@78.4]
  wire [31:0] _T_516; // @[Mux.scala 46:16:@79.4]
  wire [15:0] _GEN_193; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_194; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_195; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_196; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_197; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_198; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_199; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_200; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_201; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_202; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_203; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_204; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_205; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_206; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_207; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_209; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_210; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_211; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_212; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_213; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_214; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_215; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_216; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_217; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_218; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_219; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_220; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_221; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_222; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _GEN_223; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [16:0] _T_520; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  wire [15:0] _T_521; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@81.4]
  wire [31:0] _T_523; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@82.4]
  wire [15:0] _T_525; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@83.4]
  wire  _T_526; // @[Mux.scala 46:19:@84.4]
  wire [15:0] _T_527; // @[Mux.scala 46:16:@85.4]
  wire  _T_528; // @[Mux.scala 46:19:@86.4]
  wire [31:0] _T_529; // @[Mux.scala 46:16:@87.4]
  wire  _T_530; // @[Mux.scala 46:19:@88.4]
  wire [31:0] _T_531; // @[Mux.scala 46:16:@89.4]
  wire  _T_532; // @[Mux.scala 46:19:@90.4]
  wire [31:0] _T_533; // @[Mux.scala 46:16:@91.4]
  wire [15:0] _GEN_225; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_226; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_227; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_228; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_229; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_230; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_231; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_232; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_233; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_234; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_235; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_236; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_237; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_238; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_239; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_241; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_242; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_243; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_244; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_245; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_246; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_247; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_248; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_249; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_250; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_251; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_252; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_253; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_254; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _GEN_255; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [16:0] _T_537; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  wire [15:0] _T_538; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@93.4]
  wire [31:0] _T_540; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@94.4]
  wire [15:0] _T_542; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@95.4]
  wire  _T_543; // @[Mux.scala 46:19:@96.4]
  wire [15:0] _T_544; // @[Mux.scala 46:16:@97.4]
  wire  _T_545; // @[Mux.scala 46:19:@98.4]
  wire [31:0] _T_546; // @[Mux.scala 46:16:@99.4]
  wire  _T_547; // @[Mux.scala 46:19:@100.4]
  wire [31:0] _T_548; // @[Mux.scala 46:16:@101.4]
  wire  _T_549; // @[Mux.scala 46:19:@102.4]
  wire [31:0] _T_550; // @[Mux.scala 46:16:@103.4]
  assign _GEN_1 = 4'h1 == io_selects_0_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_2 = 4'h2 == io_selects_0_0 ? io_inputs_2 : _GEN_1; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_3 = 4'h3 == io_selects_0_0 ? io_inputs_3 : _GEN_2; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_4 = 4'h4 == io_selects_0_0 ? io_inputs_4 : _GEN_3; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_5 = 4'h5 == io_selects_0_0 ? io_inputs_5 : _GEN_4; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_6 = 4'h6 == io_selects_0_0 ? io_inputs_6 : _GEN_5; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_7 = 4'h7 == io_selects_0_0 ? io_inputs_7 : _GEN_6; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_8 = 4'h8 == io_selects_0_0 ? io_inputs_8 : _GEN_7; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_9 = 4'h9 == io_selects_0_0 ? io_inputs_9 : _GEN_8; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_10 = 4'ha == io_selects_0_0 ? io_inputs_10 : _GEN_9; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_11 = 4'hb == io_selects_0_0 ? io_inputs_11 : _GEN_10; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_12 = 4'hc == io_selects_0_0 ? io_inputs_12 : _GEN_11; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_13 = 4'hd == io_selects_0_0 ? io_inputs_13 : _GEN_12; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_14 = 4'he == io_selects_0_0 ? io_inputs_14 : _GEN_13; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_15 = 4'hf == io_selects_0_0 ? io_inputs_15 : _GEN_14; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_17 = 4'h1 == io_selects_0_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_18 = 4'h2 == io_selects_0_1 ? io_inputs_2 : _GEN_17; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_19 = 4'h3 == io_selects_0_1 ? io_inputs_3 : _GEN_18; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_20 = 4'h4 == io_selects_0_1 ? io_inputs_4 : _GEN_19; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_21 = 4'h5 == io_selects_0_1 ? io_inputs_5 : _GEN_20; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_22 = 4'h6 == io_selects_0_1 ? io_inputs_6 : _GEN_21; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_23 = 4'h7 == io_selects_0_1 ? io_inputs_7 : _GEN_22; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_24 = 4'h8 == io_selects_0_1 ? io_inputs_8 : _GEN_23; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_25 = 4'h9 == io_selects_0_1 ? io_inputs_9 : _GEN_24; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_26 = 4'ha == io_selects_0_1 ? io_inputs_10 : _GEN_25; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_27 = 4'hb == io_selects_0_1 ? io_inputs_11 : _GEN_26; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_28 = 4'hc == io_selects_0_1 ? io_inputs_12 : _GEN_27; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_29 = 4'hd == io_selects_0_1 ? io_inputs_13 : _GEN_28; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_30 = 4'he == io_selects_0_1 ? io_inputs_14 : _GEN_29; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_31 = 4'hf == io_selects_0_1 ? io_inputs_15 : _GEN_30; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _T_418 = _GEN_15 + _GEN_31; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _T_419 = _GEN_15 + _GEN_31; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@9.4]
  assign _T_421 = _GEN_15 * _GEN_31; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@10.4]
  assign _T_423 = _GEN_15 / _GEN_31; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@11.4]
  assign _T_424 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_425 = _T_424 ? _T_423 : 16'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_426 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_427 = _T_426 ? _T_421 : {{16'd0}, _T_425}; // @[Mux.scala 46:16:@15.4]
  assign _T_428 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_429 = _T_428 ? {{16'd0}, _T_419} : _T_427; // @[Mux.scala 46:16:@17.4]
  assign _T_430 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _T_431 = _T_430 ? {{16'd0}, _GEN_15} : _T_429; // @[Mux.scala 46:16:@19.4]
  assign _GEN_33 = 4'h1 == io_selects_1_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_34 = 4'h2 == io_selects_1_0 ? io_inputs_2 : _GEN_33; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_35 = 4'h3 == io_selects_1_0 ? io_inputs_3 : _GEN_34; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_36 = 4'h4 == io_selects_1_0 ? io_inputs_4 : _GEN_35; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_37 = 4'h5 == io_selects_1_0 ? io_inputs_5 : _GEN_36; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_38 = 4'h6 == io_selects_1_0 ? io_inputs_6 : _GEN_37; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_39 = 4'h7 == io_selects_1_0 ? io_inputs_7 : _GEN_38; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_40 = 4'h8 == io_selects_1_0 ? io_inputs_8 : _GEN_39; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_41 = 4'h9 == io_selects_1_0 ? io_inputs_9 : _GEN_40; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_42 = 4'ha == io_selects_1_0 ? io_inputs_10 : _GEN_41; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_43 = 4'hb == io_selects_1_0 ? io_inputs_11 : _GEN_42; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_44 = 4'hc == io_selects_1_0 ? io_inputs_12 : _GEN_43; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_45 = 4'hd == io_selects_1_0 ? io_inputs_13 : _GEN_44; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_46 = 4'he == io_selects_1_0 ? io_inputs_14 : _GEN_45; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_47 = 4'hf == io_selects_1_0 ? io_inputs_15 : _GEN_46; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_49 = 4'h1 == io_selects_1_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_50 = 4'h2 == io_selects_1_1 ? io_inputs_2 : _GEN_49; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_51 = 4'h3 == io_selects_1_1 ? io_inputs_3 : _GEN_50; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_52 = 4'h4 == io_selects_1_1 ? io_inputs_4 : _GEN_51; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_53 = 4'h5 == io_selects_1_1 ? io_inputs_5 : _GEN_52; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_54 = 4'h6 == io_selects_1_1 ? io_inputs_6 : _GEN_53; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_55 = 4'h7 == io_selects_1_1 ? io_inputs_7 : _GEN_54; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_56 = 4'h8 == io_selects_1_1 ? io_inputs_8 : _GEN_55; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_57 = 4'h9 == io_selects_1_1 ? io_inputs_9 : _GEN_56; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_58 = 4'ha == io_selects_1_1 ? io_inputs_10 : _GEN_57; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_59 = 4'hb == io_selects_1_1 ? io_inputs_11 : _GEN_58; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_60 = 4'hc == io_selects_1_1 ? io_inputs_12 : _GEN_59; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_61 = 4'hd == io_selects_1_1 ? io_inputs_13 : _GEN_60; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_62 = 4'he == io_selects_1_1 ? io_inputs_14 : _GEN_61; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_63 = 4'hf == io_selects_1_1 ? io_inputs_15 : _GEN_62; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _T_435 = _GEN_47 + _GEN_63; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@20.4]
  assign _T_436 = _GEN_47 + _GEN_63; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@21.4]
  assign _T_438 = _GEN_47 * _GEN_63; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@22.4]
  assign _T_440 = _GEN_47 / _GEN_63; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@23.4]
  assign _T_441 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_442 = _T_441 ? _T_440 : 16'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_443 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_444 = _T_443 ? _T_438 : {{16'd0}, _T_442}; // @[Mux.scala 46:16:@27.4]
  assign _T_445 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_446 = _T_445 ? {{16'd0}, _T_436} : _T_444; // @[Mux.scala 46:16:@29.4]
  assign _T_447 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _T_448 = _T_447 ? {{16'd0}, _GEN_47} : _T_446; // @[Mux.scala 46:16:@31.4]
  assign _GEN_65 = 4'h1 == io_selects_2_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_66 = 4'h2 == io_selects_2_0 ? io_inputs_2 : _GEN_65; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_67 = 4'h3 == io_selects_2_0 ? io_inputs_3 : _GEN_66; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_68 = 4'h4 == io_selects_2_0 ? io_inputs_4 : _GEN_67; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_69 = 4'h5 == io_selects_2_0 ? io_inputs_5 : _GEN_68; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_70 = 4'h6 == io_selects_2_0 ? io_inputs_6 : _GEN_69; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_71 = 4'h7 == io_selects_2_0 ? io_inputs_7 : _GEN_70; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_72 = 4'h8 == io_selects_2_0 ? io_inputs_8 : _GEN_71; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_73 = 4'h9 == io_selects_2_0 ? io_inputs_9 : _GEN_72; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_74 = 4'ha == io_selects_2_0 ? io_inputs_10 : _GEN_73; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_75 = 4'hb == io_selects_2_0 ? io_inputs_11 : _GEN_74; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_76 = 4'hc == io_selects_2_0 ? io_inputs_12 : _GEN_75; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_77 = 4'hd == io_selects_2_0 ? io_inputs_13 : _GEN_76; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_78 = 4'he == io_selects_2_0 ? io_inputs_14 : _GEN_77; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_79 = 4'hf == io_selects_2_0 ? io_inputs_15 : _GEN_78; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_81 = 4'h1 == io_selects_2_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_82 = 4'h2 == io_selects_2_1 ? io_inputs_2 : _GEN_81; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_83 = 4'h3 == io_selects_2_1 ? io_inputs_3 : _GEN_82; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_84 = 4'h4 == io_selects_2_1 ? io_inputs_4 : _GEN_83; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_85 = 4'h5 == io_selects_2_1 ? io_inputs_5 : _GEN_84; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_86 = 4'h6 == io_selects_2_1 ? io_inputs_6 : _GEN_85; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_87 = 4'h7 == io_selects_2_1 ? io_inputs_7 : _GEN_86; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_88 = 4'h8 == io_selects_2_1 ? io_inputs_8 : _GEN_87; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_89 = 4'h9 == io_selects_2_1 ? io_inputs_9 : _GEN_88; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_90 = 4'ha == io_selects_2_1 ? io_inputs_10 : _GEN_89; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_91 = 4'hb == io_selects_2_1 ? io_inputs_11 : _GEN_90; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_92 = 4'hc == io_selects_2_1 ? io_inputs_12 : _GEN_91; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_93 = 4'hd == io_selects_2_1 ? io_inputs_13 : _GEN_92; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_94 = 4'he == io_selects_2_1 ? io_inputs_14 : _GEN_93; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_95 = 4'hf == io_selects_2_1 ? io_inputs_15 : _GEN_94; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _T_452 = _GEN_79 + _GEN_95; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@32.4]
  assign _T_453 = _GEN_79 + _GEN_95; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@33.4]
  assign _T_455 = _GEN_79 * _GEN_95; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@34.4]
  assign _T_457 = _GEN_79 / _GEN_95; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@35.4]
  assign _T_458 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_459 = _T_458 ? _T_457 : 16'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_460 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_461 = _T_460 ? _T_455 : {{16'd0}, _T_459}; // @[Mux.scala 46:16:@39.4]
  assign _T_462 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_463 = _T_462 ? {{16'd0}, _T_453} : _T_461; // @[Mux.scala 46:16:@41.4]
  assign _T_464 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _T_465 = _T_464 ? {{16'd0}, _GEN_79} : _T_463; // @[Mux.scala 46:16:@43.4]
  assign _GEN_97 = 4'h1 == io_selects_3_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_98 = 4'h2 == io_selects_3_0 ? io_inputs_2 : _GEN_97; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_99 = 4'h3 == io_selects_3_0 ? io_inputs_3 : _GEN_98; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_100 = 4'h4 == io_selects_3_0 ? io_inputs_4 : _GEN_99; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_101 = 4'h5 == io_selects_3_0 ? io_inputs_5 : _GEN_100; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_102 = 4'h6 == io_selects_3_0 ? io_inputs_6 : _GEN_101; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_103 = 4'h7 == io_selects_3_0 ? io_inputs_7 : _GEN_102; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_104 = 4'h8 == io_selects_3_0 ? io_inputs_8 : _GEN_103; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_105 = 4'h9 == io_selects_3_0 ? io_inputs_9 : _GEN_104; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_106 = 4'ha == io_selects_3_0 ? io_inputs_10 : _GEN_105; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_107 = 4'hb == io_selects_3_0 ? io_inputs_11 : _GEN_106; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_108 = 4'hc == io_selects_3_0 ? io_inputs_12 : _GEN_107; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_109 = 4'hd == io_selects_3_0 ? io_inputs_13 : _GEN_108; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_110 = 4'he == io_selects_3_0 ? io_inputs_14 : _GEN_109; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_111 = 4'hf == io_selects_3_0 ? io_inputs_15 : _GEN_110; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_113 = 4'h1 == io_selects_3_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_114 = 4'h2 == io_selects_3_1 ? io_inputs_2 : _GEN_113; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_115 = 4'h3 == io_selects_3_1 ? io_inputs_3 : _GEN_114; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_116 = 4'h4 == io_selects_3_1 ? io_inputs_4 : _GEN_115; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_117 = 4'h5 == io_selects_3_1 ? io_inputs_5 : _GEN_116; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_118 = 4'h6 == io_selects_3_1 ? io_inputs_6 : _GEN_117; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_119 = 4'h7 == io_selects_3_1 ? io_inputs_7 : _GEN_118; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_120 = 4'h8 == io_selects_3_1 ? io_inputs_8 : _GEN_119; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_121 = 4'h9 == io_selects_3_1 ? io_inputs_9 : _GEN_120; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_122 = 4'ha == io_selects_3_1 ? io_inputs_10 : _GEN_121; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_123 = 4'hb == io_selects_3_1 ? io_inputs_11 : _GEN_122; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_124 = 4'hc == io_selects_3_1 ? io_inputs_12 : _GEN_123; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_125 = 4'hd == io_selects_3_1 ? io_inputs_13 : _GEN_124; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_126 = 4'he == io_selects_3_1 ? io_inputs_14 : _GEN_125; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_127 = 4'hf == io_selects_3_1 ? io_inputs_15 : _GEN_126; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _T_469 = _GEN_111 + _GEN_127; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@44.4]
  assign _T_470 = _GEN_111 + _GEN_127; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@45.4]
  assign _T_472 = _GEN_111 * _GEN_127; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@46.4]
  assign _T_474 = _GEN_111 / _GEN_127; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@47.4]
  assign _T_475 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_476 = _T_475 ? _T_474 : 16'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_477 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_478 = _T_477 ? _T_472 : {{16'd0}, _T_476}; // @[Mux.scala 46:16:@51.4]
  assign _T_479 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_480 = _T_479 ? {{16'd0}, _T_470} : _T_478; // @[Mux.scala 46:16:@53.4]
  assign _T_481 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _T_482 = _T_481 ? {{16'd0}, _GEN_111} : _T_480; // @[Mux.scala 46:16:@55.4]
  assign _GEN_129 = 4'h1 == io_selects_4_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_130 = 4'h2 == io_selects_4_0 ? io_inputs_2 : _GEN_129; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_131 = 4'h3 == io_selects_4_0 ? io_inputs_3 : _GEN_130; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_132 = 4'h4 == io_selects_4_0 ? io_inputs_4 : _GEN_131; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_133 = 4'h5 == io_selects_4_0 ? io_inputs_5 : _GEN_132; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_134 = 4'h6 == io_selects_4_0 ? io_inputs_6 : _GEN_133; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_135 = 4'h7 == io_selects_4_0 ? io_inputs_7 : _GEN_134; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_136 = 4'h8 == io_selects_4_0 ? io_inputs_8 : _GEN_135; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_137 = 4'h9 == io_selects_4_0 ? io_inputs_9 : _GEN_136; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_138 = 4'ha == io_selects_4_0 ? io_inputs_10 : _GEN_137; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_139 = 4'hb == io_selects_4_0 ? io_inputs_11 : _GEN_138; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_140 = 4'hc == io_selects_4_0 ? io_inputs_12 : _GEN_139; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_141 = 4'hd == io_selects_4_0 ? io_inputs_13 : _GEN_140; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_142 = 4'he == io_selects_4_0 ? io_inputs_14 : _GEN_141; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_143 = 4'hf == io_selects_4_0 ? io_inputs_15 : _GEN_142; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_145 = 4'h1 == io_selects_4_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_146 = 4'h2 == io_selects_4_1 ? io_inputs_2 : _GEN_145; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_147 = 4'h3 == io_selects_4_1 ? io_inputs_3 : _GEN_146; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_148 = 4'h4 == io_selects_4_1 ? io_inputs_4 : _GEN_147; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_149 = 4'h5 == io_selects_4_1 ? io_inputs_5 : _GEN_148; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_150 = 4'h6 == io_selects_4_1 ? io_inputs_6 : _GEN_149; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_151 = 4'h7 == io_selects_4_1 ? io_inputs_7 : _GEN_150; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_152 = 4'h8 == io_selects_4_1 ? io_inputs_8 : _GEN_151; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_153 = 4'h9 == io_selects_4_1 ? io_inputs_9 : _GEN_152; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_154 = 4'ha == io_selects_4_1 ? io_inputs_10 : _GEN_153; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_155 = 4'hb == io_selects_4_1 ? io_inputs_11 : _GEN_154; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_156 = 4'hc == io_selects_4_1 ? io_inputs_12 : _GEN_155; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_157 = 4'hd == io_selects_4_1 ? io_inputs_13 : _GEN_156; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_158 = 4'he == io_selects_4_1 ? io_inputs_14 : _GEN_157; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_159 = 4'hf == io_selects_4_1 ? io_inputs_15 : _GEN_158; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _T_486 = _GEN_143 + _GEN_159; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@56.4]
  assign _T_487 = _GEN_143 + _GEN_159; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@57.4]
  assign _T_489 = _GEN_143 * _GEN_159; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@58.4]
  assign _T_491 = _GEN_143 / _GEN_159; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@59.4]
  assign _T_492 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_493 = _T_492 ? _T_491 : 16'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_494 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_495 = _T_494 ? _T_489 : {{16'd0}, _T_493}; // @[Mux.scala 46:16:@63.4]
  assign _T_496 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_497 = _T_496 ? {{16'd0}, _T_487} : _T_495; // @[Mux.scala 46:16:@65.4]
  assign _T_498 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _T_499 = _T_498 ? {{16'd0}, _GEN_143} : _T_497; // @[Mux.scala 46:16:@67.4]
  assign _GEN_161 = 4'h1 == io_selects_5_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_162 = 4'h2 == io_selects_5_0 ? io_inputs_2 : _GEN_161; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_163 = 4'h3 == io_selects_5_0 ? io_inputs_3 : _GEN_162; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_164 = 4'h4 == io_selects_5_0 ? io_inputs_4 : _GEN_163; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_165 = 4'h5 == io_selects_5_0 ? io_inputs_5 : _GEN_164; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_166 = 4'h6 == io_selects_5_0 ? io_inputs_6 : _GEN_165; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_167 = 4'h7 == io_selects_5_0 ? io_inputs_7 : _GEN_166; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_168 = 4'h8 == io_selects_5_0 ? io_inputs_8 : _GEN_167; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_169 = 4'h9 == io_selects_5_0 ? io_inputs_9 : _GEN_168; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_170 = 4'ha == io_selects_5_0 ? io_inputs_10 : _GEN_169; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_171 = 4'hb == io_selects_5_0 ? io_inputs_11 : _GEN_170; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_172 = 4'hc == io_selects_5_0 ? io_inputs_12 : _GEN_171; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_173 = 4'hd == io_selects_5_0 ? io_inputs_13 : _GEN_172; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_174 = 4'he == io_selects_5_0 ? io_inputs_14 : _GEN_173; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_175 = 4'hf == io_selects_5_0 ? io_inputs_15 : _GEN_174; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_177 = 4'h1 == io_selects_5_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_178 = 4'h2 == io_selects_5_1 ? io_inputs_2 : _GEN_177; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_179 = 4'h3 == io_selects_5_1 ? io_inputs_3 : _GEN_178; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_180 = 4'h4 == io_selects_5_1 ? io_inputs_4 : _GEN_179; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_181 = 4'h5 == io_selects_5_1 ? io_inputs_5 : _GEN_180; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_182 = 4'h6 == io_selects_5_1 ? io_inputs_6 : _GEN_181; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_183 = 4'h7 == io_selects_5_1 ? io_inputs_7 : _GEN_182; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_184 = 4'h8 == io_selects_5_1 ? io_inputs_8 : _GEN_183; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_185 = 4'h9 == io_selects_5_1 ? io_inputs_9 : _GEN_184; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_186 = 4'ha == io_selects_5_1 ? io_inputs_10 : _GEN_185; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_187 = 4'hb == io_selects_5_1 ? io_inputs_11 : _GEN_186; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_188 = 4'hc == io_selects_5_1 ? io_inputs_12 : _GEN_187; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_189 = 4'hd == io_selects_5_1 ? io_inputs_13 : _GEN_188; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_190 = 4'he == io_selects_5_1 ? io_inputs_14 : _GEN_189; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_191 = 4'hf == io_selects_5_1 ? io_inputs_15 : _GEN_190; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _T_503 = _GEN_175 + _GEN_191; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@68.4]
  assign _T_504 = _GEN_175 + _GEN_191; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@69.4]
  assign _T_506 = _GEN_175 * _GEN_191; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@70.4]
  assign _T_508 = _GEN_175 / _GEN_191; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@71.4]
  assign _T_509 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_510 = _T_509 ? _T_508 : 16'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_511 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_512 = _T_511 ? _T_506 : {{16'd0}, _T_510}; // @[Mux.scala 46:16:@75.4]
  assign _T_513 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_514 = _T_513 ? {{16'd0}, _T_504} : _T_512; // @[Mux.scala 46:16:@77.4]
  assign _T_515 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _T_516 = _T_515 ? {{16'd0}, _GEN_175} : _T_514; // @[Mux.scala 46:16:@79.4]
  assign _GEN_193 = 4'h1 == io_selects_6_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_194 = 4'h2 == io_selects_6_0 ? io_inputs_2 : _GEN_193; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_195 = 4'h3 == io_selects_6_0 ? io_inputs_3 : _GEN_194; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_196 = 4'h4 == io_selects_6_0 ? io_inputs_4 : _GEN_195; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_197 = 4'h5 == io_selects_6_0 ? io_inputs_5 : _GEN_196; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_198 = 4'h6 == io_selects_6_0 ? io_inputs_6 : _GEN_197; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_199 = 4'h7 == io_selects_6_0 ? io_inputs_7 : _GEN_198; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_200 = 4'h8 == io_selects_6_0 ? io_inputs_8 : _GEN_199; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_201 = 4'h9 == io_selects_6_0 ? io_inputs_9 : _GEN_200; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_202 = 4'ha == io_selects_6_0 ? io_inputs_10 : _GEN_201; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_203 = 4'hb == io_selects_6_0 ? io_inputs_11 : _GEN_202; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_204 = 4'hc == io_selects_6_0 ? io_inputs_12 : _GEN_203; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_205 = 4'hd == io_selects_6_0 ? io_inputs_13 : _GEN_204; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_206 = 4'he == io_selects_6_0 ? io_inputs_14 : _GEN_205; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_207 = 4'hf == io_selects_6_0 ? io_inputs_15 : _GEN_206; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_209 = 4'h1 == io_selects_6_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_210 = 4'h2 == io_selects_6_1 ? io_inputs_2 : _GEN_209; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_211 = 4'h3 == io_selects_6_1 ? io_inputs_3 : _GEN_210; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_212 = 4'h4 == io_selects_6_1 ? io_inputs_4 : _GEN_211; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_213 = 4'h5 == io_selects_6_1 ? io_inputs_5 : _GEN_212; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_214 = 4'h6 == io_selects_6_1 ? io_inputs_6 : _GEN_213; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_215 = 4'h7 == io_selects_6_1 ? io_inputs_7 : _GEN_214; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_216 = 4'h8 == io_selects_6_1 ? io_inputs_8 : _GEN_215; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_217 = 4'h9 == io_selects_6_1 ? io_inputs_9 : _GEN_216; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_218 = 4'ha == io_selects_6_1 ? io_inputs_10 : _GEN_217; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_219 = 4'hb == io_selects_6_1 ? io_inputs_11 : _GEN_218; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_220 = 4'hc == io_selects_6_1 ? io_inputs_12 : _GEN_219; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_221 = 4'hd == io_selects_6_1 ? io_inputs_13 : _GEN_220; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_222 = 4'he == io_selects_6_1 ? io_inputs_14 : _GEN_221; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_223 = 4'hf == io_selects_6_1 ? io_inputs_15 : _GEN_222; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _T_520 = _GEN_207 + _GEN_223; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@80.4]
  assign _T_521 = _GEN_207 + _GEN_223; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@81.4]
  assign _T_523 = _GEN_207 * _GEN_223; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@82.4]
  assign _T_525 = _GEN_207 / _GEN_223; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@83.4]
  assign _T_526 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_527 = _T_526 ? _T_525 : 16'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_528 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_529 = _T_528 ? _T_523 : {{16'd0}, _T_527}; // @[Mux.scala 46:16:@87.4]
  assign _T_530 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_531 = _T_530 ? {{16'd0}, _T_521} : _T_529; // @[Mux.scala 46:16:@89.4]
  assign _T_532 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _T_533 = _T_532 ? {{16'd0}, _GEN_207} : _T_531; // @[Mux.scala 46:16:@91.4]
  assign _GEN_225 = 4'h1 == io_selects_7_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_226 = 4'h2 == io_selects_7_0 ? io_inputs_2 : _GEN_225; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_227 = 4'h3 == io_selects_7_0 ? io_inputs_3 : _GEN_226; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_228 = 4'h4 == io_selects_7_0 ? io_inputs_4 : _GEN_227; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_229 = 4'h5 == io_selects_7_0 ? io_inputs_5 : _GEN_228; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_230 = 4'h6 == io_selects_7_0 ? io_inputs_6 : _GEN_229; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_231 = 4'h7 == io_selects_7_0 ? io_inputs_7 : _GEN_230; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_232 = 4'h8 == io_selects_7_0 ? io_inputs_8 : _GEN_231; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_233 = 4'h9 == io_selects_7_0 ? io_inputs_9 : _GEN_232; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_234 = 4'ha == io_selects_7_0 ? io_inputs_10 : _GEN_233; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_235 = 4'hb == io_selects_7_0 ? io_inputs_11 : _GEN_234; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_236 = 4'hc == io_selects_7_0 ? io_inputs_12 : _GEN_235; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_237 = 4'hd == io_selects_7_0 ? io_inputs_13 : _GEN_236; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_238 = 4'he == io_selects_7_0 ? io_inputs_14 : _GEN_237; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_239 = 4'hf == io_selects_7_0 ? io_inputs_15 : _GEN_238; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_241 = 4'h1 == io_selects_7_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_242 = 4'h2 == io_selects_7_1 ? io_inputs_2 : _GEN_241; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_243 = 4'h3 == io_selects_7_1 ? io_inputs_3 : _GEN_242; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_244 = 4'h4 == io_selects_7_1 ? io_inputs_4 : _GEN_243; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_245 = 4'h5 == io_selects_7_1 ? io_inputs_5 : _GEN_244; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_246 = 4'h6 == io_selects_7_1 ? io_inputs_6 : _GEN_245; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_247 = 4'h7 == io_selects_7_1 ? io_inputs_7 : _GEN_246; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_248 = 4'h8 == io_selects_7_1 ? io_inputs_8 : _GEN_247; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_249 = 4'h9 == io_selects_7_1 ? io_inputs_9 : _GEN_248; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_250 = 4'ha == io_selects_7_1 ? io_inputs_10 : _GEN_249; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_251 = 4'hb == io_selects_7_1 ? io_inputs_11 : _GEN_250; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_252 = 4'hc == io_selects_7_1 ? io_inputs_12 : _GEN_251; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_253 = 4'hd == io_selects_7_1 ? io_inputs_13 : _GEN_252; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_254 = 4'he == io_selects_7_1 ? io_inputs_14 : _GEN_253; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_255 = 4'hf == io_selects_7_1 ? io_inputs_15 : _GEN_254; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _T_537 = _GEN_239 + _GEN_255; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@92.4]
  assign _T_538 = _GEN_239 + _GEN_255; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 32:53:@93.4]
  assign _T_540 = _GEN_239 * _GEN_255; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 33:58:@94.4]
  assign _T_542 = _GEN_239 / _GEN_255; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 34:56:@95.4]
  assign _T_543 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_544 = _T_543 ? _T_542 : 16'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_545 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_546 = _T_545 ? _T_540 : {{16'd0}, _T_544}; // @[Mux.scala 46:16:@99.4]
  assign _T_547 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_548 = _T_547 ? {{16'd0}, _T_538} : _T_546; // @[Mux.scala 46:16:@101.4]
  assign _T_549 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign _T_550 = _T_549 ? {{16'd0}, _GEN_239} : _T_548; // @[Mux.scala 46:16:@103.4]
  assign io_outputs_0 = _T_431[15:0]; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 23:14:@104.4]
  assign io_outputs_1 = _T_448[15:0]; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 23:14:@105.4]
  assign io_outputs_2 = _T_465[15:0]; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 23:14:@106.4]
  assign io_outputs_3 = _T_482[15:0]; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 23:14:@107.4]
  assign io_outputs_4 = _T_499[15:0]; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 23:14:@108.4]
  assign io_outputs_5 = _T_516[15:0]; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 23:14:@109.4]
  assign io_outputs_6 = _T_533[15:0]; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 23:14:@110.4]
  assign io_outputs_7 = _T_550[15:0]; // @[MuxTest_width_16_inputs_16_outputs_8_pipeline_0s.scala 23:14:@111.4]
endmodule
