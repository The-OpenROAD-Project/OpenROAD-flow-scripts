(* blackbox *) module ASYNC_DFFHx1_ASAP7_75t_SL (QN, D, RESET, SET, CLK);
	output QN;
	input D, RESET, SET, CLK;
endmodule
(* blackbox *) module DFFHQNx1_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQNx2_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQNx3_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFHQx4_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx1_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx2_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQNx3_ASAP7_75t_SL (QN, D, CLK);
	output QN;
	input D, CLK;
endmodule
(* blackbox *) module DFFLQx4_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx1_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx2_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DHLx3_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx1_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx2_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module DLLx3_ASAP7_75t_SL (Q, D, CLK);
	output Q;
	input D, CLK;
endmodule
(* blackbox *) module ICGx1_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx2_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx2p67DC_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx3_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx4DC_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx4_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx5_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx5p33DC_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx6p67DC_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module ICGx8DC_ASAP7_75t_SL (GCLK, ENA, SE, CLK);
	output GCLK;
	input ENA, SE, CLK;
endmodule
(* blackbox *) module SDFHx1_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx2_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx3_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFHx4_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx1_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx2_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx3_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
(* blackbox *) module SDFLx4_ASAP7_75t_SL (QN, D, SE, SI, CLK);
	output QN;
	input D, SE, SI, CLK;
endmodule
