module MockArray (clock,
    io_lsbs_0,
    io_lsbs_1,
    io_lsbs_10,
    io_lsbs_11,
    io_lsbs_12,
    io_lsbs_13,
    io_lsbs_14,
    io_lsbs_15,
    io_lsbs_16,
    io_lsbs_17,
    io_lsbs_18,
    io_lsbs_19,
    io_lsbs_2,
    io_lsbs_20,
    io_lsbs_21,
    io_lsbs_22,
    io_lsbs_23,
    io_lsbs_24,
    io_lsbs_25,
    io_lsbs_26,
    io_lsbs_27,
    io_lsbs_28,
    io_lsbs_29,
    io_lsbs_3,
    io_lsbs_30,
    io_lsbs_31,
    io_lsbs_32,
    io_lsbs_33,
    io_lsbs_34,
    io_lsbs_35,
    io_lsbs_36,
    io_lsbs_37,
    io_lsbs_38,
    io_lsbs_39,
    io_lsbs_4,
    io_lsbs_40,
    io_lsbs_41,
    io_lsbs_42,
    io_lsbs_43,
    io_lsbs_44,
    io_lsbs_45,
    io_lsbs_46,
    io_lsbs_47,
    io_lsbs_48,
    io_lsbs_49,
    io_lsbs_5,
    io_lsbs_50,
    io_lsbs_51,
    io_lsbs_52,
    io_lsbs_53,
    io_lsbs_54,
    io_lsbs_55,
    io_lsbs_56,
    io_lsbs_57,
    io_lsbs_58,
    io_lsbs_59,
    io_lsbs_6,
    io_lsbs_60,
    io_lsbs_61,
    io_lsbs_62,
    io_lsbs_63,
    io_lsbs_7,
    io_lsbs_8,
    io_lsbs_9,
    reset,
    io_ins_down_0,
    io_ins_down_1,
    io_ins_down_2,
    io_ins_down_3,
    io_ins_down_4,
    io_ins_down_5,
    io_ins_down_6,
    io_ins_down_7,
    io_ins_left_0,
    io_ins_left_1,
    io_ins_left_2,
    io_ins_left_3,
    io_ins_left_4,
    io_ins_left_5,
    io_ins_left_6,
    io_ins_left_7,
    io_ins_right_0,
    io_ins_right_1,
    io_ins_right_2,
    io_ins_right_3,
    io_ins_right_4,
    io_ins_right_5,
    io_ins_right_6,
    io_ins_right_7,
    io_ins_up_0,
    io_ins_up_1,
    io_ins_up_2,
    io_ins_up_3,
    io_ins_up_4,
    io_ins_up_5,
    io_ins_up_6,
    io_ins_up_7,
    io_outs_down_0,
    io_outs_down_1,
    io_outs_down_2,
    io_outs_down_3,
    io_outs_down_4,
    io_outs_down_5,
    io_outs_down_6,
    io_outs_down_7,
    io_outs_left_0,
    io_outs_left_1,
    io_outs_left_2,
    io_outs_left_3,
    io_outs_left_4,
    io_outs_left_5,
    io_outs_left_6,
    io_outs_left_7,
    io_outs_right_0,
    io_outs_right_1,
    io_outs_right_2,
    io_outs_right_3,
    io_outs_right_4,
    io_outs_right_5,
    io_outs_right_6,
    io_outs_right_7,
    io_outs_up_0,
    io_outs_up_1,
    io_outs_up_2,
    io_outs_up_3,
    io_outs_up_4,
    io_outs_up_5,
    io_outs_up_6,
    io_outs_up_7);
 input clock;
 output io_lsbs_0;
 output io_lsbs_1;
 output io_lsbs_10;
 output io_lsbs_11;
 output io_lsbs_12;
 output io_lsbs_13;
 output io_lsbs_14;
 output io_lsbs_15;
 output io_lsbs_16;
 output io_lsbs_17;
 output io_lsbs_18;
 output io_lsbs_19;
 output io_lsbs_2;
 output io_lsbs_20;
 output io_lsbs_21;
 output io_lsbs_22;
 output io_lsbs_23;
 output io_lsbs_24;
 output io_lsbs_25;
 output io_lsbs_26;
 output io_lsbs_27;
 output io_lsbs_28;
 output io_lsbs_29;
 output io_lsbs_3;
 output io_lsbs_30;
 output io_lsbs_31;
 output io_lsbs_32;
 output io_lsbs_33;
 output io_lsbs_34;
 output io_lsbs_35;
 output io_lsbs_36;
 output io_lsbs_37;
 output io_lsbs_38;
 output io_lsbs_39;
 output io_lsbs_4;
 output io_lsbs_40;
 output io_lsbs_41;
 output io_lsbs_42;
 output io_lsbs_43;
 output io_lsbs_44;
 output io_lsbs_45;
 output io_lsbs_46;
 output io_lsbs_47;
 output io_lsbs_48;
 output io_lsbs_49;
 output io_lsbs_5;
 output io_lsbs_50;
 output io_lsbs_51;
 output io_lsbs_52;
 output io_lsbs_53;
 output io_lsbs_54;
 output io_lsbs_55;
 output io_lsbs_56;
 output io_lsbs_57;
 output io_lsbs_58;
 output io_lsbs_59;
 output io_lsbs_6;
 output io_lsbs_60;
 output io_lsbs_61;
 output io_lsbs_62;
 output io_lsbs_63;
 output io_lsbs_7;
 output io_lsbs_8;
 output io_lsbs_9;
 input reset;
 input [63:0] io_ins_down_0;
 input [63:0] io_ins_down_1;
 input [63:0] io_ins_down_2;
 input [63:0] io_ins_down_3;
 input [63:0] io_ins_down_4;
 input [63:0] io_ins_down_5;
 input [63:0] io_ins_down_6;
 input [63:0] io_ins_down_7;
 input [63:0] io_ins_left_0;
 input [63:0] io_ins_left_1;
 input [63:0] io_ins_left_2;
 input [63:0] io_ins_left_3;
 input [63:0] io_ins_left_4;
 input [63:0] io_ins_left_5;
 input [63:0] io_ins_left_6;
 input [63:0] io_ins_left_7;
 input [63:0] io_ins_right_0;
 input [63:0] io_ins_right_1;
 input [63:0] io_ins_right_2;
 input [63:0] io_ins_right_3;
 input [63:0] io_ins_right_4;
 input [63:0] io_ins_right_5;
 input [63:0] io_ins_right_6;
 input [63:0] io_ins_right_7;
 input [63:0] io_ins_up_0;
 input [63:0] io_ins_up_1;
 input [63:0] io_ins_up_2;
 input [63:0] io_ins_up_3;
 input [63:0] io_ins_up_4;
 input [63:0] io_ins_up_5;
 input [63:0] io_ins_up_6;
 input [63:0] io_ins_up_7;
 output [63:0] io_outs_down_0;
 output [63:0] io_outs_down_1;
 output [63:0] io_outs_down_2;
 output [63:0] io_outs_down_3;
 output [63:0] io_outs_down_4;
 output [63:0] io_outs_down_5;
 output [63:0] io_outs_down_6;
 output [63:0] io_outs_down_7;
 output [63:0] io_outs_left_0;
 output [63:0] io_outs_left_1;
 output [63:0] io_outs_left_2;
 output [63:0] io_outs_left_3;
 output [63:0] io_outs_left_4;
 output [63:0] io_outs_left_5;
 output [63:0] io_outs_left_6;
 output [63:0] io_outs_left_7;
 output [63:0] io_outs_right_0;
 output [63:0] io_outs_right_1;
 output [63:0] io_outs_right_2;
 output [63:0] io_outs_right_3;
 output [63:0] io_outs_right_4;
 output [63:0] io_outs_right_5;
 output [63:0] io_outs_right_6;
 output [63:0] io_outs_right_7;
 output [63:0] io_outs_up_0;
 output [63:0] io_outs_up_1;
 output [63:0] io_outs_up_2;
 output [63:0] io_outs_up_3;
 output [63:0] io_outs_up_4;
 output [63:0] io_outs_up_5;
 output [63:0] io_outs_up_6;
 output [63:0] io_outs_up_7;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire clock_regs;
 wire \ces_0_0_io_ins_down[0] ;
 wire \ces_0_0_io_ins_down[10] ;
 wire \ces_0_0_io_ins_down[11] ;
 wire \ces_0_0_io_ins_down[12] ;
 wire \ces_0_0_io_ins_down[13] ;
 wire \ces_0_0_io_ins_down[14] ;
 wire \ces_0_0_io_ins_down[15] ;
 wire \ces_0_0_io_ins_down[16] ;
 wire \ces_0_0_io_ins_down[17] ;
 wire \ces_0_0_io_ins_down[18] ;
 wire \ces_0_0_io_ins_down[19] ;
 wire \ces_0_0_io_ins_down[1] ;
 wire \ces_0_0_io_ins_down[20] ;
 wire \ces_0_0_io_ins_down[21] ;
 wire \ces_0_0_io_ins_down[22] ;
 wire \ces_0_0_io_ins_down[23] ;
 wire \ces_0_0_io_ins_down[24] ;
 wire \ces_0_0_io_ins_down[25] ;
 wire \ces_0_0_io_ins_down[26] ;
 wire \ces_0_0_io_ins_down[27] ;
 wire \ces_0_0_io_ins_down[28] ;
 wire \ces_0_0_io_ins_down[29] ;
 wire \ces_0_0_io_ins_down[2] ;
 wire \ces_0_0_io_ins_down[30] ;
 wire \ces_0_0_io_ins_down[31] ;
 wire \ces_0_0_io_ins_down[32] ;
 wire \ces_0_0_io_ins_down[33] ;
 wire \ces_0_0_io_ins_down[34] ;
 wire \ces_0_0_io_ins_down[35] ;
 wire \ces_0_0_io_ins_down[36] ;
 wire \ces_0_0_io_ins_down[37] ;
 wire \ces_0_0_io_ins_down[38] ;
 wire \ces_0_0_io_ins_down[39] ;
 wire \ces_0_0_io_ins_down[3] ;
 wire \ces_0_0_io_ins_down[40] ;
 wire \ces_0_0_io_ins_down[41] ;
 wire \ces_0_0_io_ins_down[42] ;
 wire \ces_0_0_io_ins_down[43] ;
 wire \ces_0_0_io_ins_down[44] ;
 wire \ces_0_0_io_ins_down[45] ;
 wire \ces_0_0_io_ins_down[46] ;
 wire \ces_0_0_io_ins_down[47] ;
 wire \ces_0_0_io_ins_down[48] ;
 wire \ces_0_0_io_ins_down[49] ;
 wire \ces_0_0_io_ins_down[4] ;
 wire \ces_0_0_io_ins_down[50] ;
 wire \ces_0_0_io_ins_down[51] ;
 wire \ces_0_0_io_ins_down[52] ;
 wire \ces_0_0_io_ins_down[53] ;
 wire \ces_0_0_io_ins_down[54] ;
 wire \ces_0_0_io_ins_down[55] ;
 wire \ces_0_0_io_ins_down[56] ;
 wire \ces_0_0_io_ins_down[57] ;
 wire \ces_0_0_io_ins_down[58] ;
 wire \ces_0_0_io_ins_down[59] ;
 wire \ces_0_0_io_ins_down[5] ;
 wire \ces_0_0_io_ins_down[60] ;
 wire \ces_0_0_io_ins_down[61] ;
 wire \ces_0_0_io_ins_down[62] ;
 wire \ces_0_0_io_ins_down[63] ;
 wire \ces_0_0_io_ins_down[6] ;
 wire \ces_0_0_io_ins_down[7] ;
 wire \ces_0_0_io_ins_down[8] ;
 wire \ces_0_0_io_ins_down[9] ;
 wire \ces_0_0_io_ins_left[0] ;
 wire \ces_0_0_io_ins_left[10] ;
 wire \ces_0_0_io_ins_left[11] ;
 wire \ces_0_0_io_ins_left[12] ;
 wire \ces_0_0_io_ins_left[13] ;
 wire \ces_0_0_io_ins_left[14] ;
 wire \ces_0_0_io_ins_left[15] ;
 wire \ces_0_0_io_ins_left[16] ;
 wire \ces_0_0_io_ins_left[17] ;
 wire \ces_0_0_io_ins_left[18] ;
 wire \ces_0_0_io_ins_left[19] ;
 wire \ces_0_0_io_ins_left[1] ;
 wire \ces_0_0_io_ins_left[20] ;
 wire \ces_0_0_io_ins_left[21] ;
 wire \ces_0_0_io_ins_left[22] ;
 wire \ces_0_0_io_ins_left[23] ;
 wire \ces_0_0_io_ins_left[24] ;
 wire \ces_0_0_io_ins_left[25] ;
 wire \ces_0_0_io_ins_left[26] ;
 wire \ces_0_0_io_ins_left[27] ;
 wire \ces_0_0_io_ins_left[28] ;
 wire \ces_0_0_io_ins_left[29] ;
 wire \ces_0_0_io_ins_left[2] ;
 wire \ces_0_0_io_ins_left[30] ;
 wire \ces_0_0_io_ins_left[31] ;
 wire \ces_0_0_io_ins_left[32] ;
 wire \ces_0_0_io_ins_left[33] ;
 wire \ces_0_0_io_ins_left[34] ;
 wire \ces_0_0_io_ins_left[35] ;
 wire \ces_0_0_io_ins_left[36] ;
 wire \ces_0_0_io_ins_left[37] ;
 wire \ces_0_0_io_ins_left[38] ;
 wire \ces_0_0_io_ins_left[39] ;
 wire \ces_0_0_io_ins_left[3] ;
 wire \ces_0_0_io_ins_left[40] ;
 wire \ces_0_0_io_ins_left[41] ;
 wire \ces_0_0_io_ins_left[42] ;
 wire \ces_0_0_io_ins_left[43] ;
 wire \ces_0_0_io_ins_left[44] ;
 wire \ces_0_0_io_ins_left[45] ;
 wire \ces_0_0_io_ins_left[46] ;
 wire \ces_0_0_io_ins_left[47] ;
 wire \ces_0_0_io_ins_left[48] ;
 wire \ces_0_0_io_ins_left[49] ;
 wire \ces_0_0_io_ins_left[4] ;
 wire \ces_0_0_io_ins_left[50] ;
 wire \ces_0_0_io_ins_left[51] ;
 wire \ces_0_0_io_ins_left[52] ;
 wire \ces_0_0_io_ins_left[53] ;
 wire \ces_0_0_io_ins_left[54] ;
 wire \ces_0_0_io_ins_left[55] ;
 wire \ces_0_0_io_ins_left[56] ;
 wire \ces_0_0_io_ins_left[57] ;
 wire \ces_0_0_io_ins_left[58] ;
 wire \ces_0_0_io_ins_left[59] ;
 wire \ces_0_0_io_ins_left[5] ;
 wire \ces_0_0_io_ins_left[60] ;
 wire \ces_0_0_io_ins_left[61] ;
 wire \ces_0_0_io_ins_left[62] ;
 wire \ces_0_0_io_ins_left[63] ;
 wire \ces_0_0_io_ins_left[6] ;
 wire \ces_0_0_io_ins_left[7] ;
 wire \ces_0_0_io_ins_left[8] ;
 wire \ces_0_0_io_ins_left[9] ;
 wire ces_0_0_io_lsbOuts_0;
 wire ces_0_0_io_lsbOuts_1;
 wire ces_0_0_io_lsbOuts_2;
 wire ces_0_0_io_lsbOuts_3;
 wire ces_0_0_io_lsbOuts_4;
 wire ces_0_0_io_lsbOuts_5;
 wire ces_0_0_io_lsbOuts_6;
 wire ces_0_0_io_lsbOuts_7;
 wire \ces_0_0_io_outs_right[0] ;
 wire \ces_0_0_io_outs_right[10] ;
 wire \ces_0_0_io_outs_right[11] ;
 wire \ces_0_0_io_outs_right[12] ;
 wire \ces_0_0_io_outs_right[13] ;
 wire \ces_0_0_io_outs_right[14] ;
 wire \ces_0_0_io_outs_right[15] ;
 wire \ces_0_0_io_outs_right[16] ;
 wire \ces_0_0_io_outs_right[17] ;
 wire \ces_0_0_io_outs_right[18] ;
 wire \ces_0_0_io_outs_right[19] ;
 wire \ces_0_0_io_outs_right[1] ;
 wire \ces_0_0_io_outs_right[20] ;
 wire \ces_0_0_io_outs_right[21] ;
 wire \ces_0_0_io_outs_right[22] ;
 wire \ces_0_0_io_outs_right[23] ;
 wire \ces_0_0_io_outs_right[24] ;
 wire \ces_0_0_io_outs_right[25] ;
 wire \ces_0_0_io_outs_right[26] ;
 wire \ces_0_0_io_outs_right[27] ;
 wire \ces_0_0_io_outs_right[28] ;
 wire \ces_0_0_io_outs_right[29] ;
 wire \ces_0_0_io_outs_right[2] ;
 wire \ces_0_0_io_outs_right[30] ;
 wire \ces_0_0_io_outs_right[31] ;
 wire \ces_0_0_io_outs_right[32] ;
 wire \ces_0_0_io_outs_right[33] ;
 wire \ces_0_0_io_outs_right[34] ;
 wire \ces_0_0_io_outs_right[35] ;
 wire \ces_0_0_io_outs_right[36] ;
 wire \ces_0_0_io_outs_right[37] ;
 wire \ces_0_0_io_outs_right[38] ;
 wire \ces_0_0_io_outs_right[39] ;
 wire \ces_0_0_io_outs_right[3] ;
 wire \ces_0_0_io_outs_right[40] ;
 wire \ces_0_0_io_outs_right[41] ;
 wire \ces_0_0_io_outs_right[42] ;
 wire \ces_0_0_io_outs_right[43] ;
 wire \ces_0_0_io_outs_right[44] ;
 wire \ces_0_0_io_outs_right[45] ;
 wire \ces_0_0_io_outs_right[46] ;
 wire \ces_0_0_io_outs_right[47] ;
 wire \ces_0_0_io_outs_right[48] ;
 wire \ces_0_0_io_outs_right[49] ;
 wire \ces_0_0_io_outs_right[4] ;
 wire \ces_0_0_io_outs_right[50] ;
 wire \ces_0_0_io_outs_right[51] ;
 wire \ces_0_0_io_outs_right[52] ;
 wire \ces_0_0_io_outs_right[53] ;
 wire \ces_0_0_io_outs_right[54] ;
 wire \ces_0_0_io_outs_right[55] ;
 wire \ces_0_0_io_outs_right[56] ;
 wire \ces_0_0_io_outs_right[57] ;
 wire \ces_0_0_io_outs_right[58] ;
 wire \ces_0_0_io_outs_right[59] ;
 wire \ces_0_0_io_outs_right[5] ;
 wire \ces_0_0_io_outs_right[60] ;
 wire \ces_0_0_io_outs_right[61] ;
 wire \ces_0_0_io_outs_right[62] ;
 wire \ces_0_0_io_outs_right[63] ;
 wire \ces_0_0_io_outs_right[6] ;
 wire \ces_0_0_io_outs_right[7] ;
 wire \ces_0_0_io_outs_right[8] ;
 wire \ces_0_0_io_outs_right[9] ;
 wire \ces_0_0_io_outs_up[0] ;
 wire \ces_0_0_io_outs_up[10] ;
 wire \ces_0_0_io_outs_up[11] ;
 wire \ces_0_0_io_outs_up[12] ;
 wire \ces_0_0_io_outs_up[13] ;
 wire \ces_0_0_io_outs_up[14] ;
 wire \ces_0_0_io_outs_up[15] ;
 wire \ces_0_0_io_outs_up[16] ;
 wire \ces_0_0_io_outs_up[17] ;
 wire \ces_0_0_io_outs_up[18] ;
 wire \ces_0_0_io_outs_up[19] ;
 wire \ces_0_0_io_outs_up[1] ;
 wire \ces_0_0_io_outs_up[20] ;
 wire \ces_0_0_io_outs_up[21] ;
 wire \ces_0_0_io_outs_up[22] ;
 wire \ces_0_0_io_outs_up[23] ;
 wire \ces_0_0_io_outs_up[24] ;
 wire \ces_0_0_io_outs_up[25] ;
 wire \ces_0_0_io_outs_up[26] ;
 wire \ces_0_0_io_outs_up[27] ;
 wire \ces_0_0_io_outs_up[28] ;
 wire \ces_0_0_io_outs_up[29] ;
 wire \ces_0_0_io_outs_up[2] ;
 wire \ces_0_0_io_outs_up[30] ;
 wire \ces_0_0_io_outs_up[31] ;
 wire \ces_0_0_io_outs_up[32] ;
 wire \ces_0_0_io_outs_up[33] ;
 wire \ces_0_0_io_outs_up[34] ;
 wire \ces_0_0_io_outs_up[35] ;
 wire \ces_0_0_io_outs_up[36] ;
 wire \ces_0_0_io_outs_up[37] ;
 wire \ces_0_0_io_outs_up[38] ;
 wire \ces_0_0_io_outs_up[39] ;
 wire \ces_0_0_io_outs_up[3] ;
 wire \ces_0_0_io_outs_up[40] ;
 wire \ces_0_0_io_outs_up[41] ;
 wire \ces_0_0_io_outs_up[42] ;
 wire \ces_0_0_io_outs_up[43] ;
 wire \ces_0_0_io_outs_up[44] ;
 wire \ces_0_0_io_outs_up[45] ;
 wire \ces_0_0_io_outs_up[46] ;
 wire \ces_0_0_io_outs_up[47] ;
 wire \ces_0_0_io_outs_up[48] ;
 wire \ces_0_0_io_outs_up[49] ;
 wire \ces_0_0_io_outs_up[4] ;
 wire \ces_0_0_io_outs_up[50] ;
 wire \ces_0_0_io_outs_up[51] ;
 wire \ces_0_0_io_outs_up[52] ;
 wire \ces_0_0_io_outs_up[53] ;
 wire \ces_0_0_io_outs_up[54] ;
 wire \ces_0_0_io_outs_up[55] ;
 wire \ces_0_0_io_outs_up[56] ;
 wire \ces_0_0_io_outs_up[57] ;
 wire \ces_0_0_io_outs_up[58] ;
 wire \ces_0_0_io_outs_up[59] ;
 wire \ces_0_0_io_outs_up[5] ;
 wire \ces_0_0_io_outs_up[60] ;
 wire \ces_0_0_io_outs_up[61] ;
 wire \ces_0_0_io_outs_up[62] ;
 wire \ces_0_0_io_outs_up[63] ;
 wire \ces_0_0_io_outs_up[6] ;
 wire \ces_0_0_io_outs_up[7] ;
 wire \ces_0_0_io_outs_up[8] ;
 wire \ces_0_0_io_outs_up[9] ;
 wire \ces_0_1_io_ins_down[0] ;
 wire \ces_0_1_io_ins_down[10] ;
 wire \ces_0_1_io_ins_down[11] ;
 wire \ces_0_1_io_ins_down[12] ;
 wire \ces_0_1_io_ins_down[13] ;
 wire \ces_0_1_io_ins_down[14] ;
 wire \ces_0_1_io_ins_down[15] ;
 wire \ces_0_1_io_ins_down[16] ;
 wire \ces_0_1_io_ins_down[17] ;
 wire \ces_0_1_io_ins_down[18] ;
 wire \ces_0_1_io_ins_down[19] ;
 wire \ces_0_1_io_ins_down[1] ;
 wire \ces_0_1_io_ins_down[20] ;
 wire \ces_0_1_io_ins_down[21] ;
 wire \ces_0_1_io_ins_down[22] ;
 wire \ces_0_1_io_ins_down[23] ;
 wire \ces_0_1_io_ins_down[24] ;
 wire \ces_0_1_io_ins_down[25] ;
 wire \ces_0_1_io_ins_down[26] ;
 wire \ces_0_1_io_ins_down[27] ;
 wire \ces_0_1_io_ins_down[28] ;
 wire \ces_0_1_io_ins_down[29] ;
 wire \ces_0_1_io_ins_down[2] ;
 wire \ces_0_1_io_ins_down[30] ;
 wire \ces_0_1_io_ins_down[31] ;
 wire \ces_0_1_io_ins_down[32] ;
 wire \ces_0_1_io_ins_down[33] ;
 wire \ces_0_1_io_ins_down[34] ;
 wire \ces_0_1_io_ins_down[35] ;
 wire \ces_0_1_io_ins_down[36] ;
 wire \ces_0_1_io_ins_down[37] ;
 wire \ces_0_1_io_ins_down[38] ;
 wire \ces_0_1_io_ins_down[39] ;
 wire \ces_0_1_io_ins_down[3] ;
 wire \ces_0_1_io_ins_down[40] ;
 wire \ces_0_1_io_ins_down[41] ;
 wire \ces_0_1_io_ins_down[42] ;
 wire \ces_0_1_io_ins_down[43] ;
 wire \ces_0_1_io_ins_down[44] ;
 wire \ces_0_1_io_ins_down[45] ;
 wire \ces_0_1_io_ins_down[46] ;
 wire \ces_0_1_io_ins_down[47] ;
 wire \ces_0_1_io_ins_down[48] ;
 wire \ces_0_1_io_ins_down[49] ;
 wire \ces_0_1_io_ins_down[4] ;
 wire \ces_0_1_io_ins_down[50] ;
 wire \ces_0_1_io_ins_down[51] ;
 wire \ces_0_1_io_ins_down[52] ;
 wire \ces_0_1_io_ins_down[53] ;
 wire \ces_0_1_io_ins_down[54] ;
 wire \ces_0_1_io_ins_down[55] ;
 wire \ces_0_1_io_ins_down[56] ;
 wire \ces_0_1_io_ins_down[57] ;
 wire \ces_0_1_io_ins_down[58] ;
 wire \ces_0_1_io_ins_down[59] ;
 wire \ces_0_1_io_ins_down[5] ;
 wire \ces_0_1_io_ins_down[60] ;
 wire \ces_0_1_io_ins_down[61] ;
 wire \ces_0_1_io_ins_down[62] ;
 wire \ces_0_1_io_ins_down[63] ;
 wire \ces_0_1_io_ins_down[6] ;
 wire \ces_0_1_io_ins_down[7] ;
 wire \ces_0_1_io_ins_down[8] ;
 wire \ces_0_1_io_ins_down[9] ;
 wire \ces_0_1_io_ins_left[0] ;
 wire \ces_0_1_io_ins_left[10] ;
 wire \ces_0_1_io_ins_left[11] ;
 wire \ces_0_1_io_ins_left[12] ;
 wire \ces_0_1_io_ins_left[13] ;
 wire \ces_0_1_io_ins_left[14] ;
 wire \ces_0_1_io_ins_left[15] ;
 wire \ces_0_1_io_ins_left[16] ;
 wire \ces_0_1_io_ins_left[17] ;
 wire \ces_0_1_io_ins_left[18] ;
 wire \ces_0_1_io_ins_left[19] ;
 wire \ces_0_1_io_ins_left[1] ;
 wire \ces_0_1_io_ins_left[20] ;
 wire \ces_0_1_io_ins_left[21] ;
 wire \ces_0_1_io_ins_left[22] ;
 wire \ces_0_1_io_ins_left[23] ;
 wire \ces_0_1_io_ins_left[24] ;
 wire \ces_0_1_io_ins_left[25] ;
 wire \ces_0_1_io_ins_left[26] ;
 wire \ces_0_1_io_ins_left[27] ;
 wire \ces_0_1_io_ins_left[28] ;
 wire \ces_0_1_io_ins_left[29] ;
 wire \ces_0_1_io_ins_left[2] ;
 wire \ces_0_1_io_ins_left[30] ;
 wire \ces_0_1_io_ins_left[31] ;
 wire \ces_0_1_io_ins_left[32] ;
 wire \ces_0_1_io_ins_left[33] ;
 wire \ces_0_1_io_ins_left[34] ;
 wire \ces_0_1_io_ins_left[35] ;
 wire \ces_0_1_io_ins_left[36] ;
 wire \ces_0_1_io_ins_left[37] ;
 wire \ces_0_1_io_ins_left[38] ;
 wire \ces_0_1_io_ins_left[39] ;
 wire \ces_0_1_io_ins_left[3] ;
 wire \ces_0_1_io_ins_left[40] ;
 wire \ces_0_1_io_ins_left[41] ;
 wire \ces_0_1_io_ins_left[42] ;
 wire \ces_0_1_io_ins_left[43] ;
 wire \ces_0_1_io_ins_left[44] ;
 wire \ces_0_1_io_ins_left[45] ;
 wire \ces_0_1_io_ins_left[46] ;
 wire \ces_0_1_io_ins_left[47] ;
 wire \ces_0_1_io_ins_left[48] ;
 wire \ces_0_1_io_ins_left[49] ;
 wire \ces_0_1_io_ins_left[4] ;
 wire \ces_0_1_io_ins_left[50] ;
 wire \ces_0_1_io_ins_left[51] ;
 wire \ces_0_1_io_ins_left[52] ;
 wire \ces_0_1_io_ins_left[53] ;
 wire \ces_0_1_io_ins_left[54] ;
 wire \ces_0_1_io_ins_left[55] ;
 wire \ces_0_1_io_ins_left[56] ;
 wire \ces_0_1_io_ins_left[57] ;
 wire \ces_0_1_io_ins_left[58] ;
 wire \ces_0_1_io_ins_left[59] ;
 wire \ces_0_1_io_ins_left[5] ;
 wire \ces_0_1_io_ins_left[60] ;
 wire \ces_0_1_io_ins_left[61] ;
 wire \ces_0_1_io_ins_left[62] ;
 wire \ces_0_1_io_ins_left[63] ;
 wire \ces_0_1_io_ins_left[6] ;
 wire \ces_0_1_io_ins_left[7] ;
 wire \ces_0_1_io_ins_left[8] ;
 wire \ces_0_1_io_ins_left[9] ;
 wire ces_0_1_io_lsbOuts_0;
 wire ces_0_1_io_lsbOuts_1;
 wire ces_0_1_io_lsbOuts_2;
 wire ces_0_1_io_lsbOuts_3;
 wire ces_0_1_io_lsbOuts_4;
 wire ces_0_1_io_lsbOuts_5;
 wire ces_0_1_io_lsbOuts_6;
 wire ces_0_1_io_lsbOuts_7;
 wire \ces_0_1_io_outs_right[0] ;
 wire \ces_0_1_io_outs_right[10] ;
 wire \ces_0_1_io_outs_right[11] ;
 wire \ces_0_1_io_outs_right[12] ;
 wire \ces_0_1_io_outs_right[13] ;
 wire \ces_0_1_io_outs_right[14] ;
 wire \ces_0_1_io_outs_right[15] ;
 wire \ces_0_1_io_outs_right[16] ;
 wire \ces_0_1_io_outs_right[17] ;
 wire \ces_0_1_io_outs_right[18] ;
 wire \ces_0_1_io_outs_right[19] ;
 wire \ces_0_1_io_outs_right[1] ;
 wire \ces_0_1_io_outs_right[20] ;
 wire \ces_0_1_io_outs_right[21] ;
 wire \ces_0_1_io_outs_right[22] ;
 wire \ces_0_1_io_outs_right[23] ;
 wire \ces_0_1_io_outs_right[24] ;
 wire \ces_0_1_io_outs_right[25] ;
 wire \ces_0_1_io_outs_right[26] ;
 wire \ces_0_1_io_outs_right[27] ;
 wire \ces_0_1_io_outs_right[28] ;
 wire \ces_0_1_io_outs_right[29] ;
 wire \ces_0_1_io_outs_right[2] ;
 wire \ces_0_1_io_outs_right[30] ;
 wire \ces_0_1_io_outs_right[31] ;
 wire \ces_0_1_io_outs_right[32] ;
 wire \ces_0_1_io_outs_right[33] ;
 wire \ces_0_1_io_outs_right[34] ;
 wire \ces_0_1_io_outs_right[35] ;
 wire \ces_0_1_io_outs_right[36] ;
 wire \ces_0_1_io_outs_right[37] ;
 wire \ces_0_1_io_outs_right[38] ;
 wire \ces_0_1_io_outs_right[39] ;
 wire \ces_0_1_io_outs_right[3] ;
 wire \ces_0_1_io_outs_right[40] ;
 wire \ces_0_1_io_outs_right[41] ;
 wire \ces_0_1_io_outs_right[42] ;
 wire \ces_0_1_io_outs_right[43] ;
 wire \ces_0_1_io_outs_right[44] ;
 wire \ces_0_1_io_outs_right[45] ;
 wire \ces_0_1_io_outs_right[46] ;
 wire \ces_0_1_io_outs_right[47] ;
 wire \ces_0_1_io_outs_right[48] ;
 wire \ces_0_1_io_outs_right[49] ;
 wire \ces_0_1_io_outs_right[4] ;
 wire \ces_0_1_io_outs_right[50] ;
 wire \ces_0_1_io_outs_right[51] ;
 wire \ces_0_1_io_outs_right[52] ;
 wire \ces_0_1_io_outs_right[53] ;
 wire \ces_0_1_io_outs_right[54] ;
 wire \ces_0_1_io_outs_right[55] ;
 wire \ces_0_1_io_outs_right[56] ;
 wire \ces_0_1_io_outs_right[57] ;
 wire \ces_0_1_io_outs_right[58] ;
 wire \ces_0_1_io_outs_right[59] ;
 wire \ces_0_1_io_outs_right[5] ;
 wire \ces_0_1_io_outs_right[60] ;
 wire \ces_0_1_io_outs_right[61] ;
 wire \ces_0_1_io_outs_right[62] ;
 wire \ces_0_1_io_outs_right[63] ;
 wire \ces_0_1_io_outs_right[6] ;
 wire \ces_0_1_io_outs_right[7] ;
 wire \ces_0_1_io_outs_right[8] ;
 wire \ces_0_1_io_outs_right[9] ;
 wire \ces_0_1_io_outs_up[0] ;
 wire \ces_0_1_io_outs_up[10] ;
 wire \ces_0_1_io_outs_up[11] ;
 wire \ces_0_1_io_outs_up[12] ;
 wire \ces_0_1_io_outs_up[13] ;
 wire \ces_0_1_io_outs_up[14] ;
 wire \ces_0_1_io_outs_up[15] ;
 wire \ces_0_1_io_outs_up[16] ;
 wire \ces_0_1_io_outs_up[17] ;
 wire \ces_0_1_io_outs_up[18] ;
 wire \ces_0_1_io_outs_up[19] ;
 wire \ces_0_1_io_outs_up[1] ;
 wire \ces_0_1_io_outs_up[20] ;
 wire \ces_0_1_io_outs_up[21] ;
 wire \ces_0_1_io_outs_up[22] ;
 wire \ces_0_1_io_outs_up[23] ;
 wire \ces_0_1_io_outs_up[24] ;
 wire \ces_0_1_io_outs_up[25] ;
 wire \ces_0_1_io_outs_up[26] ;
 wire \ces_0_1_io_outs_up[27] ;
 wire \ces_0_1_io_outs_up[28] ;
 wire \ces_0_1_io_outs_up[29] ;
 wire \ces_0_1_io_outs_up[2] ;
 wire \ces_0_1_io_outs_up[30] ;
 wire \ces_0_1_io_outs_up[31] ;
 wire \ces_0_1_io_outs_up[32] ;
 wire \ces_0_1_io_outs_up[33] ;
 wire \ces_0_1_io_outs_up[34] ;
 wire \ces_0_1_io_outs_up[35] ;
 wire \ces_0_1_io_outs_up[36] ;
 wire \ces_0_1_io_outs_up[37] ;
 wire \ces_0_1_io_outs_up[38] ;
 wire \ces_0_1_io_outs_up[39] ;
 wire \ces_0_1_io_outs_up[3] ;
 wire \ces_0_1_io_outs_up[40] ;
 wire \ces_0_1_io_outs_up[41] ;
 wire \ces_0_1_io_outs_up[42] ;
 wire \ces_0_1_io_outs_up[43] ;
 wire \ces_0_1_io_outs_up[44] ;
 wire \ces_0_1_io_outs_up[45] ;
 wire \ces_0_1_io_outs_up[46] ;
 wire \ces_0_1_io_outs_up[47] ;
 wire \ces_0_1_io_outs_up[48] ;
 wire \ces_0_1_io_outs_up[49] ;
 wire \ces_0_1_io_outs_up[4] ;
 wire \ces_0_1_io_outs_up[50] ;
 wire \ces_0_1_io_outs_up[51] ;
 wire \ces_0_1_io_outs_up[52] ;
 wire \ces_0_1_io_outs_up[53] ;
 wire \ces_0_1_io_outs_up[54] ;
 wire \ces_0_1_io_outs_up[55] ;
 wire \ces_0_1_io_outs_up[56] ;
 wire \ces_0_1_io_outs_up[57] ;
 wire \ces_0_1_io_outs_up[58] ;
 wire \ces_0_1_io_outs_up[59] ;
 wire \ces_0_1_io_outs_up[5] ;
 wire \ces_0_1_io_outs_up[60] ;
 wire \ces_0_1_io_outs_up[61] ;
 wire \ces_0_1_io_outs_up[62] ;
 wire \ces_0_1_io_outs_up[63] ;
 wire \ces_0_1_io_outs_up[6] ;
 wire \ces_0_1_io_outs_up[7] ;
 wire \ces_0_1_io_outs_up[8] ;
 wire \ces_0_1_io_outs_up[9] ;
 wire \ces_0_2_io_ins_down[0] ;
 wire \ces_0_2_io_ins_down[10] ;
 wire \ces_0_2_io_ins_down[11] ;
 wire \ces_0_2_io_ins_down[12] ;
 wire \ces_0_2_io_ins_down[13] ;
 wire \ces_0_2_io_ins_down[14] ;
 wire \ces_0_2_io_ins_down[15] ;
 wire \ces_0_2_io_ins_down[16] ;
 wire \ces_0_2_io_ins_down[17] ;
 wire \ces_0_2_io_ins_down[18] ;
 wire \ces_0_2_io_ins_down[19] ;
 wire \ces_0_2_io_ins_down[1] ;
 wire \ces_0_2_io_ins_down[20] ;
 wire \ces_0_2_io_ins_down[21] ;
 wire \ces_0_2_io_ins_down[22] ;
 wire \ces_0_2_io_ins_down[23] ;
 wire \ces_0_2_io_ins_down[24] ;
 wire \ces_0_2_io_ins_down[25] ;
 wire \ces_0_2_io_ins_down[26] ;
 wire \ces_0_2_io_ins_down[27] ;
 wire \ces_0_2_io_ins_down[28] ;
 wire \ces_0_2_io_ins_down[29] ;
 wire \ces_0_2_io_ins_down[2] ;
 wire \ces_0_2_io_ins_down[30] ;
 wire \ces_0_2_io_ins_down[31] ;
 wire \ces_0_2_io_ins_down[32] ;
 wire \ces_0_2_io_ins_down[33] ;
 wire \ces_0_2_io_ins_down[34] ;
 wire \ces_0_2_io_ins_down[35] ;
 wire \ces_0_2_io_ins_down[36] ;
 wire \ces_0_2_io_ins_down[37] ;
 wire \ces_0_2_io_ins_down[38] ;
 wire \ces_0_2_io_ins_down[39] ;
 wire \ces_0_2_io_ins_down[3] ;
 wire \ces_0_2_io_ins_down[40] ;
 wire \ces_0_2_io_ins_down[41] ;
 wire \ces_0_2_io_ins_down[42] ;
 wire \ces_0_2_io_ins_down[43] ;
 wire \ces_0_2_io_ins_down[44] ;
 wire \ces_0_2_io_ins_down[45] ;
 wire \ces_0_2_io_ins_down[46] ;
 wire \ces_0_2_io_ins_down[47] ;
 wire \ces_0_2_io_ins_down[48] ;
 wire \ces_0_2_io_ins_down[49] ;
 wire \ces_0_2_io_ins_down[4] ;
 wire \ces_0_2_io_ins_down[50] ;
 wire \ces_0_2_io_ins_down[51] ;
 wire \ces_0_2_io_ins_down[52] ;
 wire \ces_0_2_io_ins_down[53] ;
 wire \ces_0_2_io_ins_down[54] ;
 wire \ces_0_2_io_ins_down[55] ;
 wire \ces_0_2_io_ins_down[56] ;
 wire \ces_0_2_io_ins_down[57] ;
 wire \ces_0_2_io_ins_down[58] ;
 wire \ces_0_2_io_ins_down[59] ;
 wire \ces_0_2_io_ins_down[5] ;
 wire \ces_0_2_io_ins_down[60] ;
 wire \ces_0_2_io_ins_down[61] ;
 wire \ces_0_2_io_ins_down[62] ;
 wire \ces_0_2_io_ins_down[63] ;
 wire \ces_0_2_io_ins_down[6] ;
 wire \ces_0_2_io_ins_down[7] ;
 wire \ces_0_2_io_ins_down[8] ;
 wire \ces_0_2_io_ins_down[9] ;
 wire \ces_0_2_io_ins_left[0] ;
 wire \ces_0_2_io_ins_left[10] ;
 wire \ces_0_2_io_ins_left[11] ;
 wire \ces_0_2_io_ins_left[12] ;
 wire \ces_0_2_io_ins_left[13] ;
 wire \ces_0_2_io_ins_left[14] ;
 wire \ces_0_2_io_ins_left[15] ;
 wire \ces_0_2_io_ins_left[16] ;
 wire \ces_0_2_io_ins_left[17] ;
 wire \ces_0_2_io_ins_left[18] ;
 wire \ces_0_2_io_ins_left[19] ;
 wire \ces_0_2_io_ins_left[1] ;
 wire \ces_0_2_io_ins_left[20] ;
 wire \ces_0_2_io_ins_left[21] ;
 wire \ces_0_2_io_ins_left[22] ;
 wire \ces_0_2_io_ins_left[23] ;
 wire \ces_0_2_io_ins_left[24] ;
 wire \ces_0_2_io_ins_left[25] ;
 wire \ces_0_2_io_ins_left[26] ;
 wire \ces_0_2_io_ins_left[27] ;
 wire \ces_0_2_io_ins_left[28] ;
 wire \ces_0_2_io_ins_left[29] ;
 wire \ces_0_2_io_ins_left[2] ;
 wire \ces_0_2_io_ins_left[30] ;
 wire \ces_0_2_io_ins_left[31] ;
 wire \ces_0_2_io_ins_left[32] ;
 wire \ces_0_2_io_ins_left[33] ;
 wire \ces_0_2_io_ins_left[34] ;
 wire \ces_0_2_io_ins_left[35] ;
 wire \ces_0_2_io_ins_left[36] ;
 wire \ces_0_2_io_ins_left[37] ;
 wire \ces_0_2_io_ins_left[38] ;
 wire \ces_0_2_io_ins_left[39] ;
 wire \ces_0_2_io_ins_left[3] ;
 wire \ces_0_2_io_ins_left[40] ;
 wire \ces_0_2_io_ins_left[41] ;
 wire \ces_0_2_io_ins_left[42] ;
 wire \ces_0_2_io_ins_left[43] ;
 wire \ces_0_2_io_ins_left[44] ;
 wire \ces_0_2_io_ins_left[45] ;
 wire \ces_0_2_io_ins_left[46] ;
 wire \ces_0_2_io_ins_left[47] ;
 wire \ces_0_2_io_ins_left[48] ;
 wire \ces_0_2_io_ins_left[49] ;
 wire \ces_0_2_io_ins_left[4] ;
 wire \ces_0_2_io_ins_left[50] ;
 wire \ces_0_2_io_ins_left[51] ;
 wire \ces_0_2_io_ins_left[52] ;
 wire \ces_0_2_io_ins_left[53] ;
 wire \ces_0_2_io_ins_left[54] ;
 wire \ces_0_2_io_ins_left[55] ;
 wire \ces_0_2_io_ins_left[56] ;
 wire \ces_0_2_io_ins_left[57] ;
 wire \ces_0_2_io_ins_left[58] ;
 wire \ces_0_2_io_ins_left[59] ;
 wire \ces_0_2_io_ins_left[5] ;
 wire \ces_0_2_io_ins_left[60] ;
 wire \ces_0_2_io_ins_left[61] ;
 wire \ces_0_2_io_ins_left[62] ;
 wire \ces_0_2_io_ins_left[63] ;
 wire \ces_0_2_io_ins_left[6] ;
 wire \ces_0_2_io_ins_left[7] ;
 wire \ces_0_2_io_ins_left[8] ;
 wire \ces_0_2_io_ins_left[9] ;
 wire ces_0_2_io_lsbOuts_0;
 wire ces_0_2_io_lsbOuts_1;
 wire ces_0_2_io_lsbOuts_2;
 wire ces_0_2_io_lsbOuts_3;
 wire ces_0_2_io_lsbOuts_4;
 wire ces_0_2_io_lsbOuts_5;
 wire ces_0_2_io_lsbOuts_6;
 wire ces_0_2_io_lsbOuts_7;
 wire \ces_0_2_io_outs_right[0] ;
 wire \ces_0_2_io_outs_right[10] ;
 wire \ces_0_2_io_outs_right[11] ;
 wire \ces_0_2_io_outs_right[12] ;
 wire \ces_0_2_io_outs_right[13] ;
 wire \ces_0_2_io_outs_right[14] ;
 wire \ces_0_2_io_outs_right[15] ;
 wire \ces_0_2_io_outs_right[16] ;
 wire \ces_0_2_io_outs_right[17] ;
 wire \ces_0_2_io_outs_right[18] ;
 wire \ces_0_2_io_outs_right[19] ;
 wire \ces_0_2_io_outs_right[1] ;
 wire \ces_0_2_io_outs_right[20] ;
 wire \ces_0_2_io_outs_right[21] ;
 wire \ces_0_2_io_outs_right[22] ;
 wire \ces_0_2_io_outs_right[23] ;
 wire \ces_0_2_io_outs_right[24] ;
 wire \ces_0_2_io_outs_right[25] ;
 wire \ces_0_2_io_outs_right[26] ;
 wire \ces_0_2_io_outs_right[27] ;
 wire \ces_0_2_io_outs_right[28] ;
 wire \ces_0_2_io_outs_right[29] ;
 wire \ces_0_2_io_outs_right[2] ;
 wire \ces_0_2_io_outs_right[30] ;
 wire \ces_0_2_io_outs_right[31] ;
 wire \ces_0_2_io_outs_right[32] ;
 wire \ces_0_2_io_outs_right[33] ;
 wire \ces_0_2_io_outs_right[34] ;
 wire \ces_0_2_io_outs_right[35] ;
 wire \ces_0_2_io_outs_right[36] ;
 wire \ces_0_2_io_outs_right[37] ;
 wire \ces_0_2_io_outs_right[38] ;
 wire \ces_0_2_io_outs_right[39] ;
 wire \ces_0_2_io_outs_right[3] ;
 wire \ces_0_2_io_outs_right[40] ;
 wire \ces_0_2_io_outs_right[41] ;
 wire \ces_0_2_io_outs_right[42] ;
 wire \ces_0_2_io_outs_right[43] ;
 wire \ces_0_2_io_outs_right[44] ;
 wire \ces_0_2_io_outs_right[45] ;
 wire \ces_0_2_io_outs_right[46] ;
 wire \ces_0_2_io_outs_right[47] ;
 wire \ces_0_2_io_outs_right[48] ;
 wire \ces_0_2_io_outs_right[49] ;
 wire \ces_0_2_io_outs_right[4] ;
 wire \ces_0_2_io_outs_right[50] ;
 wire \ces_0_2_io_outs_right[51] ;
 wire \ces_0_2_io_outs_right[52] ;
 wire \ces_0_2_io_outs_right[53] ;
 wire \ces_0_2_io_outs_right[54] ;
 wire \ces_0_2_io_outs_right[55] ;
 wire \ces_0_2_io_outs_right[56] ;
 wire \ces_0_2_io_outs_right[57] ;
 wire \ces_0_2_io_outs_right[58] ;
 wire \ces_0_2_io_outs_right[59] ;
 wire \ces_0_2_io_outs_right[5] ;
 wire \ces_0_2_io_outs_right[60] ;
 wire \ces_0_2_io_outs_right[61] ;
 wire \ces_0_2_io_outs_right[62] ;
 wire \ces_0_2_io_outs_right[63] ;
 wire \ces_0_2_io_outs_right[6] ;
 wire \ces_0_2_io_outs_right[7] ;
 wire \ces_0_2_io_outs_right[8] ;
 wire \ces_0_2_io_outs_right[9] ;
 wire \ces_0_2_io_outs_up[0] ;
 wire \ces_0_2_io_outs_up[10] ;
 wire \ces_0_2_io_outs_up[11] ;
 wire \ces_0_2_io_outs_up[12] ;
 wire \ces_0_2_io_outs_up[13] ;
 wire \ces_0_2_io_outs_up[14] ;
 wire \ces_0_2_io_outs_up[15] ;
 wire \ces_0_2_io_outs_up[16] ;
 wire \ces_0_2_io_outs_up[17] ;
 wire \ces_0_2_io_outs_up[18] ;
 wire \ces_0_2_io_outs_up[19] ;
 wire \ces_0_2_io_outs_up[1] ;
 wire \ces_0_2_io_outs_up[20] ;
 wire \ces_0_2_io_outs_up[21] ;
 wire \ces_0_2_io_outs_up[22] ;
 wire \ces_0_2_io_outs_up[23] ;
 wire \ces_0_2_io_outs_up[24] ;
 wire \ces_0_2_io_outs_up[25] ;
 wire \ces_0_2_io_outs_up[26] ;
 wire \ces_0_2_io_outs_up[27] ;
 wire \ces_0_2_io_outs_up[28] ;
 wire \ces_0_2_io_outs_up[29] ;
 wire \ces_0_2_io_outs_up[2] ;
 wire \ces_0_2_io_outs_up[30] ;
 wire \ces_0_2_io_outs_up[31] ;
 wire \ces_0_2_io_outs_up[32] ;
 wire \ces_0_2_io_outs_up[33] ;
 wire \ces_0_2_io_outs_up[34] ;
 wire \ces_0_2_io_outs_up[35] ;
 wire \ces_0_2_io_outs_up[36] ;
 wire \ces_0_2_io_outs_up[37] ;
 wire \ces_0_2_io_outs_up[38] ;
 wire \ces_0_2_io_outs_up[39] ;
 wire \ces_0_2_io_outs_up[3] ;
 wire \ces_0_2_io_outs_up[40] ;
 wire \ces_0_2_io_outs_up[41] ;
 wire \ces_0_2_io_outs_up[42] ;
 wire \ces_0_2_io_outs_up[43] ;
 wire \ces_0_2_io_outs_up[44] ;
 wire \ces_0_2_io_outs_up[45] ;
 wire \ces_0_2_io_outs_up[46] ;
 wire \ces_0_2_io_outs_up[47] ;
 wire \ces_0_2_io_outs_up[48] ;
 wire \ces_0_2_io_outs_up[49] ;
 wire \ces_0_2_io_outs_up[4] ;
 wire \ces_0_2_io_outs_up[50] ;
 wire \ces_0_2_io_outs_up[51] ;
 wire \ces_0_2_io_outs_up[52] ;
 wire \ces_0_2_io_outs_up[53] ;
 wire \ces_0_2_io_outs_up[54] ;
 wire \ces_0_2_io_outs_up[55] ;
 wire \ces_0_2_io_outs_up[56] ;
 wire \ces_0_2_io_outs_up[57] ;
 wire \ces_0_2_io_outs_up[58] ;
 wire \ces_0_2_io_outs_up[59] ;
 wire \ces_0_2_io_outs_up[5] ;
 wire \ces_0_2_io_outs_up[60] ;
 wire \ces_0_2_io_outs_up[61] ;
 wire \ces_0_2_io_outs_up[62] ;
 wire \ces_0_2_io_outs_up[63] ;
 wire \ces_0_2_io_outs_up[6] ;
 wire \ces_0_2_io_outs_up[7] ;
 wire \ces_0_2_io_outs_up[8] ;
 wire \ces_0_2_io_outs_up[9] ;
 wire \ces_0_3_io_ins_down[0] ;
 wire \ces_0_3_io_ins_down[10] ;
 wire \ces_0_3_io_ins_down[11] ;
 wire \ces_0_3_io_ins_down[12] ;
 wire \ces_0_3_io_ins_down[13] ;
 wire \ces_0_3_io_ins_down[14] ;
 wire \ces_0_3_io_ins_down[15] ;
 wire \ces_0_3_io_ins_down[16] ;
 wire \ces_0_3_io_ins_down[17] ;
 wire \ces_0_3_io_ins_down[18] ;
 wire \ces_0_3_io_ins_down[19] ;
 wire \ces_0_3_io_ins_down[1] ;
 wire \ces_0_3_io_ins_down[20] ;
 wire \ces_0_3_io_ins_down[21] ;
 wire \ces_0_3_io_ins_down[22] ;
 wire \ces_0_3_io_ins_down[23] ;
 wire \ces_0_3_io_ins_down[24] ;
 wire \ces_0_3_io_ins_down[25] ;
 wire \ces_0_3_io_ins_down[26] ;
 wire \ces_0_3_io_ins_down[27] ;
 wire \ces_0_3_io_ins_down[28] ;
 wire \ces_0_3_io_ins_down[29] ;
 wire \ces_0_3_io_ins_down[2] ;
 wire \ces_0_3_io_ins_down[30] ;
 wire \ces_0_3_io_ins_down[31] ;
 wire \ces_0_3_io_ins_down[32] ;
 wire \ces_0_3_io_ins_down[33] ;
 wire \ces_0_3_io_ins_down[34] ;
 wire \ces_0_3_io_ins_down[35] ;
 wire \ces_0_3_io_ins_down[36] ;
 wire \ces_0_3_io_ins_down[37] ;
 wire \ces_0_3_io_ins_down[38] ;
 wire \ces_0_3_io_ins_down[39] ;
 wire \ces_0_3_io_ins_down[3] ;
 wire \ces_0_3_io_ins_down[40] ;
 wire \ces_0_3_io_ins_down[41] ;
 wire \ces_0_3_io_ins_down[42] ;
 wire \ces_0_3_io_ins_down[43] ;
 wire \ces_0_3_io_ins_down[44] ;
 wire \ces_0_3_io_ins_down[45] ;
 wire \ces_0_3_io_ins_down[46] ;
 wire \ces_0_3_io_ins_down[47] ;
 wire \ces_0_3_io_ins_down[48] ;
 wire \ces_0_3_io_ins_down[49] ;
 wire \ces_0_3_io_ins_down[4] ;
 wire \ces_0_3_io_ins_down[50] ;
 wire \ces_0_3_io_ins_down[51] ;
 wire \ces_0_3_io_ins_down[52] ;
 wire \ces_0_3_io_ins_down[53] ;
 wire \ces_0_3_io_ins_down[54] ;
 wire \ces_0_3_io_ins_down[55] ;
 wire \ces_0_3_io_ins_down[56] ;
 wire \ces_0_3_io_ins_down[57] ;
 wire \ces_0_3_io_ins_down[58] ;
 wire \ces_0_3_io_ins_down[59] ;
 wire \ces_0_3_io_ins_down[5] ;
 wire \ces_0_3_io_ins_down[60] ;
 wire \ces_0_3_io_ins_down[61] ;
 wire \ces_0_3_io_ins_down[62] ;
 wire \ces_0_3_io_ins_down[63] ;
 wire \ces_0_3_io_ins_down[6] ;
 wire \ces_0_3_io_ins_down[7] ;
 wire \ces_0_3_io_ins_down[8] ;
 wire \ces_0_3_io_ins_down[9] ;
 wire \ces_0_3_io_ins_left[0] ;
 wire \ces_0_3_io_ins_left[10] ;
 wire \ces_0_3_io_ins_left[11] ;
 wire \ces_0_3_io_ins_left[12] ;
 wire \ces_0_3_io_ins_left[13] ;
 wire \ces_0_3_io_ins_left[14] ;
 wire \ces_0_3_io_ins_left[15] ;
 wire \ces_0_3_io_ins_left[16] ;
 wire \ces_0_3_io_ins_left[17] ;
 wire \ces_0_3_io_ins_left[18] ;
 wire \ces_0_3_io_ins_left[19] ;
 wire \ces_0_3_io_ins_left[1] ;
 wire \ces_0_3_io_ins_left[20] ;
 wire \ces_0_3_io_ins_left[21] ;
 wire \ces_0_3_io_ins_left[22] ;
 wire \ces_0_3_io_ins_left[23] ;
 wire \ces_0_3_io_ins_left[24] ;
 wire \ces_0_3_io_ins_left[25] ;
 wire \ces_0_3_io_ins_left[26] ;
 wire \ces_0_3_io_ins_left[27] ;
 wire \ces_0_3_io_ins_left[28] ;
 wire \ces_0_3_io_ins_left[29] ;
 wire \ces_0_3_io_ins_left[2] ;
 wire \ces_0_3_io_ins_left[30] ;
 wire \ces_0_3_io_ins_left[31] ;
 wire \ces_0_3_io_ins_left[32] ;
 wire \ces_0_3_io_ins_left[33] ;
 wire \ces_0_3_io_ins_left[34] ;
 wire \ces_0_3_io_ins_left[35] ;
 wire \ces_0_3_io_ins_left[36] ;
 wire \ces_0_3_io_ins_left[37] ;
 wire \ces_0_3_io_ins_left[38] ;
 wire \ces_0_3_io_ins_left[39] ;
 wire \ces_0_3_io_ins_left[3] ;
 wire \ces_0_3_io_ins_left[40] ;
 wire \ces_0_3_io_ins_left[41] ;
 wire \ces_0_3_io_ins_left[42] ;
 wire \ces_0_3_io_ins_left[43] ;
 wire \ces_0_3_io_ins_left[44] ;
 wire \ces_0_3_io_ins_left[45] ;
 wire \ces_0_3_io_ins_left[46] ;
 wire \ces_0_3_io_ins_left[47] ;
 wire \ces_0_3_io_ins_left[48] ;
 wire \ces_0_3_io_ins_left[49] ;
 wire \ces_0_3_io_ins_left[4] ;
 wire \ces_0_3_io_ins_left[50] ;
 wire \ces_0_3_io_ins_left[51] ;
 wire \ces_0_3_io_ins_left[52] ;
 wire \ces_0_3_io_ins_left[53] ;
 wire \ces_0_3_io_ins_left[54] ;
 wire \ces_0_3_io_ins_left[55] ;
 wire \ces_0_3_io_ins_left[56] ;
 wire \ces_0_3_io_ins_left[57] ;
 wire \ces_0_3_io_ins_left[58] ;
 wire \ces_0_3_io_ins_left[59] ;
 wire \ces_0_3_io_ins_left[5] ;
 wire \ces_0_3_io_ins_left[60] ;
 wire \ces_0_3_io_ins_left[61] ;
 wire \ces_0_3_io_ins_left[62] ;
 wire \ces_0_3_io_ins_left[63] ;
 wire \ces_0_3_io_ins_left[6] ;
 wire \ces_0_3_io_ins_left[7] ;
 wire \ces_0_3_io_ins_left[8] ;
 wire \ces_0_3_io_ins_left[9] ;
 wire ces_0_3_io_lsbOuts_0;
 wire ces_0_3_io_lsbOuts_1;
 wire ces_0_3_io_lsbOuts_2;
 wire ces_0_3_io_lsbOuts_3;
 wire ces_0_3_io_lsbOuts_4;
 wire ces_0_3_io_lsbOuts_5;
 wire ces_0_3_io_lsbOuts_6;
 wire ces_0_3_io_lsbOuts_7;
 wire \ces_0_3_io_outs_right[0] ;
 wire \ces_0_3_io_outs_right[10] ;
 wire \ces_0_3_io_outs_right[11] ;
 wire \ces_0_3_io_outs_right[12] ;
 wire \ces_0_3_io_outs_right[13] ;
 wire \ces_0_3_io_outs_right[14] ;
 wire \ces_0_3_io_outs_right[15] ;
 wire \ces_0_3_io_outs_right[16] ;
 wire \ces_0_3_io_outs_right[17] ;
 wire \ces_0_3_io_outs_right[18] ;
 wire \ces_0_3_io_outs_right[19] ;
 wire \ces_0_3_io_outs_right[1] ;
 wire \ces_0_3_io_outs_right[20] ;
 wire \ces_0_3_io_outs_right[21] ;
 wire \ces_0_3_io_outs_right[22] ;
 wire \ces_0_3_io_outs_right[23] ;
 wire \ces_0_3_io_outs_right[24] ;
 wire \ces_0_3_io_outs_right[25] ;
 wire \ces_0_3_io_outs_right[26] ;
 wire \ces_0_3_io_outs_right[27] ;
 wire \ces_0_3_io_outs_right[28] ;
 wire \ces_0_3_io_outs_right[29] ;
 wire \ces_0_3_io_outs_right[2] ;
 wire \ces_0_3_io_outs_right[30] ;
 wire \ces_0_3_io_outs_right[31] ;
 wire \ces_0_3_io_outs_right[32] ;
 wire \ces_0_3_io_outs_right[33] ;
 wire \ces_0_3_io_outs_right[34] ;
 wire \ces_0_3_io_outs_right[35] ;
 wire \ces_0_3_io_outs_right[36] ;
 wire \ces_0_3_io_outs_right[37] ;
 wire \ces_0_3_io_outs_right[38] ;
 wire \ces_0_3_io_outs_right[39] ;
 wire \ces_0_3_io_outs_right[3] ;
 wire \ces_0_3_io_outs_right[40] ;
 wire \ces_0_3_io_outs_right[41] ;
 wire \ces_0_3_io_outs_right[42] ;
 wire \ces_0_3_io_outs_right[43] ;
 wire \ces_0_3_io_outs_right[44] ;
 wire \ces_0_3_io_outs_right[45] ;
 wire \ces_0_3_io_outs_right[46] ;
 wire \ces_0_3_io_outs_right[47] ;
 wire \ces_0_3_io_outs_right[48] ;
 wire \ces_0_3_io_outs_right[49] ;
 wire \ces_0_3_io_outs_right[4] ;
 wire \ces_0_3_io_outs_right[50] ;
 wire \ces_0_3_io_outs_right[51] ;
 wire \ces_0_3_io_outs_right[52] ;
 wire \ces_0_3_io_outs_right[53] ;
 wire \ces_0_3_io_outs_right[54] ;
 wire \ces_0_3_io_outs_right[55] ;
 wire \ces_0_3_io_outs_right[56] ;
 wire \ces_0_3_io_outs_right[57] ;
 wire \ces_0_3_io_outs_right[58] ;
 wire \ces_0_3_io_outs_right[59] ;
 wire \ces_0_3_io_outs_right[5] ;
 wire \ces_0_3_io_outs_right[60] ;
 wire \ces_0_3_io_outs_right[61] ;
 wire \ces_0_3_io_outs_right[62] ;
 wire \ces_0_3_io_outs_right[63] ;
 wire \ces_0_3_io_outs_right[6] ;
 wire \ces_0_3_io_outs_right[7] ;
 wire \ces_0_3_io_outs_right[8] ;
 wire \ces_0_3_io_outs_right[9] ;
 wire \ces_0_3_io_outs_up[0] ;
 wire \ces_0_3_io_outs_up[10] ;
 wire \ces_0_3_io_outs_up[11] ;
 wire \ces_0_3_io_outs_up[12] ;
 wire \ces_0_3_io_outs_up[13] ;
 wire \ces_0_3_io_outs_up[14] ;
 wire \ces_0_3_io_outs_up[15] ;
 wire \ces_0_3_io_outs_up[16] ;
 wire \ces_0_3_io_outs_up[17] ;
 wire \ces_0_3_io_outs_up[18] ;
 wire \ces_0_3_io_outs_up[19] ;
 wire \ces_0_3_io_outs_up[1] ;
 wire \ces_0_3_io_outs_up[20] ;
 wire \ces_0_3_io_outs_up[21] ;
 wire \ces_0_3_io_outs_up[22] ;
 wire \ces_0_3_io_outs_up[23] ;
 wire \ces_0_3_io_outs_up[24] ;
 wire \ces_0_3_io_outs_up[25] ;
 wire \ces_0_3_io_outs_up[26] ;
 wire \ces_0_3_io_outs_up[27] ;
 wire \ces_0_3_io_outs_up[28] ;
 wire \ces_0_3_io_outs_up[29] ;
 wire \ces_0_3_io_outs_up[2] ;
 wire \ces_0_3_io_outs_up[30] ;
 wire \ces_0_3_io_outs_up[31] ;
 wire \ces_0_3_io_outs_up[32] ;
 wire \ces_0_3_io_outs_up[33] ;
 wire \ces_0_3_io_outs_up[34] ;
 wire \ces_0_3_io_outs_up[35] ;
 wire \ces_0_3_io_outs_up[36] ;
 wire \ces_0_3_io_outs_up[37] ;
 wire \ces_0_3_io_outs_up[38] ;
 wire \ces_0_3_io_outs_up[39] ;
 wire \ces_0_3_io_outs_up[3] ;
 wire \ces_0_3_io_outs_up[40] ;
 wire \ces_0_3_io_outs_up[41] ;
 wire \ces_0_3_io_outs_up[42] ;
 wire \ces_0_3_io_outs_up[43] ;
 wire \ces_0_3_io_outs_up[44] ;
 wire \ces_0_3_io_outs_up[45] ;
 wire \ces_0_3_io_outs_up[46] ;
 wire \ces_0_3_io_outs_up[47] ;
 wire \ces_0_3_io_outs_up[48] ;
 wire \ces_0_3_io_outs_up[49] ;
 wire \ces_0_3_io_outs_up[4] ;
 wire \ces_0_3_io_outs_up[50] ;
 wire \ces_0_3_io_outs_up[51] ;
 wire \ces_0_3_io_outs_up[52] ;
 wire \ces_0_3_io_outs_up[53] ;
 wire \ces_0_3_io_outs_up[54] ;
 wire \ces_0_3_io_outs_up[55] ;
 wire \ces_0_3_io_outs_up[56] ;
 wire \ces_0_3_io_outs_up[57] ;
 wire \ces_0_3_io_outs_up[58] ;
 wire \ces_0_3_io_outs_up[59] ;
 wire \ces_0_3_io_outs_up[5] ;
 wire \ces_0_3_io_outs_up[60] ;
 wire \ces_0_3_io_outs_up[61] ;
 wire \ces_0_3_io_outs_up[62] ;
 wire \ces_0_3_io_outs_up[63] ;
 wire \ces_0_3_io_outs_up[6] ;
 wire \ces_0_3_io_outs_up[7] ;
 wire \ces_0_3_io_outs_up[8] ;
 wire \ces_0_3_io_outs_up[9] ;
 wire \ces_0_4_io_ins_down[0] ;
 wire \ces_0_4_io_ins_down[10] ;
 wire \ces_0_4_io_ins_down[11] ;
 wire \ces_0_4_io_ins_down[12] ;
 wire \ces_0_4_io_ins_down[13] ;
 wire \ces_0_4_io_ins_down[14] ;
 wire \ces_0_4_io_ins_down[15] ;
 wire \ces_0_4_io_ins_down[16] ;
 wire \ces_0_4_io_ins_down[17] ;
 wire \ces_0_4_io_ins_down[18] ;
 wire \ces_0_4_io_ins_down[19] ;
 wire \ces_0_4_io_ins_down[1] ;
 wire \ces_0_4_io_ins_down[20] ;
 wire \ces_0_4_io_ins_down[21] ;
 wire \ces_0_4_io_ins_down[22] ;
 wire \ces_0_4_io_ins_down[23] ;
 wire \ces_0_4_io_ins_down[24] ;
 wire \ces_0_4_io_ins_down[25] ;
 wire \ces_0_4_io_ins_down[26] ;
 wire \ces_0_4_io_ins_down[27] ;
 wire \ces_0_4_io_ins_down[28] ;
 wire \ces_0_4_io_ins_down[29] ;
 wire \ces_0_4_io_ins_down[2] ;
 wire \ces_0_4_io_ins_down[30] ;
 wire \ces_0_4_io_ins_down[31] ;
 wire \ces_0_4_io_ins_down[32] ;
 wire \ces_0_4_io_ins_down[33] ;
 wire \ces_0_4_io_ins_down[34] ;
 wire \ces_0_4_io_ins_down[35] ;
 wire \ces_0_4_io_ins_down[36] ;
 wire \ces_0_4_io_ins_down[37] ;
 wire \ces_0_4_io_ins_down[38] ;
 wire \ces_0_4_io_ins_down[39] ;
 wire \ces_0_4_io_ins_down[3] ;
 wire \ces_0_4_io_ins_down[40] ;
 wire \ces_0_4_io_ins_down[41] ;
 wire \ces_0_4_io_ins_down[42] ;
 wire \ces_0_4_io_ins_down[43] ;
 wire \ces_0_4_io_ins_down[44] ;
 wire \ces_0_4_io_ins_down[45] ;
 wire \ces_0_4_io_ins_down[46] ;
 wire \ces_0_4_io_ins_down[47] ;
 wire \ces_0_4_io_ins_down[48] ;
 wire \ces_0_4_io_ins_down[49] ;
 wire \ces_0_4_io_ins_down[4] ;
 wire \ces_0_4_io_ins_down[50] ;
 wire \ces_0_4_io_ins_down[51] ;
 wire \ces_0_4_io_ins_down[52] ;
 wire \ces_0_4_io_ins_down[53] ;
 wire \ces_0_4_io_ins_down[54] ;
 wire \ces_0_4_io_ins_down[55] ;
 wire \ces_0_4_io_ins_down[56] ;
 wire \ces_0_4_io_ins_down[57] ;
 wire \ces_0_4_io_ins_down[58] ;
 wire \ces_0_4_io_ins_down[59] ;
 wire \ces_0_4_io_ins_down[5] ;
 wire \ces_0_4_io_ins_down[60] ;
 wire \ces_0_4_io_ins_down[61] ;
 wire \ces_0_4_io_ins_down[62] ;
 wire \ces_0_4_io_ins_down[63] ;
 wire \ces_0_4_io_ins_down[6] ;
 wire \ces_0_4_io_ins_down[7] ;
 wire \ces_0_4_io_ins_down[8] ;
 wire \ces_0_4_io_ins_down[9] ;
 wire \ces_0_4_io_ins_left[0] ;
 wire \ces_0_4_io_ins_left[10] ;
 wire \ces_0_4_io_ins_left[11] ;
 wire \ces_0_4_io_ins_left[12] ;
 wire \ces_0_4_io_ins_left[13] ;
 wire \ces_0_4_io_ins_left[14] ;
 wire \ces_0_4_io_ins_left[15] ;
 wire \ces_0_4_io_ins_left[16] ;
 wire \ces_0_4_io_ins_left[17] ;
 wire \ces_0_4_io_ins_left[18] ;
 wire \ces_0_4_io_ins_left[19] ;
 wire \ces_0_4_io_ins_left[1] ;
 wire \ces_0_4_io_ins_left[20] ;
 wire \ces_0_4_io_ins_left[21] ;
 wire \ces_0_4_io_ins_left[22] ;
 wire \ces_0_4_io_ins_left[23] ;
 wire \ces_0_4_io_ins_left[24] ;
 wire \ces_0_4_io_ins_left[25] ;
 wire \ces_0_4_io_ins_left[26] ;
 wire \ces_0_4_io_ins_left[27] ;
 wire \ces_0_4_io_ins_left[28] ;
 wire \ces_0_4_io_ins_left[29] ;
 wire \ces_0_4_io_ins_left[2] ;
 wire \ces_0_4_io_ins_left[30] ;
 wire \ces_0_4_io_ins_left[31] ;
 wire \ces_0_4_io_ins_left[32] ;
 wire \ces_0_4_io_ins_left[33] ;
 wire \ces_0_4_io_ins_left[34] ;
 wire \ces_0_4_io_ins_left[35] ;
 wire \ces_0_4_io_ins_left[36] ;
 wire \ces_0_4_io_ins_left[37] ;
 wire \ces_0_4_io_ins_left[38] ;
 wire \ces_0_4_io_ins_left[39] ;
 wire \ces_0_4_io_ins_left[3] ;
 wire \ces_0_4_io_ins_left[40] ;
 wire \ces_0_4_io_ins_left[41] ;
 wire \ces_0_4_io_ins_left[42] ;
 wire \ces_0_4_io_ins_left[43] ;
 wire \ces_0_4_io_ins_left[44] ;
 wire \ces_0_4_io_ins_left[45] ;
 wire \ces_0_4_io_ins_left[46] ;
 wire \ces_0_4_io_ins_left[47] ;
 wire \ces_0_4_io_ins_left[48] ;
 wire \ces_0_4_io_ins_left[49] ;
 wire \ces_0_4_io_ins_left[4] ;
 wire \ces_0_4_io_ins_left[50] ;
 wire \ces_0_4_io_ins_left[51] ;
 wire \ces_0_4_io_ins_left[52] ;
 wire \ces_0_4_io_ins_left[53] ;
 wire \ces_0_4_io_ins_left[54] ;
 wire \ces_0_4_io_ins_left[55] ;
 wire \ces_0_4_io_ins_left[56] ;
 wire \ces_0_4_io_ins_left[57] ;
 wire \ces_0_4_io_ins_left[58] ;
 wire \ces_0_4_io_ins_left[59] ;
 wire \ces_0_4_io_ins_left[5] ;
 wire \ces_0_4_io_ins_left[60] ;
 wire \ces_0_4_io_ins_left[61] ;
 wire \ces_0_4_io_ins_left[62] ;
 wire \ces_0_4_io_ins_left[63] ;
 wire \ces_0_4_io_ins_left[6] ;
 wire \ces_0_4_io_ins_left[7] ;
 wire \ces_0_4_io_ins_left[8] ;
 wire \ces_0_4_io_ins_left[9] ;
 wire ces_0_4_io_lsbOuts_0;
 wire ces_0_4_io_lsbOuts_1;
 wire ces_0_4_io_lsbOuts_2;
 wire ces_0_4_io_lsbOuts_3;
 wire ces_0_4_io_lsbOuts_4;
 wire ces_0_4_io_lsbOuts_5;
 wire ces_0_4_io_lsbOuts_6;
 wire ces_0_4_io_lsbOuts_7;
 wire \ces_0_4_io_outs_right[0] ;
 wire \ces_0_4_io_outs_right[10] ;
 wire \ces_0_4_io_outs_right[11] ;
 wire \ces_0_4_io_outs_right[12] ;
 wire \ces_0_4_io_outs_right[13] ;
 wire \ces_0_4_io_outs_right[14] ;
 wire \ces_0_4_io_outs_right[15] ;
 wire \ces_0_4_io_outs_right[16] ;
 wire \ces_0_4_io_outs_right[17] ;
 wire \ces_0_4_io_outs_right[18] ;
 wire \ces_0_4_io_outs_right[19] ;
 wire \ces_0_4_io_outs_right[1] ;
 wire \ces_0_4_io_outs_right[20] ;
 wire \ces_0_4_io_outs_right[21] ;
 wire \ces_0_4_io_outs_right[22] ;
 wire \ces_0_4_io_outs_right[23] ;
 wire \ces_0_4_io_outs_right[24] ;
 wire \ces_0_4_io_outs_right[25] ;
 wire \ces_0_4_io_outs_right[26] ;
 wire \ces_0_4_io_outs_right[27] ;
 wire \ces_0_4_io_outs_right[28] ;
 wire \ces_0_4_io_outs_right[29] ;
 wire \ces_0_4_io_outs_right[2] ;
 wire \ces_0_4_io_outs_right[30] ;
 wire \ces_0_4_io_outs_right[31] ;
 wire \ces_0_4_io_outs_right[32] ;
 wire \ces_0_4_io_outs_right[33] ;
 wire \ces_0_4_io_outs_right[34] ;
 wire \ces_0_4_io_outs_right[35] ;
 wire \ces_0_4_io_outs_right[36] ;
 wire \ces_0_4_io_outs_right[37] ;
 wire \ces_0_4_io_outs_right[38] ;
 wire \ces_0_4_io_outs_right[39] ;
 wire \ces_0_4_io_outs_right[3] ;
 wire \ces_0_4_io_outs_right[40] ;
 wire \ces_0_4_io_outs_right[41] ;
 wire \ces_0_4_io_outs_right[42] ;
 wire \ces_0_4_io_outs_right[43] ;
 wire \ces_0_4_io_outs_right[44] ;
 wire \ces_0_4_io_outs_right[45] ;
 wire \ces_0_4_io_outs_right[46] ;
 wire \ces_0_4_io_outs_right[47] ;
 wire \ces_0_4_io_outs_right[48] ;
 wire \ces_0_4_io_outs_right[49] ;
 wire \ces_0_4_io_outs_right[4] ;
 wire \ces_0_4_io_outs_right[50] ;
 wire \ces_0_4_io_outs_right[51] ;
 wire \ces_0_4_io_outs_right[52] ;
 wire \ces_0_4_io_outs_right[53] ;
 wire \ces_0_4_io_outs_right[54] ;
 wire \ces_0_4_io_outs_right[55] ;
 wire \ces_0_4_io_outs_right[56] ;
 wire \ces_0_4_io_outs_right[57] ;
 wire \ces_0_4_io_outs_right[58] ;
 wire \ces_0_4_io_outs_right[59] ;
 wire \ces_0_4_io_outs_right[5] ;
 wire \ces_0_4_io_outs_right[60] ;
 wire \ces_0_4_io_outs_right[61] ;
 wire \ces_0_4_io_outs_right[62] ;
 wire \ces_0_4_io_outs_right[63] ;
 wire \ces_0_4_io_outs_right[6] ;
 wire \ces_0_4_io_outs_right[7] ;
 wire \ces_0_4_io_outs_right[8] ;
 wire \ces_0_4_io_outs_right[9] ;
 wire \ces_0_4_io_outs_up[0] ;
 wire \ces_0_4_io_outs_up[10] ;
 wire \ces_0_4_io_outs_up[11] ;
 wire \ces_0_4_io_outs_up[12] ;
 wire \ces_0_4_io_outs_up[13] ;
 wire \ces_0_4_io_outs_up[14] ;
 wire \ces_0_4_io_outs_up[15] ;
 wire \ces_0_4_io_outs_up[16] ;
 wire \ces_0_4_io_outs_up[17] ;
 wire \ces_0_4_io_outs_up[18] ;
 wire \ces_0_4_io_outs_up[19] ;
 wire \ces_0_4_io_outs_up[1] ;
 wire \ces_0_4_io_outs_up[20] ;
 wire \ces_0_4_io_outs_up[21] ;
 wire \ces_0_4_io_outs_up[22] ;
 wire \ces_0_4_io_outs_up[23] ;
 wire \ces_0_4_io_outs_up[24] ;
 wire \ces_0_4_io_outs_up[25] ;
 wire \ces_0_4_io_outs_up[26] ;
 wire \ces_0_4_io_outs_up[27] ;
 wire \ces_0_4_io_outs_up[28] ;
 wire \ces_0_4_io_outs_up[29] ;
 wire \ces_0_4_io_outs_up[2] ;
 wire \ces_0_4_io_outs_up[30] ;
 wire \ces_0_4_io_outs_up[31] ;
 wire \ces_0_4_io_outs_up[32] ;
 wire \ces_0_4_io_outs_up[33] ;
 wire \ces_0_4_io_outs_up[34] ;
 wire \ces_0_4_io_outs_up[35] ;
 wire \ces_0_4_io_outs_up[36] ;
 wire \ces_0_4_io_outs_up[37] ;
 wire \ces_0_4_io_outs_up[38] ;
 wire \ces_0_4_io_outs_up[39] ;
 wire \ces_0_4_io_outs_up[3] ;
 wire \ces_0_4_io_outs_up[40] ;
 wire \ces_0_4_io_outs_up[41] ;
 wire \ces_0_4_io_outs_up[42] ;
 wire \ces_0_4_io_outs_up[43] ;
 wire \ces_0_4_io_outs_up[44] ;
 wire \ces_0_4_io_outs_up[45] ;
 wire \ces_0_4_io_outs_up[46] ;
 wire \ces_0_4_io_outs_up[47] ;
 wire \ces_0_4_io_outs_up[48] ;
 wire \ces_0_4_io_outs_up[49] ;
 wire \ces_0_4_io_outs_up[4] ;
 wire \ces_0_4_io_outs_up[50] ;
 wire \ces_0_4_io_outs_up[51] ;
 wire \ces_0_4_io_outs_up[52] ;
 wire \ces_0_4_io_outs_up[53] ;
 wire \ces_0_4_io_outs_up[54] ;
 wire \ces_0_4_io_outs_up[55] ;
 wire \ces_0_4_io_outs_up[56] ;
 wire \ces_0_4_io_outs_up[57] ;
 wire \ces_0_4_io_outs_up[58] ;
 wire \ces_0_4_io_outs_up[59] ;
 wire \ces_0_4_io_outs_up[5] ;
 wire \ces_0_4_io_outs_up[60] ;
 wire \ces_0_4_io_outs_up[61] ;
 wire \ces_0_4_io_outs_up[62] ;
 wire \ces_0_4_io_outs_up[63] ;
 wire \ces_0_4_io_outs_up[6] ;
 wire \ces_0_4_io_outs_up[7] ;
 wire \ces_0_4_io_outs_up[8] ;
 wire \ces_0_4_io_outs_up[9] ;
 wire \ces_0_5_io_ins_down[0] ;
 wire \ces_0_5_io_ins_down[10] ;
 wire \ces_0_5_io_ins_down[11] ;
 wire \ces_0_5_io_ins_down[12] ;
 wire \ces_0_5_io_ins_down[13] ;
 wire \ces_0_5_io_ins_down[14] ;
 wire \ces_0_5_io_ins_down[15] ;
 wire \ces_0_5_io_ins_down[16] ;
 wire \ces_0_5_io_ins_down[17] ;
 wire \ces_0_5_io_ins_down[18] ;
 wire \ces_0_5_io_ins_down[19] ;
 wire \ces_0_5_io_ins_down[1] ;
 wire \ces_0_5_io_ins_down[20] ;
 wire \ces_0_5_io_ins_down[21] ;
 wire \ces_0_5_io_ins_down[22] ;
 wire \ces_0_5_io_ins_down[23] ;
 wire \ces_0_5_io_ins_down[24] ;
 wire \ces_0_5_io_ins_down[25] ;
 wire \ces_0_5_io_ins_down[26] ;
 wire \ces_0_5_io_ins_down[27] ;
 wire \ces_0_5_io_ins_down[28] ;
 wire \ces_0_5_io_ins_down[29] ;
 wire \ces_0_5_io_ins_down[2] ;
 wire \ces_0_5_io_ins_down[30] ;
 wire \ces_0_5_io_ins_down[31] ;
 wire \ces_0_5_io_ins_down[32] ;
 wire \ces_0_5_io_ins_down[33] ;
 wire \ces_0_5_io_ins_down[34] ;
 wire \ces_0_5_io_ins_down[35] ;
 wire \ces_0_5_io_ins_down[36] ;
 wire \ces_0_5_io_ins_down[37] ;
 wire \ces_0_5_io_ins_down[38] ;
 wire \ces_0_5_io_ins_down[39] ;
 wire \ces_0_5_io_ins_down[3] ;
 wire \ces_0_5_io_ins_down[40] ;
 wire \ces_0_5_io_ins_down[41] ;
 wire \ces_0_5_io_ins_down[42] ;
 wire \ces_0_5_io_ins_down[43] ;
 wire \ces_0_5_io_ins_down[44] ;
 wire \ces_0_5_io_ins_down[45] ;
 wire \ces_0_5_io_ins_down[46] ;
 wire \ces_0_5_io_ins_down[47] ;
 wire \ces_0_5_io_ins_down[48] ;
 wire \ces_0_5_io_ins_down[49] ;
 wire \ces_0_5_io_ins_down[4] ;
 wire \ces_0_5_io_ins_down[50] ;
 wire \ces_0_5_io_ins_down[51] ;
 wire \ces_0_5_io_ins_down[52] ;
 wire \ces_0_5_io_ins_down[53] ;
 wire \ces_0_5_io_ins_down[54] ;
 wire \ces_0_5_io_ins_down[55] ;
 wire \ces_0_5_io_ins_down[56] ;
 wire \ces_0_5_io_ins_down[57] ;
 wire \ces_0_5_io_ins_down[58] ;
 wire \ces_0_5_io_ins_down[59] ;
 wire \ces_0_5_io_ins_down[5] ;
 wire \ces_0_5_io_ins_down[60] ;
 wire \ces_0_5_io_ins_down[61] ;
 wire \ces_0_5_io_ins_down[62] ;
 wire \ces_0_5_io_ins_down[63] ;
 wire \ces_0_5_io_ins_down[6] ;
 wire \ces_0_5_io_ins_down[7] ;
 wire \ces_0_5_io_ins_down[8] ;
 wire \ces_0_5_io_ins_down[9] ;
 wire \ces_0_5_io_ins_left[0] ;
 wire \ces_0_5_io_ins_left[10] ;
 wire \ces_0_5_io_ins_left[11] ;
 wire \ces_0_5_io_ins_left[12] ;
 wire \ces_0_5_io_ins_left[13] ;
 wire \ces_0_5_io_ins_left[14] ;
 wire \ces_0_5_io_ins_left[15] ;
 wire \ces_0_5_io_ins_left[16] ;
 wire \ces_0_5_io_ins_left[17] ;
 wire \ces_0_5_io_ins_left[18] ;
 wire \ces_0_5_io_ins_left[19] ;
 wire \ces_0_5_io_ins_left[1] ;
 wire \ces_0_5_io_ins_left[20] ;
 wire \ces_0_5_io_ins_left[21] ;
 wire \ces_0_5_io_ins_left[22] ;
 wire \ces_0_5_io_ins_left[23] ;
 wire \ces_0_5_io_ins_left[24] ;
 wire \ces_0_5_io_ins_left[25] ;
 wire \ces_0_5_io_ins_left[26] ;
 wire \ces_0_5_io_ins_left[27] ;
 wire \ces_0_5_io_ins_left[28] ;
 wire \ces_0_5_io_ins_left[29] ;
 wire \ces_0_5_io_ins_left[2] ;
 wire \ces_0_5_io_ins_left[30] ;
 wire \ces_0_5_io_ins_left[31] ;
 wire \ces_0_5_io_ins_left[32] ;
 wire \ces_0_5_io_ins_left[33] ;
 wire \ces_0_5_io_ins_left[34] ;
 wire \ces_0_5_io_ins_left[35] ;
 wire \ces_0_5_io_ins_left[36] ;
 wire \ces_0_5_io_ins_left[37] ;
 wire \ces_0_5_io_ins_left[38] ;
 wire \ces_0_5_io_ins_left[39] ;
 wire \ces_0_5_io_ins_left[3] ;
 wire \ces_0_5_io_ins_left[40] ;
 wire \ces_0_5_io_ins_left[41] ;
 wire \ces_0_5_io_ins_left[42] ;
 wire \ces_0_5_io_ins_left[43] ;
 wire \ces_0_5_io_ins_left[44] ;
 wire \ces_0_5_io_ins_left[45] ;
 wire \ces_0_5_io_ins_left[46] ;
 wire \ces_0_5_io_ins_left[47] ;
 wire \ces_0_5_io_ins_left[48] ;
 wire \ces_0_5_io_ins_left[49] ;
 wire \ces_0_5_io_ins_left[4] ;
 wire \ces_0_5_io_ins_left[50] ;
 wire \ces_0_5_io_ins_left[51] ;
 wire \ces_0_5_io_ins_left[52] ;
 wire \ces_0_5_io_ins_left[53] ;
 wire \ces_0_5_io_ins_left[54] ;
 wire \ces_0_5_io_ins_left[55] ;
 wire \ces_0_5_io_ins_left[56] ;
 wire \ces_0_5_io_ins_left[57] ;
 wire \ces_0_5_io_ins_left[58] ;
 wire \ces_0_5_io_ins_left[59] ;
 wire \ces_0_5_io_ins_left[5] ;
 wire \ces_0_5_io_ins_left[60] ;
 wire \ces_0_5_io_ins_left[61] ;
 wire \ces_0_5_io_ins_left[62] ;
 wire \ces_0_5_io_ins_left[63] ;
 wire \ces_0_5_io_ins_left[6] ;
 wire \ces_0_5_io_ins_left[7] ;
 wire \ces_0_5_io_ins_left[8] ;
 wire \ces_0_5_io_ins_left[9] ;
 wire ces_0_5_io_lsbOuts_0;
 wire ces_0_5_io_lsbOuts_1;
 wire ces_0_5_io_lsbOuts_2;
 wire ces_0_5_io_lsbOuts_3;
 wire ces_0_5_io_lsbOuts_4;
 wire ces_0_5_io_lsbOuts_5;
 wire ces_0_5_io_lsbOuts_6;
 wire ces_0_5_io_lsbOuts_7;
 wire \ces_0_5_io_outs_right[0] ;
 wire \ces_0_5_io_outs_right[10] ;
 wire \ces_0_5_io_outs_right[11] ;
 wire \ces_0_5_io_outs_right[12] ;
 wire \ces_0_5_io_outs_right[13] ;
 wire \ces_0_5_io_outs_right[14] ;
 wire \ces_0_5_io_outs_right[15] ;
 wire \ces_0_5_io_outs_right[16] ;
 wire \ces_0_5_io_outs_right[17] ;
 wire \ces_0_5_io_outs_right[18] ;
 wire \ces_0_5_io_outs_right[19] ;
 wire \ces_0_5_io_outs_right[1] ;
 wire \ces_0_5_io_outs_right[20] ;
 wire \ces_0_5_io_outs_right[21] ;
 wire \ces_0_5_io_outs_right[22] ;
 wire \ces_0_5_io_outs_right[23] ;
 wire \ces_0_5_io_outs_right[24] ;
 wire \ces_0_5_io_outs_right[25] ;
 wire \ces_0_5_io_outs_right[26] ;
 wire \ces_0_5_io_outs_right[27] ;
 wire \ces_0_5_io_outs_right[28] ;
 wire \ces_0_5_io_outs_right[29] ;
 wire \ces_0_5_io_outs_right[2] ;
 wire \ces_0_5_io_outs_right[30] ;
 wire \ces_0_5_io_outs_right[31] ;
 wire \ces_0_5_io_outs_right[32] ;
 wire \ces_0_5_io_outs_right[33] ;
 wire \ces_0_5_io_outs_right[34] ;
 wire \ces_0_5_io_outs_right[35] ;
 wire \ces_0_5_io_outs_right[36] ;
 wire \ces_0_5_io_outs_right[37] ;
 wire \ces_0_5_io_outs_right[38] ;
 wire \ces_0_5_io_outs_right[39] ;
 wire \ces_0_5_io_outs_right[3] ;
 wire \ces_0_5_io_outs_right[40] ;
 wire \ces_0_5_io_outs_right[41] ;
 wire \ces_0_5_io_outs_right[42] ;
 wire \ces_0_5_io_outs_right[43] ;
 wire \ces_0_5_io_outs_right[44] ;
 wire \ces_0_5_io_outs_right[45] ;
 wire \ces_0_5_io_outs_right[46] ;
 wire \ces_0_5_io_outs_right[47] ;
 wire \ces_0_5_io_outs_right[48] ;
 wire \ces_0_5_io_outs_right[49] ;
 wire \ces_0_5_io_outs_right[4] ;
 wire \ces_0_5_io_outs_right[50] ;
 wire \ces_0_5_io_outs_right[51] ;
 wire \ces_0_5_io_outs_right[52] ;
 wire \ces_0_5_io_outs_right[53] ;
 wire \ces_0_5_io_outs_right[54] ;
 wire \ces_0_5_io_outs_right[55] ;
 wire \ces_0_5_io_outs_right[56] ;
 wire \ces_0_5_io_outs_right[57] ;
 wire \ces_0_5_io_outs_right[58] ;
 wire \ces_0_5_io_outs_right[59] ;
 wire \ces_0_5_io_outs_right[5] ;
 wire \ces_0_5_io_outs_right[60] ;
 wire \ces_0_5_io_outs_right[61] ;
 wire \ces_0_5_io_outs_right[62] ;
 wire \ces_0_5_io_outs_right[63] ;
 wire \ces_0_5_io_outs_right[6] ;
 wire \ces_0_5_io_outs_right[7] ;
 wire \ces_0_5_io_outs_right[8] ;
 wire \ces_0_5_io_outs_right[9] ;
 wire \ces_0_5_io_outs_up[0] ;
 wire \ces_0_5_io_outs_up[10] ;
 wire \ces_0_5_io_outs_up[11] ;
 wire \ces_0_5_io_outs_up[12] ;
 wire \ces_0_5_io_outs_up[13] ;
 wire \ces_0_5_io_outs_up[14] ;
 wire \ces_0_5_io_outs_up[15] ;
 wire \ces_0_5_io_outs_up[16] ;
 wire \ces_0_5_io_outs_up[17] ;
 wire \ces_0_5_io_outs_up[18] ;
 wire \ces_0_5_io_outs_up[19] ;
 wire \ces_0_5_io_outs_up[1] ;
 wire \ces_0_5_io_outs_up[20] ;
 wire \ces_0_5_io_outs_up[21] ;
 wire \ces_0_5_io_outs_up[22] ;
 wire \ces_0_5_io_outs_up[23] ;
 wire \ces_0_5_io_outs_up[24] ;
 wire \ces_0_5_io_outs_up[25] ;
 wire \ces_0_5_io_outs_up[26] ;
 wire \ces_0_5_io_outs_up[27] ;
 wire \ces_0_5_io_outs_up[28] ;
 wire \ces_0_5_io_outs_up[29] ;
 wire \ces_0_5_io_outs_up[2] ;
 wire \ces_0_5_io_outs_up[30] ;
 wire \ces_0_5_io_outs_up[31] ;
 wire \ces_0_5_io_outs_up[32] ;
 wire \ces_0_5_io_outs_up[33] ;
 wire \ces_0_5_io_outs_up[34] ;
 wire \ces_0_5_io_outs_up[35] ;
 wire \ces_0_5_io_outs_up[36] ;
 wire \ces_0_5_io_outs_up[37] ;
 wire \ces_0_5_io_outs_up[38] ;
 wire \ces_0_5_io_outs_up[39] ;
 wire \ces_0_5_io_outs_up[3] ;
 wire \ces_0_5_io_outs_up[40] ;
 wire \ces_0_5_io_outs_up[41] ;
 wire \ces_0_5_io_outs_up[42] ;
 wire \ces_0_5_io_outs_up[43] ;
 wire \ces_0_5_io_outs_up[44] ;
 wire \ces_0_5_io_outs_up[45] ;
 wire \ces_0_5_io_outs_up[46] ;
 wire \ces_0_5_io_outs_up[47] ;
 wire \ces_0_5_io_outs_up[48] ;
 wire \ces_0_5_io_outs_up[49] ;
 wire \ces_0_5_io_outs_up[4] ;
 wire \ces_0_5_io_outs_up[50] ;
 wire \ces_0_5_io_outs_up[51] ;
 wire \ces_0_5_io_outs_up[52] ;
 wire \ces_0_5_io_outs_up[53] ;
 wire \ces_0_5_io_outs_up[54] ;
 wire \ces_0_5_io_outs_up[55] ;
 wire \ces_0_5_io_outs_up[56] ;
 wire \ces_0_5_io_outs_up[57] ;
 wire \ces_0_5_io_outs_up[58] ;
 wire \ces_0_5_io_outs_up[59] ;
 wire \ces_0_5_io_outs_up[5] ;
 wire \ces_0_5_io_outs_up[60] ;
 wire \ces_0_5_io_outs_up[61] ;
 wire \ces_0_5_io_outs_up[62] ;
 wire \ces_0_5_io_outs_up[63] ;
 wire \ces_0_5_io_outs_up[6] ;
 wire \ces_0_5_io_outs_up[7] ;
 wire \ces_0_5_io_outs_up[8] ;
 wire \ces_0_5_io_outs_up[9] ;
 wire \ces_0_6_io_ins_down[0] ;
 wire \ces_0_6_io_ins_down[10] ;
 wire \ces_0_6_io_ins_down[11] ;
 wire \ces_0_6_io_ins_down[12] ;
 wire \ces_0_6_io_ins_down[13] ;
 wire \ces_0_6_io_ins_down[14] ;
 wire \ces_0_6_io_ins_down[15] ;
 wire \ces_0_6_io_ins_down[16] ;
 wire \ces_0_6_io_ins_down[17] ;
 wire \ces_0_6_io_ins_down[18] ;
 wire \ces_0_6_io_ins_down[19] ;
 wire \ces_0_6_io_ins_down[1] ;
 wire \ces_0_6_io_ins_down[20] ;
 wire \ces_0_6_io_ins_down[21] ;
 wire \ces_0_6_io_ins_down[22] ;
 wire \ces_0_6_io_ins_down[23] ;
 wire \ces_0_6_io_ins_down[24] ;
 wire \ces_0_6_io_ins_down[25] ;
 wire \ces_0_6_io_ins_down[26] ;
 wire \ces_0_6_io_ins_down[27] ;
 wire \ces_0_6_io_ins_down[28] ;
 wire \ces_0_6_io_ins_down[29] ;
 wire \ces_0_6_io_ins_down[2] ;
 wire \ces_0_6_io_ins_down[30] ;
 wire \ces_0_6_io_ins_down[31] ;
 wire \ces_0_6_io_ins_down[32] ;
 wire \ces_0_6_io_ins_down[33] ;
 wire \ces_0_6_io_ins_down[34] ;
 wire \ces_0_6_io_ins_down[35] ;
 wire \ces_0_6_io_ins_down[36] ;
 wire \ces_0_6_io_ins_down[37] ;
 wire \ces_0_6_io_ins_down[38] ;
 wire \ces_0_6_io_ins_down[39] ;
 wire \ces_0_6_io_ins_down[3] ;
 wire \ces_0_6_io_ins_down[40] ;
 wire \ces_0_6_io_ins_down[41] ;
 wire \ces_0_6_io_ins_down[42] ;
 wire \ces_0_6_io_ins_down[43] ;
 wire \ces_0_6_io_ins_down[44] ;
 wire \ces_0_6_io_ins_down[45] ;
 wire \ces_0_6_io_ins_down[46] ;
 wire \ces_0_6_io_ins_down[47] ;
 wire \ces_0_6_io_ins_down[48] ;
 wire \ces_0_6_io_ins_down[49] ;
 wire \ces_0_6_io_ins_down[4] ;
 wire \ces_0_6_io_ins_down[50] ;
 wire \ces_0_6_io_ins_down[51] ;
 wire \ces_0_6_io_ins_down[52] ;
 wire \ces_0_6_io_ins_down[53] ;
 wire \ces_0_6_io_ins_down[54] ;
 wire \ces_0_6_io_ins_down[55] ;
 wire \ces_0_6_io_ins_down[56] ;
 wire \ces_0_6_io_ins_down[57] ;
 wire \ces_0_6_io_ins_down[58] ;
 wire \ces_0_6_io_ins_down[59] ;
 wire \ces_0_6_io_ins_down[5] ;
 wire \ces_0_6_io_ins_down[60] ;
 wire \ces_0_6_io_ins_down[61] ;
 wire \ces_0_6_io_ins_down[62] ;
 wire \ces_0_6_io_ins_down[63] ;
 wire \ces_0_6_io_ins_down[6] ;
 wire \ces_0_6_io_ins_down[7] ;
 wire \ces_0_6_io_ins_down[8] ;
 wire \ces_0_6_io_ins_down[9] ;
 wire \ces_0_6_io_ins_left[0] ;
 wire \ces_0_6_io_ins_left[10] ;
 wire \ces_0_6_io_ins_left[11] ;
 wire \ces_0_6_io_ins_left[12] ;
 wire \ces_0_6_io_ins_left[13] ;
 wire \ces_0_6_io_ins_left[14] ;
 wire \ces_0_6_io_ins_left[15] ;
 wire \ces_0_6_io_ins_left[16] ;
 wire \ces_0_6_io_ins_left[17] ;
 wire \ces_0_6_io_ins_left[18] ;
 wire \ces_0_6_io_ins_left[19] ;
 wire \ces_0_6_io_ins_left[1] ;
 wire \ces_0_6_io_ins_left[20] ;
 wire \ces_0_6_io_ins_left[21] ;
 wire \ces_0_6_io_ins_left[22] ;
 wire \ces_0_6_io_ins_left[23] ;
 wire \ces_0_6_io_ins_left[24] ;
 wire \ces_0_6_io_ins_left[25] ;
 wire \ces_0_6_io_ins_left[26] ;
 wire \ces_0_6_io_ins_left[27] ;
 wire \ces_0_6_io_ins_left[28] ;
 wire \ces_0_6_io_ins_left[29] ;
 wire \ces_0_6_io_ins_left[2] ;
 wire \ces_0_6_io_ins_left[30] ;
 wire \ces_0_6_io_ins_left[31] ;
 wire \ces_0_6_io_ins_left[32] ;
 wire \ces_0_6_io_ins_left[33] ;
 wire \ces_0_6_io_ins_left[34] ;
 wire \ces_0_6_io_ins_left[35] ;
 wire \ces_0_6_io_ins_left[36] ;
 wire \ces_0_6_io_ins_left[37] ;
 wire \ces_0_6_io_ins_left[38] ;
 wire \ces_0_6_io_ins_left[39] ;
 wire \ces_0_6_io_ins_left[3] ;
 wire \ces_0_6_io_ins_left[40] ;
 wire \ces_0_6_io_ins_left[41] ;
 wire \ces_0_6_io_ins_left[42] ;
 wire \ces_0_6_io_ins_left[43] ;
 wire \ces_0_6_io_ins_left[44] ;
 wire \ces_0_6_io_ins_left[45] ;
 wire \ces_0_6_io_ins_left[46] ;
 wire \ces_0_6_io_ins_left[47] ;
 wire \ces_0_6_io_ins_left[48] ;
 wire \ces_0_6_io_ins_left[49] ;
 wire \ces_0_6_io_ins_left[4] ;
 wire \ces_0_6_io_ins_left[50] ;
 wire \ces_0_6_io_ins_left[51] ;
 wire \ces_0_6_io_ins_left[52] ;
 wire \ces_0_6_io_ins_left[53] ;
 wire \ces_0_6_io_ins_left[54] ;
 wire \ces_0_6_io_ins_left[55] ;
 wire \ces_0_6_io_ins_left[56] ;
 wire \ces_0_6_io_ins_left[57] ;
 wire \ces_0_6_io_ins_left[58] ;
 wire \ces_0_6_io_ins_left[59] ;
 wire \ces_0_6_io_ins_left[5] ;
 wire \ces_0_6_io_ins_left[60] ;
 wire \ces_0_6_io_ins_left[61] ;
 wire \ces_0_6_io_ins_left[62] ;
 wire \ces_0_6_io_ins_left[63] ;
 wire \ces_0_6_io_ins_left[6] ;
 wire \ces_0_6_io_ins_left[7] ;
 wire \ces_0_6_io_ins_left[8] ;
 wire \ces_0_6_io_ins_left[9] ;
 wire ces_0_6_io_lsbOuts_0;
 wire ces_0_6_io_lsbOuts_1;
 wire ces_0_6_io_lsbOuts_2;
 wire ces_0_6_io_lsbOuts_3;
 wire ces_0_6_io_lsbOuts_4;
 wire ces_0_6_io_lsbOuts_5;
 wire ces_0_6_io_lsbOuts_6;
 wire ces_0_6_io_lsbOuts_7;
 wire \ces_0_6_io_outs_right[0] ;
 wire \ces_0_6_io_outs_right[10] ;
 wire \ces_0_6_io_outs_right[11] ;
 wire \ces_0_6_io_outs_right[12] ;
 wire \ces_0_6_io_outs_right[13] ;
 wire \ces_0_6_io_outs_right[14] ;
 wire \ces_0_6_io_outs_right[15] ;
 wire \ces_0_6_io_outs_right[16] ;
 wire \ces_0_6_io_outs_right[17] ;
 wire \ces_0_6_io_outs_right[18] ;
 wire \ces_0_6_io_outs_right[19] ;
 wire \ces_0_6_io_outs_right[1] ;
 wire \ces_0_6_io_outs_right[20] ;
 wire \ces_0_6_io_outs_right[21] ;
 wire \ces_0_6_io_outs_right[22] ;
 wire \ces_0_6_io_outs_right[23] ;
 wire \ces_0_6_io_outs_right[24] ;
 wire \ces_0_6_io_outs_right[25] ;
 wire \ces_0_6_io_outs_right[26] ;
 wire \ces_0_6_io_outs_right[27] ;
 wire \ces_0_6_io_outs_right[28] ;
 wire \ces_0_6_io_outs_right[29] ;
 wire \ces_0_6_io_outs_right[2] ;
 wire \ces_0_6_io_outs_right[30] ;
 wire \ces_0_6_io_outs_right[31] ;
 wire \ces_0_6_io_outs_right[32] ;
 wire \ces_0_6_io_outs_right[33] ;
 wire \ces_0_6_io_outs_right[34] ;
 wire \ces_0_6_io_outs_right[35] ;
 wire \ces_0_6_io_outs_right[36] ;
 wire \ces_0_6_io_outs_right[37] ;
 wire \ces_0_6_io_outs_right[38] ;
 wire \ces_0_6_io_outs_right[39] ;
 wire \ces_0_6_io_outs_right[3] ;
 wire \ces_0_6_io_outs_right[40] ;
 wire \ces_0_6_io_outs_right[41] ;
 wire \ces_0_6_io_outs_right[42] ;
 wire \ces_0_6_io_outs_right[43] ;
 wire \ces_0_6_io_outs_right[44] ;
 wire \ces_0_6_io_outs_right[45] ;
 wire \ces_0_6_io_outs_right[46] ;
 wire \ces_0_6_io_outs_right[47] ;
 wire \ces_0_6_io_outs_right[48] ;
 wire \ces_0_6_io_outs_right[49] ;
 wire \ces_0_6_io_outs_right[4] ;
 wire \ces_0_6_io_outs_right[50] ;
 wire \ces_0_6_io_outs_right[51] ;
 wire \ces_0_6_io_outs_right[52] ;
 wire \ces_0_6_io_outs_right[53] ;
 wire \ces_0_6_io_outs_right[54] ;
 wire \ces_0_6_io_outs_right[55] ;
 wire \ces_0_6_io_outs_right[56] ;
 wire \ces_0_6_io_outs_right[57] ;
 wire \ces_0_6_io_outs_right[58] ;
 wire \ces_0_6_io_outs_right[59] ;
 wire \ces_0_6_io_outs_right[5] ;
 wire \ces_0_6_io_outs_right[60] ;
 wire \ces_0_6_io_outs_right[61] ;
 wire \ces_0_6_io_outs_right[62] ;
 wire \ces_0_6_io_outs_right[63] ;
 wire \ces_0_6_io_outs_right[6] ;
 wire \ces_0_6_io_outs_right[7] ;
 wire \ces_0_6_io_outs_right[8] ;
 wire \ces_0_6_io_outs_right[9] ;
 wire \ces_0_6_io_outs_up[0] ;
 wire \ces_0_6_io_outs_up[10] ;
 wire \ces_0_6_io_outs_up[11] ;
 wire \ces_0_6_io_outs_up[12] ;
 wire \ces_0_6_io_outs_up[13] ;
 wire \ces_0_6_io_outs_up[14] ;
 wire \ces_0_6_io_outs_up[15] ;
 wire \ces_0_6_io_outs_up[16] ;
 wire \ces_0_6_io_outs_up[17] ;
 wire \ces_0_6_io_outs_up[18] ;
 wire \ces_0_6_io_outs_up[19] ;
 wire \ces_0_6_io_outs_up[1] ;
 wire \ces_0_6_io_outs_up[20] ;
 wire \ces_0_6_io_outs_up[21] ;
 wire \ces_0_6_io_outs_up[22] ;
 wire \ces_0_6_io_outs_up[23] ;
 wire \ces_0_6_io_outs_up[24] ;
 wire \ces_0_6_io_outs_up[25] ;
 wire \ces_0_6_io_outs_up[26] ;
 wire \ces_0_6_io_outs_up[27] ;
 wire \ces_0_6_io_outs_up[28] ;
 wire \ces_0_6_io_outs_up[29] ;
 wire \ces_0_6_io_outs_up[2] ;
 wire \ces_0_6_io_outs_up[30] ;
 wire \ces_0_6_io_outs_up[31] ;
 wire \ces_0_6_io_outs_up[32] ;
 wire \ces_0_6_io_outs_up[33] ;
 wire \ces_0_6_io_outs_up[34] ;
 wire \ces_0_6_io_outs_up[35] ;
 wire \ces_0_6_io_outs_up[36] ;
 wire \ces_0_6_io_outs_up[37] ;
 wire \ces_0_6_io_outs_up[38] ;
 wire \ces_0_6_io_outs_up[39] ;
 wire \ces_0_6_io_outs_up[3] ;
 wire \ces_0_6_io_outs_up[40] ;
 wire \ces_0_6_io_outs_up[41] ;
 wire \ces_0_6_io_outs_up[42] ;
 wire \ces_0_6_io_outs_up[43] ;
 wire \ces_0_6_io_outs_up[44] ;
 wire \ces_0_6_io_outs_up[45] ;
 wire \ces_0_6_io_outs_up[46] ;
 wire \ces_0_6_io_outs_up[47] ;
 wire \ces_0_6_io_outs_up[48] ;
 wire \ces_0_6_io_outs_up[49] ;
 wire \ces_0_6_io_outs_up[4] ;
 wire \ces_0_6_io_outs_up[50] ;
 wire \ces_0_6_io_outs_up[51] ;
 wire \ces_0_6_io_outs_up[52] ;
 wire \ces_0_6_io_outs_up[53] ;
 wire \ces_0_6_io_outs_up[54] ;
 wire \ces_0_6_io_outs_up[55] ;
 wire \ces_0_6_io_outs_up[56] ;
 wire \ces_0_6_io_outs_up[57] ;
 wire \ces_0_6_io_outs_up[58] ;
 wire \ces_0_6_io_outs_up[59] ;
 wire \ces_0_6_io_outs_up[5] ;
 wire \ces_0_6_io_outs_up[60] ;
 wire \ces_0_6_io_outs_up[61] ;
 wire \ces_0_6_io_outs_up[62] ;
 wire \ces_0_6_io_outs_up[63] ;
 wire \ces_0_6_io_outs_up[6] ;
 wire \ces_0_6_io_outs_up[7] ;
 wire \ces_0_6_io_outs_up[8] ;
 wire \ces_0_6_io_outs_up[9] ;
 wire \ces_0_7_io_ins_down[0] ;
 wire \ces_0_7_io_ins_down[10] ;
 wire \ces_0_7_io_ins_down[11] ;
 wire \ces_0_7_io_ins_down[12] ;
 wire \ces_0_7_io_ins_down[13] ;
 wire \ces_0_7_io_ins_down[14] ;
 wire \ces_0_7_io_ins_down[15] ;
 wire \ces_0_7_io_ins_down[16] ;
 wire \ces_0_7_io_ins_down[17] ;
 wire \ces_0_7_io_ins_down[18] ;
 wire \ces_0_7_io_ins_down[19] ;
 wire \ces_0_7_io_ins_down[1] ;
 wire \ces_0_7_io_ins_down[20] ;
 wire \ces_0_7_io_ins_down[21] ;
 wire \ces_0_7_io_ins_down[22] ;
 wire \ces_0_7_io_ins_down[23] ;
 wire \ces_0_7_io_ins_down[24] ;
 wire \ces_0_7_io_ins_down[25] ;
 wire \ces_0_7_io_ins_down[26] ;
 wire \ces_0_7_io_ins_down[27] ;
 wire \ces_0_7_io_ins_down[28] ;
 wire \ces_0_7_io_ins_down[29] ;
 wire \ces_0_7_io_ins_down[2] ;
 wire \ces_0_7_io_ins_down[30] ;
 wire \ces_0_7_io_ins_down[31] ;
 wire \ces_0_7_io_ins_down[32] ;
 wire \ces_0_7_io_ins_down[33] ;
 wire \ces_0_7_io_ins_down[34] ;
 wire \ces_0_7_io_ins_down[35] ;
 wire \ces_0_7_io_ins_down[36] ;
 wire \ces_0_7_io_ins_down[37] ;
 wire \ces_0_7_io_ins_down[38] ;
 wire \ces_0_7_io_ins_down[39] ;
 wire \ces_0_7_io_ins_down[3] ;
 wire \ces_0_7_io_ins_down[40] ;
 wire \ces_0_7_io_ins_down[41] ;
 wire \ces_0_7_io_ins_down[42] ;
 wire \ces_0_7_io_ins_down[43] ;
 wire \ces_0_7_io_ins_down[44] ;
 wire \ces_0_7_io_ins_down[45] ;
 wire \ces_0_7_io_ins_down[46] ;
 wire \ces_0_7_io_ins_down[47] ;
 wire \ces_0_7_io_ins_down[48] ;
 wire \ces_0_7_io_ins_down[49] ;
 wire \ces_0_7_io_ins_down[4] ;
 wire \ces_0_7_io_ins_down[50] ;
 wire \ces_0_7_io_ins_down[51] ;
 wire \ces_0_7_io_ins_down[52] ;
 wire \ces_0_7_io_ins_down[53] ;
 wire \ces_0_7_io_ins_down[54] ;
 wire \ces_0_7_io_ins_down[55] ;
 wire \ces_0_7_io_ins_down[56] ;
 wire \ces_0_7_io_ins_down[57] ;
 wire \ces_0_7_io_ins_down[58] ;
 wire \ces_0_7_io_ins_down[59] ;
 wire \ces_0_7_io_ins_down[5] ;
 wire \ces_0_7_io_ins_down[60] ;
 wire \ces_0_7_io_ins_down[61] ;
 wire \ces_0_7_io_ins_down[62] ;
 wire \ces_0_7_io_ins_down[63] ;
 wire \ces_0_7_io_ins_down[6] ;
 wire \ces_0_7_io_ins_down[7] ;
 wire \ces_0_7_io_ins_down[8] ;
 wire \ces_0_7_io_ins_down[9] ;
 wire ces_0_7_io_lsbOuts_0;
 wire ces_0_7_io_lsbOuts_1;
 wire ces_0_7_io_lsbOuts_2;
 wire ces_0_7_io_lsbOuts_3;
 wire ces_0_7_io_lsbOuts_4;
 wire ces_0_7_io_lsbOuts_5;
 wire ces_0_7_io_lsbOuts_6;
 wire ces_0_7_io_lsbOuts_7;
 wire \ces_0_7_io_outs_up[0] ;
 wire \ces_0_7_io_outs_up[10] ;
 wire \ces_0_7_io_outs_up[11] ;
 wire \ces_0_7_io_outs_up[12] ;
 wire \ces_0_7_io_outs_up[13] ;
 wire \ces_0_7_io_outs_up[14] ;
 wire \ces_0_7_io_outs_up[15] ;
 wire \ces_0_7_io_outs_up[16] ;
 wire \ces_0_7_io_outs_up[17] ;
 wire \ces_0_7_io_outs_up[18] ;
 wire \ces_0_7_io_outs_up[19] ;
 wire \ces_0_7_io_outs_up[1] ;
 wire \ces_0_7_io_outs_up[20] ;
 wire \ces_0_7_io_outs_up[21] ;
 wire \ces_0_7_io_outs_up[22] ;
 wire \ces_0_7_io_outs_up[23] ;
 wire \ces_0_7_io_outs_up[24] ;
 wire \ces_0_7_io_outs_up[25] ;
 wire \ces_0_7_io_outs_up[26] ;
 wire \ces_0_7_io_outs_up[27] ;
 wire \ces_0_7_io_outs_up[28] ;
 wire \ces_0_7_io_outs_up[29] ;
 wire \ces_0_7_io_outs_up[2] ;
 wire \ces_0_7_io_outs_up[30] ;
 wire \ces_0_7_io_outs_up[31] ;
 wire \ces_0_7_io_outs_up[32] ;
 wire \ces_0_7_io_outs_up[33] ;
 wire \ces_0_7_io_outs_up[34] ;
 wire \ces_0_7_io_outs_up[35] ;
 wire \ces_0_7_io_outs_up[36] ;
 wire \ces_0_7_io_outs_up[37] ;
 wire \ces_0_7_io_outs_up[38] ;
 wire \ces_0_7_io_outs_up[39] ;
 wire \ces_0_7_io_outs_up[3] ;
 wire \ces_0_7_io_outs_up[40] ;
 wire \ces_0_7_io_outs_up[41] ;
 wire \ces_0_7_io_outs_up[42] ;
 wire \ces_0_7_io_outs_up[43] ;
 wire \ces_0_7_io_outs_up[44] ;
 wire \ces_0_7_io_outs_up[45] ;
 wire \ces_0_7_io_outs_up[46] ;
 wire \ces_0_7_io_outs_up[47] ;
 wire \ces_0_7_io_outs_up[48] ;
 wire \ces_0_7_io_outs_up[49] ;
 wire \ces_0_7_io_outs_up[4] ;
 wire \ces_0_7_io_outs_up[50] ;
 wire \ces_0_7_io_outs_up[51] ;
 wire \ces_0_7_io_outs_up[52] ;
 wire \ces_0_7_io_outs_up[53] ;
 wire \ces_0_7_io_outs_up[54] ;
 wire \ces_0_7_io_outs_up[55] ;
 wire \ces_0_7_io_outs_up[56] ;
 wire \ces_0_7_io_outs_up[57] ;
 wire \ces_0_7_io_outs_up[58] ;
 wire \ces_0_7_io_outs_up[59] ;
 wire \ces_0_7_io_outs_up[5] ;
 wire \ces_0_7_io_outs_up[60] ;
 wire \ces_0_7_io_outs_up[61] ;
 wire \ces_0_7_io_outs_up[62] ;
 wire \ces_0_7_io_outs_up[63] ;
 wire \ces_0_7_io_outs_up[6] ;
 wire \ces_0_7_io_outs_up[7] ;
 wire \ces_0_7_io_outs_up[8] ;
 wire \ces_0_7_io_outs_up[9] ;
 wire \ces_1_0_io_ins_down[0] ;
 wire \ces_1_0_io_ins_down[10] ;
 wire \ces_1_0_io_ins_down[11] ;
 wire \ces_1_0_io_ins_down[12] ;
 wire \ces_1_0_io_ins_down[13] ;
 wire \ces_1_0_io_ins_down[14] ;
 wire \ces_1_0_io_ins_down[15] ;
 wire \ces_1_0_io_ins_down[16] ;
 wire \ces_1_0_io_ins_down[17] ;
 wire \ces_1_0_io_ins_down[18] ;
 wire \ces_1_0_io_ins_down[19] ;
 wire \ces_1_0_io_ins_down[1] ;
 wire \ces_1_0_io_ins_down[20] ;
 wire \ces_1_0_io_ins_down[21] ;
 wire \ces_1_0_io_ins_down[22] ;
 wire \ces_1_0_io_ins_down[23] ;
 wire \ces_1_0_io_ins_down[24] ;
 wire \ces_1_0_io_ins_down[25] ;
 wire \ces_1_0_io_ins_down[26] ;
 wire \ces_1_0_io_ins_down[27] ;
 wire \ces_1_0_io_ins_down[28] ;
 wire \ces_1_0_io_ins_down[29] ;
 wire \ces_1_0_io_ins_down[2] ;
 wire \ces_1_0_io_ins_down[30] ;
 wire \ces_1_0_io_ins_down[31] ;
 wire \ces_1_0_io_ins_down[32] ;
 wire \ces_1_0_io_ins_down[33] ;
 wire \ces_1_0_io_ins_down[34] ;
 wire \ces_1_0_io_ins_down[35] ;
 wire \ces_1_0_io_ins_down[36] ;
 wire \ces_1_0_io_ins_down[37] ;
 wire \ces_1_0_io_ins_down[38] ;
 wire \ces_1_0_io_ins_down[39] ;
 wire \ces_1_0_io_ins_down[3] ;
 wire \ces_1_0_io_ins_down[40] ;
 wire \ces_1_0_io_ins_down[41] ;
 wire \ces_1_0_io_ins_down[42] ;
 wire \ces_1_0_io_ins_down[43] ;
 wire \ces_1_0_io_ins_down[44] ;
 wire \ces_1_0_io_ins_down[45] ;
 wire \ces_1_0_io_ins_down[46] ;
 wire \ces_1_0_io_ins_down[47] ;
 wire \ces_1_0_io_ins_down[48] ;
 wire \ces_1_0_io_ins_down[49] ;
 wire \ces_1_0_io_ins_down[4] ;
 wire \ces_1_0_io_ins_down[50] ;
 wire \ces_1_0_io_ins_down[51] ;
 wire \ces_1_0_io_ins_down[52] ;
 wire \ces_1_0_io_ins_down[53] ;
 wire \ces_1_0_io_ins_down[54] ;
 wire \ces_1_0_io_ins_down[55] ;
 wire \ces_1_0_io_ins_down[56] ;
 wire \ces_1_0_io_ins_down[57] ;
 wire \ces_1_0_io_ins_down[58] ;
 wire \ces_1_0_io_ins_down[59] ;
 wire \ces_1_0_io_ins_down[5] ;
 wire \ces_1_0_io_ins_down[60] ;
 wire \ces_1_0_io_ins_down[61] ;
 wire \ces_1_0_io_ins_down[62] ;
 wire \ces_1_0_io_ins_down[63] ;
 wire \ces_1_0_io_ins_down[6] ;
 wire \ces_1_0_io_ins_down[7] ;
 wire \ces_1_0_io_ins_down[8] ;
 wire \ces_1_0_io_ins_down[9] ;
 wire \ces_1_0_io_ins_left[0] ;
 wire \ces_1_0_io_ins_left[10] ;
 wire \ces_1_0_io_ins_left[11] ;
 wire \ces_1_0_io_ins_left[12] ;
 wire \ces_1_0_io_ins_left[13] ;
 wire \ces_1_0_io_ins_left[14] ;
 wire \ces_1_0_io_ins_left[15] ;
 wire \ces_1_0_io_ins_left[16] ;
 wire \ces_1_0_io_ins_left[17] ;
 wire \ces_1_0_io_ins_left[18] ;
 wire \ces_1_0_io_ins_left[19] ;
 wire \ces_1_0_io_ins_left[1] ;
 wire \ces_1_0_io_ins_left[20] ;
 wire \ces_1_0_io_ins_left[21] ;
 wire \ces_1_0_io_ins_left[22] ;
 wire \ces_1_0_io_ins_left[23] ;
 wire \ces_1_0_io_ins_left[24] ;
 wire \ces_1_0_io_ins_left[25] ;
 wire \ces_1_0_io_ins_left[26] ;
 wire \ces_1_0_io_ins_left[27] ;
 wire \ces_1_0_io_ins_left[28] ;
 wire \ces_1_0_io_ins_left[29] ;
 wire \ces_1_0_io_ins_left[2] ;
 wire \ces_1_0_io_ins_left[30] ;
 wire \ces_1_0_io_ins_left[31] ;
 wire \ces_1_0_io_ins_left[32] ;
 wire \ces_1_0_io_ins_left[33] ;
 wire \ces_1_0_io_ins_left[34] ;
 wire \ces_1_0_io_ins_left[35] ;
 wire \ces_1_0_io_ins_left[36] ;
 wire \ces_1_0_io_ins_left[37] ;
 wire \ces_1_0_io_ins_left[38] ;
 wire \ces_1_0_io_ins_left[39] ;
 wire \ces_1_0_io_ins_left[3] ;
 wire \ces_1_0_io_ins_left[40] ;
 wire \ces_1_0_io_ins_left[41] ;
 wire \ces_1_0_io_ins_left[42] ;
 wire \ces_1_0_io_ins_left[43] ;
 wire \ces_1_0_io_ins_left[44] ;
 wire \ces_1_0_io_ins_left[45] ;
 wire \ces_1_0_io_ins_left[46] ;
 wire \ces_1_0_io_ins_left[47] ;
 wire \ces_1_0_io_ins_left[48] ;
 wire \ces_1_0_io_ins_left[49] ;
 wire \ces_1_0_io_ins_left[4] ;
 wire \ces_1_0_io_ins_left[50] ;
 wire \ces_1_0_io_ins_left[51] ;
 wire \ces_1_0_io_ins_left[52] ;
 wire \ces_1_0_io_ins_left[53] ;
 wire \ces_1_0_io_ins_left[54] ;
 wire \ces_1_0_io_ins_left[55] ;
 wire \ces_1_0_io_ins_left[56] ;
 wire \ces_1_0_io_ins_left[57] ;
 wire \ces_1_0_io_ins_left[58] ;
 wire \ces_1_0_io_ins_left[59] ;
 wire \ces_1_0_io_ins_left[5] ;
 wire \ces_1_0_io_ins_left[60] ;
 wire \ces_1_0_io_ins_left[61] ;
 wire \ces_1_0_io_ins_left[62] ;
 wire \ces_1_0_io_ins_left[63] ;
 wire \ces_1_0_io_ins_left[6] ;
 wire \ces_1_0_io_ins_left[7] ;
 wire \ces_1_0_io_ins_left[8] ;
 wire \ces_1_0_io_ins_left[9] ;
 wire ces_1_0_io_lsbOuts_0;
 wire ces_1_0_io_lsbOuts_1;
 wire ces_1_0_io_lsbOuts_2;
 wire ces_1_0_io_lsbOuts_3;
 wire ces_1_0_io_lsbOuts_4;
 wire ces_1_0_io_lsbOuts_5;
 wire ces_1_0_io_lsbOuts_6;
 wire ces_1_0_io_lsbOuts_7;
 wire \ces_1_0_io_outs_right[0] ;
 wire \ces_1_0_io_outs_right[10] ;
 wire \ces_1_0_io_outs_right[11] ;
 wire \ces_1_0_io_outs_right[12] ;
 wire \ces_1_0_io_outs_right[13] ;
 wire \ces_1_0_io_outs_right[14] ;
 wire \ces_1_0_io_outs_right[15] ;
 wire \ces_1_0_io_outs_right[16] ;
 wire \ces_1_0_io_outs_right[17] ;
 wire \ces_1_0_io_outs_right[18] ;
 wire \ces_1_0_io_outs_right[19] ;
 wire \ces_1_0_io_outs_right[1] ;
 wire \ces_1_0_io_outs_right[20] ;
 wire \ces_1_0_io_outs_right[21] ;
 wire \ces_1_0_io_outs_right[22] ;
 wire \ces_1_0_io_outs_right[23] ;
 wire \ces_1_0_io_outs_right[24] ;
 wire \ces_1_0_io_outs_right[25] ;
 wire \ces_1_0_io_outs_right[26] ;
 wire \ces_1_0_io_outs_right[27] ;
 wire \ces_1_0_io_outs_right[28] ;
 wire \ces_1_0_io_outs_right[29] ;
 wire \ces_1_0_io_outs_right[2] ;
 wire \ces_1_0_io_outs_right[30] ;
 wire \ces_1_0_io_outs_right[31] ;
 wire \ces_1_0_io_outs_right[32] ;
 wire \ces_1_0_io_outs_right[33] ;
 wire \ces_1_0_io_outs_right[34] ;
 wire \ces_1_0_io_outs_right[35] ;
 wire \ces_1_0_io_outs_right[36] ;
 wire \ces_1_0_io_outs_right[37] ;
 wire \ces_1_0_io_outs_right[38] ;
 wire \ces_1_0_io_outs_right[39] ;
 wire \ces_1_0_io_outs_right[3] ;
 wire \ces_1_0_io_outs_right[40] ;
 wire \ces_1_0_io_outs_right[41] ;
 wire \ces_1_0_io_outs_right[42] ;
 wire \ces_1_0_io_outs_right[43] ;
 wire \ces_1_0_io_outs_right[44] ;
 wire \ces_1_0_io_outs_right[45] ;
 wire \ces_1_0_io_outs_right[46] ;
 wire \ces_1_0_io_outs_right[47] ;
 wire \ces_1_0_io_outs_right[48] ;
 wire \ces_1_0_io_outs_right[49] ;
 wire \ces_1_0_io_outs_right[4] ;
 wire \ces_1_0_io_outs_right[50] ;
 wire \ces_1_0_io_outs_right[51] ;
 wire \ces_1_0_io_outs_right[52] ;
 wire \ces_1_0_io_outs_right[53] ;
 wire \ces_1_0_io_outs_right[54] ;
 wire \ces_1_0_io_outs_right[55] ;
 wire \ces_1_0_io_outs_right[56] ;
 wire \ces_1_0_io_outs_right[57] ;
 wire \ces_1_0_io_outs_right[58] ;
 wire \ces_1_0_io_outs_right[59] ;
 wire \ces_1_0_io_outs_right[5] ;
 wire \ces_1_0_io_outs_right[60] ;
 wire \ces_1_0_io_outs_right[61] ;
 wire \ces_1_0_io_outs_right[62] ;
 wire \ces_1_0_io_outs_right[63] ;
 wire \ces_1_0_io_outs_right[6] ;
 wire \ces_1_0_io_outs_right[7] ;
 wire \ces_1_0_io_outs_right[8] ;
 wire \ces_1_0_io_outs_right[9] ;
 wire \ces_1_0_io_outs_up[0] ;
 wire \ces_1_0_io_outs_up[10] ;
 wire \ces_1_0_io_outs_up[11] ;
 wire \ces_1_0_io_outs_up[12] ;
 wire \ces_1_0_io_outs_up[13] ;
 wire \ces_1_0_io_outs_up[14] ;
 wire \ces_1_0_io_outs_up[15] ;
 wire \ces_1_0_io_outs_up[16] ;
 wire \ces_1_0_io_outs_up[17] ;
 wire \ces_1_0_io_outs_up[18] ;
 wire \ces_1_0_io_outs_up[19] ;
 wire \ces_1_0_io_outs_up[1] ;
 wire \ces_1_0_io_outs_up[20] ;
 wire \ces_1_0_io_outs_up[21] ;
 wire \ces_1_0_io_outs_up[22] ;
 wire \ces_1_0_io_outs_up[23] ;
 wire \ces_1_0_io_outs_up[24] ;
 wire \ces_1_0_io_outs_up[25] ;
 wire \ces_1_0_io_outs_up[26] ;
 wire \ces_1_0_io_outs_up[27] ;
 wire \ces_1_0_io_outs_up[28] ;
 wire \ces_1_0_io_outs_up[29] ;
 wire \ces_1_0_io_outs_up[2] ;
 wire \ces_1_0_io_outs_up[30] ;
 wire \ces_1_0_io_outs_up[31] ;
 wire \ces_1_0_io_outs_up[32] ;
 wire \ces_1_0_io_outs_up[33] ;
 wire \ces_1_0_io_outs_up[34] ;
 wire \ces_1_0_io_outs_up[35] ;
 wire \ces_1_0_io_outs_up[36] ;
 wire \ces_1_0_io_outs_up[37] ;
 wire \ces_1_0_io_outs_up[38] ;
 wire \ces_1_0_io_outs_up[39] ;
 wire \ces_1_0_io_outs_up[3] ;
 wire \ces_1_0_io_outs_up[40] ;
 wire \ces_1_0_io_outs_up[41] ;
 wire \ces_1_0_io_outs_up[42] ;
 wire \ces_1_0_io_outs_up[43] ;
 wire \ces_1_0_io_outs_up[44] ;
 wire \ces_1_0_io_outs_up[45] ;
 wire \ces_1_0_io_outs_up[46] ;
 wire \ces_1_0_io_outs_up[47] ;
 wire \ces_1_0_io_outs_up[48] ;
 wire \ces_1_0_io_outs_up[49] ;
 wire \ces_1_0_io_outs_up[4] ;
 wire \ces_1_0_io_outs_up[50] ;
 wire \ces_1_0_io_outs_up[51] ;
 wire \ces_1_0_io_outs_up[52] ;
 wire \ces_1_0_io_outs_up[53] ;
 wire \ces_1_0_io_outs_up[54] ;
 wire \ces_1_0_io_outs_up[55] ;
 wire \ces_1_0_io_outs_up[56] ;
 wire \ces_1_0_io_outs_up[57] ;
 wire \ces_1_0_io_outs_up[58] ;
 wire \ces_1_0_io_outs_up[59] ;
 wire \ces_1_0_io_outs_up[5] ;
 wire \ces_1_0_io_outs_up[60] ;
 wire \ces_1_0_io_outs_up[61] ;
 wire \ces_1_0_io_outs_up[62] ;
 wire \ces_1_0_io_outs_up[63] ;
 wire \ces_1_0_io_outs_up[6] ;
 wire \ces_1_0_io_outs_up[7] ;
 wire \ces_1_0_io_outs_up[8] ;
 wire \ces_1_0_io_outs_up[9] ;
 wire \ces_1_1_io_ins_down[0] ;
 wire \ces_1_1_io_ins_down[10] ;
 wire \ces_1_1_io_ins_down[11] ;
 wire \ces_1_1_io_ins_down[12] ;
 wire \ces_1_1_io_ins_down[13] ;
 wire \ces_1_1_io_ins_down[14] ;
 wire \ces_1_1_io_ins_down[15] ;
 wire \ces_1_1_io_ins_down[16] ;
 wire \ces_1_1_io_ins_down[17] ;
 wire \ces_1_1_io_ins_down[18] ;
 wire \ces_1_1_io_ins_down[19] ;
 wire \ces_1_1_io_ins_down[1] ;
 wire \ces_1_1_io_ins_down[20] ;
 wire \ces_1_1_io_ins_down[21] ;
 wire \ces_1_1_io_ins_down[22] ;
 wire \ces_1_1_io_ins_down[23] ;
 wire \ces_1_1_io_ins_down[24] ;
 wire \ces_1_1_io_ins_down[25] ;
 wire \ces_1_1_io_ins_down[26] ;
 wire \ces_1_1_io_ins_down[27] ;
 wire \ces_1_1_io_ins_down[28] ;
 wire \ces_1_1_io_ins_down[29] ;
 wire \ces_1_1_io_ins_down[2] ;
 wire \ces_1_1_io_ins_down[30] ;
 wire \ces_1_1_io_ins_down[31] ;
 wire \ces_1_1_io_ins_down[32] ;
 wire \ces_1_1_io_ins_down[33] ;
 wire \ces_1_1_io_ins_down[34] ;
 wire \ces_1_1_io_ins_down[35] ;
 wire \ces_1_1_io_ins_down[36] ;
 wire \ces_1_1_io_ins_down[37] ;
 wire \ces_1_1_io_ins_down[38] ;
 wire \ces_1_1_io_ins_down[39] ;
 wire \ces_1_1_io_ins_down[3] ;
 wire \ces_1_1_io_ins_down[40] ;
 wire \ces_1_1_io_ins_down[41] ;
 wire \ces_1_1_io_ins_down[42] ;
 wire \ces_1_1_io_ins_down[43] ;
 wire \ces_1_1_io_ins_down[44] ;
 wire \ces_1_1_io_ins_down[45] ;
 wire \ces_1_1_io_ins_down[46] ;
 wire \ces_1_1_io_ins_down[47] ;
 wire \ces_1_1_io_ins_down[48] ;
 wire \ces_1_1_io_ins_down[49] ;
 wire \ces_1_1_io_ins_down[4] ;
 wire \ces_1_1_io_ins_down[50] ;
 wire \ces_1_1_io_ins_down[51] ;
 wire \ces_1_1_io_ins_down[52] ;
 wire \ces_1_1_io_ins_down[53] ;
 wire \ces_1_1_io_ins_down[54] ;
 wire \ces_1_1_io_ins_down[55] ;
 wire \ces_1_1_io_ins_down[56] ;
 wire \ces_1_1_io_ins_down[57] ;
 wire \ces_1_1_io_ins_down[58] ;
 wire \ces_1_1_io_ins_down[59] ;
 wire \ces_1_1_io_ins_down[5] ;
 wire \ces_1_1_io_ins_down[60] ;
 wire \ces_1_1_io_ins_down[61] ;
 wire \ces_1_1_io_ins_down[62] ;
 wire \ces_1_1_io_ins_down[63] ;
 wire \ces_1_1_io_ins_down[6] ;
 wire \ces_1_1_io_ins_down[7] ;
 wire \ces_1_1_io_ins_down[8] ;
 wire \ces_1_1_io_ins_down[9] ;
 wire \ces_1_1_io_ins_left[0] ;
 wire \ces_1_1_io_ins_left[10] ;
 wire \ces_1_1_io_ins_left[11] ;
 wire \ces_1_1_io_ins_left[12] ;
 wire \ces_1_1_io_ins_left[13] ;
 wire \ces_1_1_io_ins_left[14] ;
 wire \ces_1_1_io_ins_left[15] ;
 wire \ces_1_1_io_ins_left[16] ;
 wire \ces_1_1_io_ins_left[17] ;
 wire \ces_1_1_io_ins_left[18] ;
 wire \ces_1_1_io_ins_left[19] ;
 wire \ces_1_1_io_ins_left[1] ;
 wire \ces_1_1_io_ins_left[20] ;
 wire \ces_1_1_io_ins_left[21] ;
 wire \ces_1_1_io_ins_left[22] ;
 wire \ces_1_1_io_ins_left[23] ;
 wire \ces_1_1_io_ins_left[24] ;
 wire \ces_1_1_io_ins_left[25] ;
 wire \ces_1_1_io_ins_left[26] ;
 wire \ces_1_1_io_ins_left[27] ;
 wire \ces_1_1_io_ins_left[28] ;
 wire \ces_1_1_io_ins_left[29] ;
 wire \ces_1_1_io_ins_left[2] ;
 wire \ces_1_1_io_ins_left[30] ;
 wire \ces_1_1_io_ins_left[31] ;
 wire \ces_1_1_io_ins_left[32] ;
 wire \ces_1_1_io_ins_left[33] ;
 wire \ces_1_1_io_ins_left[34] ;
 wire \ces_1_1_io_ins_left[35] ;
 wire \ces_1_1_io_ins_left[36] ;
 wire \ces_1_1_io_ins_left[37] ;
 wire \ces_1_1_io_ins_left[38] ;
 wire \ces_1_1_io_ins_left[39] ;
 wire \ces_1_1_io_ins_left[3] ;
 wire \ces_1_1_io_ins_left[40] ;
 wire \ces_1_1_io_ins_left[41] ;
 wire \ces_1_1_io_ins_left[42] ;
 wire \ces_1_1_io_ins_left[43] ;
 wire \ces_1_1_io_ins_left[44] ;
 wire \ces_1_1_io_ins_left[45] ;
 wire \ces_1_1_io_ins_left[46] ;
 wire \ces_1_1_io_ins_left[47] ;
 wire \ces_1_1_io_ins_left[48] ;
 wire \ces_1_1_io_ins_left[49] ;
 wire \ces_1_1_io_ins_left[4] ;
 wire \ces_1_1_io_ins_left[50] ;
 wire \ces_1_1_io_ins_left[51] ;
 wire \ces_1_1_io_ins_left[52] ;
 wire \ces_1_1_io_ins_left[53] ;
 wire \ces_1_1_io_ins_left[54] ;
 wire \ces_1_1_io_ins_left[55] ;
 wire \ces_1_1_io_ins_left[56] ;
 wire \ces_1_1_io_ins_left[57] ;
 wire \ces_1_1_io_ins_left[58] ;
 wire \ces_1_1_io_ins_left[59] ;
 wire \ces_1_1_io_ins_left[5] ;
 wire \ces_1_1_io_ins_left[60] ;
 wire \ces_1_1_io_ins_left[61] ;
 wire \ces_1_1_io_ins_left[62] ;
 wire \ces_1_1_io_ins_left[63] ;
 wire \ces_1_1_io_ins_left[6] ;
 wire \ces_1_1_io_ins_left[7] ;
 wire \ces_1_1_io_ins_left[8] ;
 wire \ces_1_1_io_ins_left[9] ;
 wire ces_1_1_io_lsbOuts_0;
 wire ces_1_1_io_lsbOuts_1;
 wire ces_1_1_io_lsbOuts_2;
 wire ces_1_1_io_lsbOuts_3;
 wire ces_1_1_io_lsbOuts_4;
 wire ces_1_1_io_lsbOuts_5;
 wire ces_1_1_io_lsbOuts_6;
 wire ces_1_1_io_lsbOuts_7;
 wire \ces_1_1_io_outs_right[0] ;
 wire \ces_1_1_io_outs_right[10] ;
 wire \ces_1_1_io_outs_right[11] ;
 wire \ces_1_1_io_outs_right[12] ;
 wire \ces_1_1_io_outs_right[13] ;
 wire \ces_1_1_io_outs_right[14] ;
 wire \ces_1_1_io_outs_right[15] ;
 wire \ces_1_1_io_outs_right[16] ;
 wire \ces_1_1_io_outs_right[17] ;
 wire \ces_1_1_io_outs_right[18] ;
 wire \ces_1_1_io_outs_right[19] ;
 wire \ces_1_1_io_outs_right[1] ;
 wire \ces_1_1_io_outs_right[20] ;
 wire \ces_1_1_io_outs_right[21] ;
 wire \ces_1_1_io_outs_right[22] ;
 wire \ces_1_1_io_outs_right[23] ;
 wire \ces_1_1_io_outs_right[24] ;
 wire \ces_1_1_io_outs_right[25] ;
 wire \ces_1_1_io_outs_right[26] ;
 wire \ces_1_1_io_outs_right[27] ;
 wire \ces_1_1_io_outs_right[28] ;
 wire \ces_1_1_io_outs_right[29] ;
 wire \ces_1_1_io_outs_right[2] ;
 wire \ces_1_1_io_outs_right[30] ;
 wire \ces_1_1_io_outs_right[31] ;
 wire \ces_1_1_io_outs_right[32] ;
 wire \ces_1_1_io_outs_right[33] ;
 wire \ces_1_1_io_outs_right[34] ;
 wire \ces_1_1_io_outs_right[35] ;
 wire \ces_1_1_io_outs_right[36] ;
 wire \ces_1_1_io_outs_right[37] ;
 wire \ces_1_1_io_outs_right[38] ;
 wire \ces_1_1_io_outs_right[39] ;
 wire \ces_1_1_io_outs_right[3] ;
 wire \ces_1_1_io_outs_right[40] ;
 wire \ces_1_1_io_outs_right[41] ;
 wire \ces_1_1_io_outs_right[42] ;
 wire \ces_1_1_io_outs_right[43] ;
 wire \ces_1_1_io_outs_right[44] ;
 wire \ces_1_1_io_outs_right[45] ;
 wire \ces_1_1_io_outs_right[46] ;
 wire \ces_1_1_io_outs_right[47] ;
 wire \ces_1_1_io_outs_right[48] ;
 wire \ces_1_1_io_outs_right[49] ;
 wire \ces_1_1_io_outs_right[4] ;
 wire \ces_1_1_io_outs_right[50] ;
 wire \ces_1_1_io_outs_right[51] ;
 wire \ces_1_1_io_outs_right[52] ;
 wire \ces_1_1_io_outs_right[53] ;
 wire \ces_1_1_io_outs_right[54] ;
 wire \ces_1_1_io_outs_right[55] ;
 wire \ces_1_1_io_outs_right[56] ;
 wire \ces_1_1_io_outs_right[57] ;
 wire \ces_1_1_io_outs_right[58] ;
 wire \ces_1_1_io_outs_right[59] ;
 wire \ces_1_1_io_outs_right[5] ;
 wire \ces_1_1_io_outs_right[60] ;
 wire \ces_1_1_io_outs_right[61] ;
 wire \ces_1_1_io_outs_right[62] ;
 wire \ces_1_1_io_outs_right[63] ;
 wire \ces_1_1_io_outs_right[6] ;
 wire \ces_1_1_io_outs_right[7] ;
 wire \ces_1_1_io_outs_right[8] ;
 wire \ces_1_1_io_outs_right[9] ;
 wire \ces_1_1_io_outs_up[0] ;
 wire \ces_1_1_io_outs_up[10] ;
 wire \ces_1_1_io_outs_up[11] ;
 wire \ces_1_1_io_outs_up[12] ;
 wire \ces_1_1_io_outs_up[13] ;
 wire \ces_1_1_io_outs_up[14] ;
 wire \ces_1_1_io_outs_up[15] ;
 wire \ces_1_1_io_outs_up[16] ;
 wire \ces_1_1_io_outs_up[17] ;
 wire \ces_1_1_io_outs_up[18] ;
 wire \ces_1_1_io_outs_up[19] ;
 wire \ces_1_1_io_outs_up[1] ;
 wire \ces_1_1_io_outs_up[20] ;
 wire \ces_1_1_io_outs_up[21] ;
 wire \ces_1_1_io_outs_up[22] ;
 wire \ces_1_1_io_outs_up[23] ;
 wire \ces_1_1_io_outs_up[24] ;
 wire \ces_1_1_io_outs_up[25] ;
 wire \ces_1_1_io_outs_up[26] ;
 wire \ces_1_1_io_outs_up[27] ;
 wire \ces_1_1_io_outs_up[28] ;
 wire \ces_1_1_io_outs_up[29] ;
 wire \ces_1_1_io_outs_up[2] ;
 wire \ces_1_1_io_outs_up[30] ;
 wire \ces_1_1_io_outs_up[31] ;
 wire \ces_1_1_io_outs_up[32] ;
 wire \ces_1_1_io_outs_up[33] ;
 wire \ces_1_1_io_outs_up[34] ;
 wire \ces_1_1_io_outs_up[35] ;
 wire \ces_1_1_io_outs_up[36] ;
 wire \ces_1_1_io_outs_up[37] ;
 wire \ces_1_1_io_outs_up[38] ;
 wire \ces_1_1_io_outs_up[39] ;
 wire \ces_1_1_io_outs_up[3] ;
 wire \ces_1_1_io_outs_up[40] ;
 wire \ces_1_1_io_outs_up[41] ;
 wire \ces_1_1_io_outs_up[42] ;
 wire \ces_1_1_io_outs_up[43] ;
 wire \ces_1_1_io_outs_up[44] ;
 wire \ces_1_1_io_outs_up[45] ;
 wire \ces_1_1_io_outs_up[46] ;
 wire \ces_1_1_io_outs_up[47] ;
 wire \ces_1_1_io_outs_up[48] ;
 wire \ces_1_1_io_outs_up[49] ;
 wire \ces_1_1_io_outs_up[4] ;
 wire \ces_1_1_io_outs_up[50] ;
 wire \ces_1_1_io_outs_up[51] ;
 wire \ces_1_1_io_outs_up[52] ;
 wire \ces_1_1_io_outs_up[53] ;
 wire \ces_1_1_io_outs_up[54] ;
 wire \ces_1_1_io_outs_up[55] ;
 wire \ces_1_1_io_outs_up[56] ;
 wire \ces_1_1_io_outs_up[57] ;
 wire \ces_1_1_io_outs_up[58] ;
 wire \ces_1_1_io_outs_up[59] ;
 wire \ces_1_1_io_outs_up[5] ;
 wire \ces_1_1_io_outs_up[60] ;
 wire \ces_1_1_io_outs_up[61] ;
 wire \ces_1_1_io_outs_up[62] ;
 wire \ces_1_1_io_outs_up[63] ;
 wire \ces_1_1_io_outs_up[6] ;
 wire \ces_1_1_io_outs_up[7] ;
 wire \ces_1_1_io_outs_up[8] ;
 wire \ces_1_1_io_outs_up[9] ;
 wire \ces_1_2_io_ins_down[0] ;
 wire \ces_1_2_io_ins_down[10] ;
 wire \ces_1_2_io_ins_down[11] ;
 wire \ces_1_2_io_ins_down[12] ;
 wire \ces_1_2_io_ins_down[13] ;
 wire \ces_1_2_io_ins_down[14] ;
 wire \ces_1_2_io_ins_down[15] ;
 wire \ces_1_2_io_ins_down[16] ;
 wire \ces_1_2_io_ins_down[17] ;
 wire \ces_1_2_io_ins_down[18] ;
 wire \ces_1_2_io_ins_down[19] ;
 wire \ces_1_2_io_ins_down[1] ;
 wire \ces_1_2_io_ins_down[20] ;
 wire \ces_1_2_io_ins_down[21] ;
 wire \ces_1_2_io_ins_down[22] ;
 wire \ces_1_2_io_ins_down[23] ;
 wire \ces_1_2_io_ins_down[24] ;
 wire \ces_1_2_io_ins_down[25] ;
 wire \ces_1_2_io_ins_down[26] ;
 wire \ces_1_2_io_ins_down[27] ;
 wire \ces_1_2_io_ins_down[28] ;
 wire \ces_1_2_io_ins_down[29] ;
 wire \ces_1_2_io_ins_down[2] ;
 wire \ces_1_2_io_ins_down[30] ;
 wire \ces_1_2_io_ins_down[31] ;
 wire \ces_1_2_io_ins_down[32] ;
 wire \ces_1_2_io_ins_down[33] ;
 wire \ces_1_2_io_ins_down[34] ;
 wire \ces_1_2_io_ins_down[35] ;
 wire \ces_1_2_io_ins_down[36] ;
 wire \ces_1_2_io_ins_down[37] ;
 wire \ces_1_2_io_ins_down[38] ;
 wire \ces_1_2_io_ins_down[39] ;
 wire \ces_1_2_io_ins_down[3] ;
 wire \ces_1_2_io_ins_down[40] ;
 wire \ces_1_2_io_ins_down[41] ;
 wire \ces_1_2_io_ins_down[42] ;
 wire \ces_1_2_io_ins_down[43] ;
 wire \ces_1_2_io_ins_down[44] ;
 wire \ces_1_2_io_ins_down[45] ;
 wire \ces_1_2_io_ins_down[46] ;
 wire \ces_1_2_io_ins_down[47] ;
 wire \ces_1_2_io_ins_down[48] ;
 wire \ces_1_2_io_ins_down[49] ;
 wire \ces_1_2_io_ins_down[4] ;
 wire \ces_1_2_io_ins_down[50] ;
 wire \ces_1_2_io_ins_down[51] ;
 wire \ces_1_2_io_ins_down[52] ;
 wire \ces_1_2_io_ins_down[53] ;
 wire \ces_1_2_io_ins_down[54] ;
 wire \ces_1_2_io_ins_down[55] ;
 wire \ces_1_2_io_ins_down[56] ;
 wire \ces_1_2_io_ins_down[57] ;
 wire \ces_1_2_io_ins_down[58] ;
 wire \ces_1_2_io_ins_down[59] ;
 wire \ces_1_2_io_ins_down[5] ;
 wire \ces_1_2_io_ins_down[60] ;
 wire \ces_1_2_io_ins_down[61] ;
 wire \ces_1_2_io_ins_down[62] ;
 wire \ces_1_2_io_ins_down[63] ;
 wire \ces_1_2_io_ins_down[6] ;
 wire \ces_1_2_io_ins_down[7] ;
 wire \ces_1_2_io_ins_down[8] ;
 wire \ces_1_2_io_ins_down[9] ;
 wire \ces_1_2_io_ins_left[0] ;
 wire \ces_1_2_io_ins_left[10] ;
 wire \ces_1_2_io_ins_left[11] ;
 wire \ces_1_2_io_ins_left[12] ;
 wire \ces_1_2_io_ins_left[13] ;
 wire \ces_1_2_io_ins_left[14] ;
 wire \ces_1_2_io_ins_left[15] ;
 wire \ces_1_2_io_ins_left[16] ;
 wire \ces_1_2_io_ins_left[17] ;
 wire \ces_1_2_io_ins_left[18] ;
 wire \ces_1_2_io_ins_left[19] ;
 wire \ces_1_2_io_ins_left[1] ;
 wire \ces_1_2_io_ins_left[20] ;
 wire \ces_1_2_io_ins_left[21] ;
 wire \ces_1_2_io_ins_left[22] ;
 wire \ces_1_2_io_ins_left[23] ;
 wire \ces_1_2_io_ins_left[24] ;
 wire \ces_1_2_io_ins_left[25] ;
 wire \ces_1_2_io_ins_left[26] ;
 wire \ces_1_2_io_ins_left[27] ;
 wire \ces_1_2_io_ins_left[28] ;
 wire \ces_1_2_io_ins_left[29] ;
 wire \ces_1_2_io_ins_left[2] ;
 wire \ces_1_2_io_ins_left[30] ;
 wire \ces_1_2_io_ins_left[31] ;
 wire \ces_1_2_io_ins_left[32] ;
 wire \ces_1_2_io_ins_left[33] ;
 wire \ces_1_2_io_ins_left[34] ;
 wire \ces_1_2_io_ins_left[35] ;
 wire \ces_1_2_io_ins_left[36] ;
 wire \ces_1_2_io_ins_left[37] ;
 wire \ces_1_2_io_ins_left[38] ;
 wire \ces_1_2_io_ins_left[39] ;
 wire \ces_1_2_io_ins_left[3] ;
 wire \ces_1_2_io_ins_left[40] ;
 wire \ces_1_2_io_ins_left[41] ;
 wire \ces_1_2_io_ins_left[42] ;
 wire \ces_1_2_io_ins_left[43] ;
 wire \ces_1_2_io_ins_left[44] ;
 wire \ces_1_2_io_ins_left[45] ;
 wire \ces_1_2_io_ins_left[46] ;
 wire \ces_1_2_io_ins_left[47] ;
 wire \ces_1_2_io_ins_left[48] ;
 wire \ces_1_2_io_ins_left[49] ;
 wire \ces_1_2_io_ins_left[4] ;
 wire \ces_1_2_io_ins_left[50] ;
 wire \ces_1_2_io_ins_left[51] ;
 wire \ces_1_2_io_ins_left[52] ;
 wire \ces_1_2_io_ins_left[53] ;
 wire \ces_1_2_io_ins_left[54] ;
 wire \ces_1_2_io_ins_left[55] ;
 wire \ces_1_2_io_ins_left[56] ;
 wire \ces_1_2_io_ins_left[57] ;
 wire \ces_1_2_io_ins_left[58] ;
 wire \ces_1_2_io_ins_left[59] ;
 wire \ces_1_2_io_ins_left[5] ;
 wire \ces_1_2_io_ins_left[60] ;
 wire \ces_1_2_io_ins_left[61] ;
 wire \ces_1_2_io_ins_left[62] ;
 wire \ces_1_2_io_ins_left[63] ;
 wire \ces_1_2_io_ins_left[6] ;
 wire \ces_1_2_io_ins_left[7] ;
 wire \ces_1_2_io_ins_left[8] ;
 wire \ces_1_2_io_ins_left[9] ;
 wire ces_1_2_io_lsbOuts_0;
 wire ces_1_2_io_lsbOuts_1;
 wire ces_1_2_io_lsbOuts_2;
 wire ces_1_2_io_lsbOuts_3;
 wire ces_1_2_io_lsbOuts_4;
 wire ces_1_2_io_lsbOuts_5;
 wire ces_1_2_io_lsbOuts_6;
 wire ces_1_2_io_lsbOuts_7;
 wire \ces_1_2_io_outs_right[0] ;
 wire \ces_1_2_io_outs_right[10] ;
 wire \ces_1_2_io_outs_right[11] ;
 wire \ces_1_2_io_outs_right[12] ;
 wire \ces_1_2_io_outs_right[13] ;
 wire \ces_1_2_io_outs_right[14] ;
 wire \ces_1_2_io_outs_right[15] ;
 wire \ces_1_2_io_outs_right[16] ;
 wire \ces_1_2_io_outs_right[17] ;
 wire \ces_1_2_io_outs_right[18] ;
 wire \ces_1_2_io_outs_right[19] ;
 wire \ces_1_2_io_outs_right[1] ;
 wire \ces_1_2_io_outs_right[20] ;
 wire \ces_1_2_io_outs_right[21] ;
 wire \ces_1_2_io_outs_right[22] ;
 wire \ces_1_2_io_outs_right[23] ;
 wire \ces_1_2_io_outs_right[24] ;
 wire \ces_1_2_io_outs_right[25] ;
 wire \ces_1_2_io_outs_right[26] ;
 wire \ces_1_2_io_outs_right[27] ;
 wire \ces_1_2_io_outs_right[28] ;
 wire \ces_1_2_io_outs_right[29] ;
 wire \ces_1_2_io_outs_right[2] ;
 wire \ces_1_2_io_outs_right[30] ;
 wire \ces_1_2_io_outs_right[31] ;
 wire \ces_1_2_io_outs_right[32] ;
 wire \ces_1_2_io_outs_right[33] ;
 wire \ces_1_2_io_outs_right[34] ;
 wire \ces_1_2_io_outs_right[35] ;
 wire \ces_1_2_io_outs_right[36] ;
 wire \ces_1_2_io_outs_right[37] ;
 wire \ces_1_2_io_outs_right[38] ;
 wire \ces_1_2_io_outs_right[39] ;
 wire \ces_1_2_io_outs_right[3] ;
 wire \ces_1_2_io_outs_right[40] ;
 wire \ces_1_2_io_outs_right[41] ;
 wire \ces_1_2_io_outs_right[42] ;
 wire \ces_1_2_io_outs_right[43] ;
 wire \ces_1_2_io_outs_right[44] ;
 wire \ces_1_2_io_outs_right[45] ;
 wire \ces_1_2_io_outs_right[46] ;
 wire \ces_1_2_io_outs_right[47] ;
 wire \ces_1_2_io_outs_right[48] ;
 wire \ces_1_2_io_outs_right[49] ;
 wire \ces_1_2_io_outs_right[4] ;
 wire \ces_1_2_io_outs_right[50] ;
 wire \ces_1_2_io_outs_right[51] ;
 wire \ces_1_2_io_outs_right[52] ;
 wire \ces_1_2_io_outs_right[53] ;
 wire \ces_1_2_io_outs_right[54] ;
 wire \ces_1_2_io_outs_right[55] ;
 wire \ces_1_2_io_outs_right[56] ;
 wire \ces_1_2_io_outs_right[57] ;
 wire \ces_1_2_io_outs_right[58] ;
 wire \ces_1_2_io_outs_right[59] ;
 wire \ces_1_2_io_outs_right[5] ;
 wire \ces_1_2_io_outs_right[60] ;
 wire \ces_1_2_io_outs_right[61] ;
 wire \ces_1_2_io_outs_right[62] ;
 wire \ces_1_2_io_outs_right[63] ;
 wire \ces_1_2_io_outs_right[6] ;
 wire \ces_1_2_io_outs_right[7] ;
 wire \ces_1_2_io_outs_right[8] ;
 wire \ces_1_2_io_outs_right[9] ;
 wire \ces_1_2_io_outs_up[0] ;
 wire \ces_1_2_io_outs_up[10] ;
 wire \ces_1_2_io_outs_up[11] ;
 wire \ces_1_2_io_outs_up[12] ;
 wire \ces_1_2_io_outs_up[13] ;
 wire \ces_1_2_io_outs_up[14] ;
 wire \ces_1_2_io_outs_up[15] ;
 wire \ces_1_2_io_outs_up[16] ;
 wire \ces_1_2_io_outs_up[17] ;
 wire \ces_1_2_io_outs_up[18] ;
 wire \ces_1_2_io_outs_up[19] ;
 wire \ces_1_2_io_outs_up[1] ;
 wire \ces_1_2_io_outs_up[20] ;
 wire \ces_1_2_io_outs_up[21] ;
 wire \ces_1_2_io_outs_up[22] ;
 wire \ces_1_2_io_outs_up[23] ;
 wire \ces_1_2_io_outs_up[24] ;
 wire \ces_1_2_io_outs_up[25] ;
 wire \ces_1_2_io_outs_up[26] ;
 wire \ces_1_2_io_outs_up[27] ;
 wire \ces_1_2_io_outs_up[28] ;
 wire \ces_1_2_io_outs_up[29] ;
 wire \ces_1_2_io_outs_up[2] ;
 wire \ces_1_2_io_outs_up[30] ;
 wire \ces_1_2_io_outs_up[31] ;
 wire \ces_1_2_io_outs_up[32] ;
 wire \ces_1_2_io_outs_up[33] ;
 wire \ces_1_2_io_outs_up[34] ;
 wire \ces_1_2_io_outs_up[35] ;
 wire \ces_1_2_io_outs_up[36] ;
 wire \ces_1_2_io_outs_up[37] ;
 wire \ces_1_2_io_outs_up[38] ;
 wire \ces_1_2_io_outs_up[39] ;
 wire \ces_1_2_io_outs_up[3] ;
 wire \ces_1_2_io_outs_up[40] ;
 wire \ces_1_2_io_outs_up[41] ;
 wire \ces_1_2_io_outs_up[42] ;
 wire \ces_1_2_io_outs_up[43] ;
 wire \ces_1_2_io_outs_up[44] ;
 wire \ces_1_2_io_outs_up[45] ;
 wire \ces_1_2_io_outs_up[46] ;
 wire \ces_1_2_io_outs_up[47] ;
 wire \ces_1_2_io_outs_up[48] ;
 wire \ces_1_2_io_outs_up[49] ;
 wire \ces_1_2_io_outs_up[4] ;
 wire \ces_1_2_io_outs_up[50] ;
 wire \ces_1_2_io_outs_up[51] ;
 wire \ces_1_2_io_outs_up[52] ;
 wire \ces_1_2_io_outs_up[53] ;
 wire \ces_1_2_io_outs_up[54] ;
 wire \ces_1_2_io_outs_up[55] ;
 wire \ces_1_2_io_outs_up[56] ;
 wire \ces_1_2_io_outs_up[57] ;
 wire \ces_1_2_io_outs_up[58] ;
 wire \ces_1_2_io_outs_up[59] ;
 wire \ces_1_2_io_outs_up[5] ;
 wire \ces_1_2_io_outs_up[60] ;
 wire \ces_1_2_io_outs_up[61] ;
 wire \ces_1_2_io_outs_up[62] ;
 wire \ces_1_2_io_outs_up[63] ;
 wire \ces_1_2_io_outs_up[6] ;
 wire \ces_1_2_io_outs_up[7] ;
 wire \ces_1_2_io_outs_up[8] ;
 wire \ces_1_2_io_outs_up[9] ;
 wire \ces_1_3_io_ins_down[0] ;
 wire \ces_1_3_io_ins_down[10] ;
 wire \ces_1_3_io_ins_down[11] ;
 wire \ces_1_3_io_ins_down[12] ;
 wire \ces_1_3_io_ins_down[13] ;
 wire \ces_1_3_io_ins_down[14] ;
 wire \ces_1_3_io_ins_down[15] ;
 wire \ces_1_3_io_ins_down[16] ;
 wire \ces_1_3_io_ins_down[17] ;
 wire \ces_1_3_io_ins_down[18] ;
 wire \ces_1_3_io_ins_down[19] ;
 wire \ces_1_3_io_ins_down[1] ;
 wire \ces_1_3_io_ins_down[20] ;
 wire \ces_1_3_io_ins_down[21] ;
 wire \ces_1_3_io_ins_down[22] ;
 wire \ces_1_3_io_ins_down[23] ;
 wire \ces_1_3_io_ins_down[24] ;
 wire \ces_1_3_io_ins_down[25] ;
 wire \ces_1_3_io_ins_down[26] ;
 wire \ces_1_3_io_ins_down[27] ;
 wire \ces_1_3_io_ins_down[28] ;
 wire \ces_1_3_io_ins_down[29] ;
 wire \ces_1_3_io_ins_down[2] ;
 wire \ces_1_3_io_ins_down[30] ;
 wire \ces_1_3_io_ins_down[31] ;
 wire \ces_1_3_io_ins_down[32] ;
 wire \ces_1_3_io_ins_down[33] ;
 wire \ces_1_3_io_ins_down[34] ;
 wire \ces_1_3_io_ins_down[35] ;
 wire \ces_1_3_io_ins_down[36] ;
 wire \ces_1_3_io_ins_down[37] ;
 wire \ces_1_3_io_ins_down[38] ;
 wire \ces_1_3_io_ins_down[39] ;
 wire \ces_1_3_io_ins_down[3] ;
 wire \ces_1_3_io_ins_down[40] ;
 wire \ces_1_3_io_ins_down[41] ;
 wire \ces_1_3_io_ins_down[42] ;
 wire \ces_1_3_io_ins_down[43] ;
 wire \ces_1_3_io_ins_down[44] ;
 wire \ces_1_3_io_ins_down[45] ;
 wire \ces_1_3_io_ins_down[46] ;
 wire \ces_1_3_io_ins_down[47] ;
 wire \ces_1_3_io_ins_down[48] ;
 wire \ces_1_3_io_ins_down[49] ;
 wire \ces_1_3_io_ins_down[4] ;
 wire \ces_1_3_io_ins_down[50] ;
 wire \ces_1_3_io_ins_down[51] ;
 wire \ces_1_3_io_ins_down[52] ;
 wire \ces_1_3_io_ins_down[53] ;
 wire \ces_1_3_io_ins_down[54] ;
 wire \ces_1_3_io_ins_down[55] ;
 wire \ces_1_3_io_ins_down[56] ;
 wire \ces_1_3_io_ins_down[57] ;
 wire \ces_1_3_io_ins_down[58] ;
 wire \ces_1_3_io_ins_down[59] ;
 wire \ces_1_3_io_ins_down[5] ;
 wire \ces_1_3_io_ins_down[60] ;
 wire \ces_1_3_io_ins_down[61] ;
 wire \ces_1_3_io_ins_down[62] ;
 wire \ces_1_3_io_ins_down[63] ;
 wire \ces_1_3_io_ins_down[6] ;
 wire \ces_1_3_io_ins_down[7] ;
 wire \ces_1_3_io_ins_down[8] ;
 wire \ces_1_3_io_ins_down[9] ;
 wire \ces_1_3_io_ins_left[0] ;
 wire \ces_1_3_io_ins_left[10] ;
 wire \ces_1_3_io_ins_left[11] ;
 wire \ces_1_3_io_ins_left[12] ;
 wire \ces_1_3_io_ins_left[13] ;
 wire \ces_1_3_io_ins_left[14] ;
 wire \ces_1_3_io_ins_left[15] ;
 wire \ces_1_3_io_ins_left[16] ;
 wire \ces_1_3_io_ins_left[17] ;
 wire \ces_1_3_io_ins_left[18] ;
 wire \ces_1_3_io_ins_left[19] ;
 wire \ces_1_3_io_ins_left[1] ;
 wire \ces_1_3_io_ins_left[20] ;
 wire \ces_1_3_io_ins_left[21] ;
 wire \ces_1_3_io_ins_left[22] ;
 wire \ces_1_3_io_ins_left[23] ;
 wire \ces_1_3_io_ins_left[24] ;
 wire \ces_1_3_io_ins_left[25] ;
 wire \ces_1_3_io_ins_left[26] ;
 wire \ces_1_3_io_ins_left[27] ;
 wire \ces_1_3_io_ins_left[28] ;
 wire \ces_1_3_io_ins_left[29] ;
 wire \ces_1_3_io_ins_left[2] ;
 wire \ces_1_3_io_ins_left[30] ;
 wire \ces_1_3_io_ins_left[31] ;
 wire \ces_1_3_io_ins_left[32] ;
 wire \ces_1_3_io_ins_left[33] ;
 wire \ces_1_3_io_ins_left[34] ;
 wire \ces_1_3_io_ins_left[35] ;
 wire \ces_1_3_io_ins_left[36] ;
 wire \ces_1_3_io_ins_left[37] ;
 wire \ces_1_3_io_ins_left[38] ;
 wire \ces_1_3_io_ins_left[39] ;
 wire \ces_1_3_io_ins_left[3] ;
 wire \ces_1_3_io_ins_left[40] ;
 wire \ces_1_3_io_ins_left[41] ;
 wire \ces_1_3_io_ins_left[42] ;
 wire \ces_1_3_io_ins_left[43] ;
 wire \ces_1_3_io_ins_left[44] ;
 wire \ces_1_3_io_ins_left[45] ;
 wire \ces_1_3_io_ins_left[46] ;
 wire \ces_1_3_io_ins_left[47] ;
 wire \ces_1_3_io_ins_left[48] ;
 wire \ces_1_3_io_ins_left[49] ;
 wire \ces_1_3_io_ins_left[4] ;
 wire \ces_1_3_io_ins_left[50] ;
 wire \ces_1_3_io_ins_left[51] ;
 wire \ces_1_3_io_ins_left[52] ;
 wire \ces_1_3_io_ins_left[53] ;
 wire \ces_1_3_io_ins_left[54] ;
 wire \ces_1_3_io_ins_left[55] ;
 wire \ces_1_3_io_ins_left[56] ;
 wire \ces_1_3_io_ins_left[57] ;
 wire \ces_1_3_io_ins_left[58] ;
 wire \ces_1_3_io_ins_left[59] ;
 wire \ces_1_3_io_ins_left[5] ;
 wire \ces_1_3_io_ins_left[60] ;
 wire \ces_1_3_io_ins_left[61] ;
 wire \ces_1_3_io_ins_left[62] ;
 wire \ces_1_3_io_ins_left[63] ;
 wire \ces_1_3_io_ins_left[6] ;
 wire \ces_1_3_io_ins_left[7] ;
 wire \ces_1_3_io_ins_left[8] ;
 wire \ces_1_3_io_ins_left[9] ;
 wire ces_1_3_io_lsbOuts_0;
 wire ces_1_3_io_lsbOuts_1;
 wire ces_1_3_io_lsbOuts_2;
 wire ces_1_3_io_lsbOuts_3;
 wire ces_1_3_io_lsbOuts_4;
 wire ces_1_3_io_lsbOuts_5;
 wire ces_1_3_io_lsbOuts_6;
 wire ces_1_3_io_lsbOuts_7;
 wire \ces_1_3_io_outs_right[0] ;
 wire \ces_1_3_io_outs_right[10] ;
 wire \ces_1_3_io_outs_right[11] ;
 wire \ces_1_3_io_outs_right[12] ;
 wire \ces_1_3_io_outs_right[13] ;
 wire \ces_1_3_io_outs_right[14] ;
 wire \ces_1_3_io_outs_right[15] ;
 wire \ces_1_3_io_outs_right[16] ;
 wire \ces_1_3_io_outs_right[17] ;
 wire \ces_1_3_io_outs_right[18] ;
 wire \ces_1_3_io_outs_right[19] ;
 wire \ces_1_3_io_outs_right[1] ;
 wire \ces_1_3_io_outs_right[20] ;
 wire \ces_1_3_io_outs_right[21] ;
 wire \ces_1_3_io_outs_right[22] ;
 wire \ces_1_3_io_outs_right[23] ;
 wire \ces_1_3_io_outs_right[24] ;
 wire \ces_1_3_io_outs_right[25] ;
 wire \ces_1_3_io_outs_right[26] ;
 wire \ces_1_3_io_outs_right[27] ;
 wire \ces_1_3_io_outs_right[28] ;
 wire \ces_1_3_io_outs_right[29] ;
 wire \ces_1_3_io_outs_right[2] ;
 wire \ces_1_3_io_outs_right[30] ;
 wire \ces_1_3_io_outs_right[31] ;
 wire \ces_1_3_io_outs_right[32] ;
 wire \ces_1_3_io_outs_right[33] ;
 wire \ces_1_3_io_outs_right[34] ;
 wire \ces_1_3_io_outs_right[35] ;
 wire \ces_1_3_io_outs_right[36] ;
 wire \ces_1_3_io_outs_right[37] ;
 wire \ces_1_3_io_outs_right[38] ;
 wire \ces_1_3_io_outs_right[39] ;
 wire \ces_1_3_io_outs_right[3] ;
 wire \ces_1_3_io_outs_right[40] ;
 wire \ces_1_3_io_outs_right[41] ;
 wire \ces_1_3_io_outs_right[42] ;
 wire \ces_1_3_io_outs_right[43] ;
 wire \ces_1_3_io_outs_right[44] ;
 wire \ces_1_3_io_outs_right[45] ;
 wire \ces_1_3_io_outs_right[46] ;
 wire \ces_1_3_io_outs_right[47] ;
 wire \ces_1_3_io_outs_right[48] ;
 wire \ces_1_3_io_outs_right[49] ;
 wire \ces_1_3_io_outs_right[4] ;
 wire \ces_1_3_io_outs_right[50] ;
 wire \ces_1_3_io_outs_right[51] ;
 wire \ces_1_3_io_outs_right[52] ;
 wire \ces_1_3_io_outs_right[53] ;
 wire \ces_1_3_io_outs_right[54] ;
 wire \ces_1_3_io_outs_right[55] ;
 wire \ces_1_3_io_outs_right[56] ;
 wire \ces_1_3_io_outs_right[57] ;
 wire \ces_1_3_io_outs_right[58] ;
 wire \ces_1_3_io_outs_right[59] ;
 wire \ces_1_3_io_outs_right[5] ;
 wire \ces_1_3_io_outs_right[60] ;
 wire \ces_1_3_io_outs_right[61] ;
 wire \ces_1_3_io_outs_right[62] ;
 wire \ces_1_3_io_outs_right[63] ;
 wire \ces_1_3_io_outs_right[6] ;
 wire \ces_1_3_io_outs_right[7] ;
 wire \ces_1_3_io_outs_right[8] ;
 wire \ces_1_3_io_outs_right[9] ;
 wire \ces_1_3_io_outs_up[0] ;
 wire \ces_1_3_io_outs_up[10] ;
 wire \ces_1_3_io_outs_up[11] ;
 wire \ces_1_3_io_outs_up[12] ;
 wire \ces_1_3_io_outs_up[13] ;
 wire \ces_1_3_io_outs_up[14] ;
 wire \ces_1_3_io_outs_up[15] ;
 wire \ces_1_3_io_outs_up[16] ;
 wire \ces_1_3_io_outs_up[17] ;
 wire \ces_1_3_io_outs_up[18] ;
 wire \ces_1_3_io_outs_up[19] ;
 wire \ces_1_3_io_outs_up[1] ;
 wire \ces_1_3_io_outs_up[20] ;
 wire \ces_1_3_io_outs_up[21] ;
 wire \ces_1_3_io_outs_up[22] ;
 wire \ces_1_3_io_outs_up[23] ;
 wire \ces_1_3_io_outs_up[24] ;
 wire \ces_1_3_io_outs_up[25] ;
 wire \ces_1_3_io_outs_up[26] ;
 wire \ces_1_3_io_outs_up[27] ;
 wire \ces_1_3_io_outs_up[28] ;
 wire \ces_1_3_io_outs_up[29] ;
 wire \ces_1_3_io_outs_up[2] ;
 wire \ces_1_3_io_outs_up[30] ;
 wire \ces_1_3_io_outs_up[31] ;
 wire \ces_1_3_io_outs_up[32] ;
 wire \ces_1_3_io_outs_up[33] ;
 wire \ces_1_3_io_outs_up[34] ;
 wire \ces_1_3_io_outs_up[35] ;
 wire \ces_1_3_io_outs_up[36] ;
 wire \ces_1_3_io_outs_up[37] ;
 wire \ces_1_3_io_outs_up[38] ;
 wire \ces_1_3_io_outs_up[39] ;
 wire \ces_1_3_io_outs_up[3] ;
 wire \ces_1_3_io_outs_up[40] ;
 wire \ces_1_3_io_outs_up[41] ;
 wire \ces_1_3_io_outs_up[42] ;
 wire \ces_1_3_io_outs_up[43] ;
 wire \ces_1_3_io_outs_up[44] ;
 wire \ces_1_3_io_outs_up[45] ;
 wire \ces_1_3_io_outs_up[46] ;
 wire \ces_1_3_io_outs_up[47] ;
 wire \ces_1_3_io_outs_up[48] ;
 wire \ces_1_3_io_outs_up[49] ;
 wire \ces_1_3_io_outs_up[4] ;
 wire \ces_1_3_io_outs_up[50] ;
 wire \ces_1_3_io_outs_up[51] ;
 wire \ces_1_3_io_outs_up[52] ;
 wire \ces_1_3_io_outs_up[53] ;
 wire \ces_1_3_io_outs_up[54] ;
 wire \ces_1_3_io_outs_up[55] ;
 wire \ces_1_3_io_outs_up[56] ;
 wire \ces_1_3_io_outs_up[57] ;
 wire \ces_1_3_io_outs_up[58] ;
 wire \ces_1_3_io_outs_up[59] ;
 wire \ces_1_3_io_outs_up[5] ;
 wire \ces_1_3_io_outs_up[60] ;
 wire \ces_1_3_io_outs_up[61] ;
 wire \ces_1_3_io_outs_up[62] ;
 wire \ces_1_3_io_outs_up[63] ;
 wire \ces_1_3_io_outs_up[6] ;
 wire \ces_1_3_io_outs_up[7] ;
 wire \ces_1_3_io_outs_up[8] ;
 wire \ces_1_3_io_outs_up[9] ;
 wire \ces_1_4_io_ins_down[0] ;
 wire \ces_1_4_io_ins_down[10] ;
 wire \ces_1_4_io_ins_down[11] ;
 wire \ces_1_4_io_ins_down[12] ;
 wire \ces_1_4_io_ins_down[13] ;
 wire \ces_1_4_io_ins_down[14] ;
 wire \ces_1_4_io_ins_down[15] ;
 wire \ces_1_4_io_ins_down[16] ;
 wire \ces_1_4_io_ins_down[17] ;
 wire \ces_1_4_io_ins_down[18] ;
 wire \ces_1_4_io_ins_down[19] ;
 wire \ces_1_4_io_ins_down[1] ;
 wire \ces_1_4_io_ins_down[20] ;
 wire \ces_1_4_io_ins_down[21] ;
 wire \ces_1_4_io_ins_down[22] ;
 wire \ces_1_4_io_ins_down[23] ;
 wire \ces_1_4_io_ins_down[24] ;
 wire \ces_1_4_io_ins_down[25] ;
 wire \ces_1_4_io_ins_down[26] ;
 wire \ces_1_4_io_ins_down[27] ;
 wire \ces_1_4_io_ins_down[28] ;
 wire \ces_1_4_io_ins_down[29] ;
 wire \ces_1_4_io_ins_down[2] ;
 wire \ces_1_4_io_ins_down[30] ;
 wire \ces_1_4_io_ins_down[31] ;
 wire \ces_1_4_io_ins_down[32] ;
 wire \ces_1_4_io_ins_down[33] ;
 wire \ces_1_4_io_ins_down[34] ;
 wire \ces_1_4_io_ins_down[35] ;
 wire \ces_1_4_io_ins_down[36] ;
 wire \ces_1_4_io_ins_down[37] ;
 wire \ces_1_4_io_ins_down[38] ;
 wire \ces_1_4_io_ins_down[39] ;
 wire \ces_1_4_io_ins_down[3] ;
 wire \ces_1_4_io_ins_down[40] ;
 wire \ces_1_4_io_ins_down[41] ;
 wire \ces_1_4_io_ins_down[42] ;
 wire \ces_1_4_io_ins_down[43] ;
 wire \ces_1_4_io_ins_down[44] ;
 wire \ces_1_4_io_ins_down[45] ;
 wire \ces_1_4_io_ins_down[46] ;
 wire \ces_1_4_io_ins_down[47] ;
 wire \ces_1_4_io_ins_down[48] ;
 wire \ces_1_4_io_ins_down[49] ;
 wire \ces_1_4_io_ins_down[4] ;
 wire \ces_1_4_io_ins_down[50] ;
 wire \ces_1_4_io_ins_down[51] ;
 wire \ces_1_4_io_ins_down[52] ;
 wire \ces_1_4_io_ins_down[53] ;
 wire \ces_1_4_io_ins_down[54] ;
 wire \ces_1_4_io_ins_down[55] ;
 wire \ces_1_4_io_ins_down[56] ;
 wire \ces_1_4_io_ins_down[57] ;
 wire \ces_1_4_io_ins_down[58] ;
 wire \ces_1_4_io_ins_down[59] ;
 wire \ces_1_4_io_ins_down[5] ;
 wire \ces_1_4_io_ins_down[60] ;
 wire \ces_1_4_io_ins_down[61] ;
 wire \ces_1_4_io_ins_down[62] ;
 wire \ces_1_4_io_ins_down[63] ;
 wire \ces_1_4_io_ins_down[6] ;
 wire \ces_1_4_io_ins_down[7] ;
 wire \ces_1_4_io_ins_down[8] ;
 wire \ces_1_4_io_ins_down[9] ;
 wire \ces_1_4_io_ins_left[0] ;
 wire \ces_1_4_io_ins_left[10] ;
 wire \ces_1_4_io_ins_left[11] ;
 wire \ces_1_4_io_ins_left[12] ;
 wire \ces_1_4_io_ins_left[13] ;
 wire \ces_1_4_io_ins_left[14] ;
 wire \ces_1_4_io_ins_left[15] ;
 wire \ces_1_4_io_ins_left[16] ;
 wire \ces_1_4_io_ins_left[17] ;
 wire \ces_1_4_io_ins_left[18] ;
 wire \ces_1_4_io_ins_left[19] ;
 wire \ces_1_4_io_ins_left[1] ;
 wire \ces_1_4_io_ins_left[20] ;
 wire \ces_1_4_io_ins_left[21] ;
 wire \ces_1_4_io_ins_left[22] ;
 wire \ces_1_4_io_ins_left[23] ;
 wire \ces_1_4_io_ins_left[24] ;
 wire \ces_1_4_io_ins_left[25] ;
 wire \ces_1_4_io_ins_left[26] ;
 wire \ces_1_4_io_ins_left[27] ;
 wire \ces_1_4_io_ins_left[28] ;
 wire \ces_1_4_io_ins_left[29] ;
 wire \ces_1_4_io_ins_left[2] ;
 wire \ces_1_4_io_ins_left[30] ;
 wire \ces_1_4_io_ins_left[31] ;
 wire \ces_1_4_io_ins_left[32] ;
 wire \ces_1_4_io_ins_left[33] ;
 wire \ces_1_4_io_ins_left[34] ;
 wire \ces_1_4_io_ins_left[35] ;
 wire \ces_1_4_io_ins_left[36] ;
 wire \ces_1_4_io_ins_left[37] ;
 wire \ces_1_4_io_ins_left[38] ;
 wire \ces_1_4_io_ins_left[39] ;
 wire \ces_1_4_io_ins_left[3] ;
 wire \ces_1_4_io_ins_left[40] ;
 wire \ces_1_4_io_ins_left[41] ;
 wire \ces_1_4_io_ins_left[42] ;
 wire \ces_1_4_io_ins_left[43] ;
 wire \ces_1_4_io_ins_left[44] ;
 wire \ces_1_4_io_ins_left[45] ;
 wire \ces_1_4_io_ins_left[46] ;
 wire \ces_1_4_io_ins_left[47] ;
 wire \ces_1_4_io_ins_left[48] ;
 wire \ces_1_4_io_ins_left[49] ;
 wire \ces_1_4_io_ins_left[4] ;
 wire \ces_1_4_io_ins_left[50] ;
 wire \ces_1_4_io_ins_left[51] ;
 wire \ces_1_4_io_ins_left[52] ;
 wire \ces_1_4_io_ins_left[53] ;
 wire \ces_1_4_io_ins_left[54] ;
 wire \ces_1_4_io_ins_left[55] ;
 wire \ces_1_4_io_ins_left[56] ;
 wire \ces_1_4_io_ins_left[57] ;
 wire \ces_1_4_io_ins_left[58] ;
 wire \ces_1_4_io_ins_left[59] ;
 wire \ces_1_4_io_ins_left[5] ;
 wire \ces_1_4_io_ins_left[60] ;
 wire \ces_1_4_io_ins_left[61] ;
 wire \ces_1_4_io_ins_left[62] ;
 wire \ces_1_4_io_ins_left[63] ;
 wire \ces_1_4_io_ins_left[6] ;
 wire \ces_1_4_io_ins_left[7] ;
 wire \ces_1_4_io_ins_left[8] ;
 wire \ces_1_4_io_ins_left[9] ;
 wire ces_1_4_io_lsbOuts_0;
 wire ces_1_4_io_lsbOuts_1;
 wire ces_1_4_io_lsbOuts_2;
 wire ces_1_4_io_lsbOuts_3;
 wire ces_1_4_io_lsbOuts_4;
 wire ces_1_4_io_lsbOuts_5;
 wire ces_1_4_io_lsbOuts_6;
 wire ces_1_4_io_lsbOuts_7;
 wire \ces_1_4_io_outs_right[0] ;
 wire \ces_1_4_io_outs_right[10] ;
 wire \ces_1_4_io_outs_right[11] ;
 wire \ces_1_4_io_outs_right[12] ;
 wire \ces_1_4_io_outs_right[13] ;
 wire \ces_1_4_io_outs_right[14] ;
 wire \ces_1_4_io_outs_right[15] ;
 wire \ces_1_4_io_outs_right[16] ;
 wire \ces_1_4_io_outs_right[17] ;
 wire \ces_1_4_io_outs_right[18] ;
 wire \ces_1_4_io_outs_right[19] ;
 wire \ces_1_4_io_outs_right[1] ;
 wire \ces_1_4_io_outs_right[20] ;
 wire \ces_1_4_io_outs_right[21] ;
 wire \ces_1_4_io_outs_right[22] ;
 wire \ces_1_4_io_outs_right[23] ;
 wire \ces_1_4_io_outs_right[24] ;
 wire \ces_1_4_io_outs_right[25] ;
 wire \ces_1_4_io_outs_right[26] ;
 wire \ces_1_4_io_outs_right[27] ;
 wire \ces_1_4_io_outs_right[28] ;
 wire \ces_1_4_io_outs_right[29] ;
 wire \ces_1_4_io_outs_right[2] ;
 wire \ces_1_4_io_outs_right[30] ;
 wire \ces_1_4_io_outs_right[31] ;
 wire \ces_1_4_io_outs_right[32] ;
 wire \ces_1_4_io_outs_right[33] ;
 wire \ces_1_4_io_outs_right[34] ;
 wire \ces_1_4_io_outs_right[35] ;
 wire \ces_1_4_io_outs_right[36] ;
 wire \ces_1_4_io_outs_right[37] ;
 wire \ces_1_4_io_outs_right[38] ;
 wire \ces_1_4_io_outs_right[39] ;
 wire \ces_1_4_io_outs_right[3] ;
 wire \ces_1_4_io_outs_right[40] ;
 wire \ces_1_4_io_outs_right[41] ;
 wire \ces_1_4_io_outs_right[42] ;
 wire \ces_1_4_io_outs_right[43] ;
 wire \ces_1_4_io_outs_right[44] ;
 wire \ces_1_4_io_outs_right[45] ;
 wire \ces_1_4_io_outs_right[46] ;
 wire \ces_1_4_io_outs_right[47] ;
 wire \ces_1_4_io_outs_right[48] ;
 wire \ces_1_4_io_outs_right[49] ;
 wire \ces_1_4_io_outs_right[4] ;
 wire \ces_1_4_io_outs_right[50] ;
 wire \ces_1_4_io_outs_right[51] ;
 wire \ces_1_4_io_outs_right[52] ;
 wire \ces_1_4_io_outs_right[53] ;
 wire \ces_1_4_io_outs_right[54] ;
 wire \ces_1_4_io_outs_right[55] ;
 wire \ces_1_4_io_outs_right[56] ;
 wire \ces_1_4_io_outs_right[57] ;
 wire \ces_1_4_io_outs_right[58] ;
 wire \ces_1_4_io_outs_right[59] ;
 wire \ces_1_4_io_outs_right[5] ;
 wire \ces_1_4_io_outs_right[60] ;
 wire \ces_1_4_io_outs_right[61] ;
 wire \ces_1_4_io_outs_right[62] ;
 wire \ces_1_4_io_outs_right[63] ;
 wire \ces_1_4_io_outs_right[6] ;
 wire \ces_1_4_io_outs_right[7] ;
 wire \ces_1_4_io_outs_right[8] ;
 wire \ces_1_4_io_outs_right[9] ;
 wire \ces_1_4_io_outs_up[0] ;
 wire \ces_1_4_io_outs_up[10] ;
 wire \ces_1_4_io_outs_up[11] ;
 wire \ces_1_4_io_outs_up[12] ;
 wire \ces_1_4_io_outs_up[13] ;
 wire \ces_1_4_io_outs_up[14] ;
 wire \ces_1_4_io_outs_up[15] ;
 wire \ces_1_4_io_outs_up[16] ;
 wire \ces_1_4_io_outs_up[17] ;
 wire \ces_1_4_io_outs_up[18] ;
 wire \ces_1_4_io_outs_up[19] ;
 wire \ces_1_4_io_outs_up[1] ;
 wire \ces_1_4_io_outs_up[20] ;
 wire \ces_1_4_io_outs_up[21] ;
 wire \ces_1_4_io_outs_up[22] ;
 wire \ces_1_4_io_outs_up[23] ;
 wire \ces_1_4_io_outs_up[24] ;
 wire \ces_1_4_io_outs_up[25] ;
 wire \ces_1_4_io_outs_up[26] ;
 wire \ces_1_4_io_outs_up[27] ;
 wire \ces_1_4_io_outs_up[28] ;
 wire \ces_1_4_io_outs_up[29] ;
 wire \ces_1_4_io_outs_up[2] ;
 wire \ces_1_4_io_outs_up[30] ;
 wire \ces_1_4_io_outs_up[31] ;
 wire \ces_1_4_io_outs_up[32] ;
 wire \ces_1_4_io_outs_up[33] ;
 wire \ces_1_4_io_outs_up[34] ;
 wire \ces_1_4_io_outs_up[35] ;
 wire \ces_1_4_io_outs_up[36] ;
 wire \ces_1_4_io_outs_up[37] ;
 wire \ces_1_4_io_outs_up[38] ;
 wire \ces_1_4_io_outs_up[39] ;
 wire \ces_1_4_io_outs_up[3] ;
 wire \ces_1_4_io_outs_up[40] ;
 wire \ces_1_4_io_outs_up[41] ;
 wire \ces_1_4_io_outs_up[42] ;
 wire \ces_1_4_io_outs_up[43] ;
 wire \ces_1_4_io_outs_up[44] ;
 wire \ces_1_4_io_outs_up[45] ;
 wire \ces_1_4_io_outs_up[46] ;
 wire \ces_1_4_io_outs_up[47] ;
 wire \ces_1_4_io_outs_up[48] ;
 wire \ces_1_4_io_outs_up[49] ;
 wire \ces_1_4_io_outs_up[4] ;
 wire \ces_1_4_io_outs_up[50] ;
 wire \ces_1_4_io_outs_up[51] ;
 wire \ces_1_4_io_outs_up[52] ;
 wire \ces_1_4_io_outs_up[53] ;
 wire \ces_1_4_io_outs_up[54] ;
 wire \ces_1_4_io_outs_up[55] ;
 wire \ces_1_4_io_outs_up[56] ;
 wire \ces_1_4_io_outs_up[57] ;
 wire \ces_1_4_io_outs_up[58] ;
 wire \ces_1_4_io_outs_up[59] ;
 wire \ces_1_4_io_outs_up[5] ;
 wire \ces_1_4_io_outs_up[60] ;
 wire \ces_1_4_io_outs_up[61] ;
 wire \ces_1_4_io_outs_up[62] ;
 wire \ces_1_4_io_outs_up[63] ;
 wire \ces_1_4_io_outs_up[6] ;
 wire \ces_1_4_io_outs_up[7] ;
 wire \ces_1_4_io_outs_up[8] ;
 wire \ces_1_4_io_outs_up[9] ;
 wire \ces_1_5_io_ins_down[0] ;
 wire \ces_1_5_io_ins_down[10] ;
 wire \ces_1_5_io_ins_down[11] ;
 wire \ces_1_5_io_ins_down[12] ;
 wire \ces_1_5_io_ins_down[13] ;
 wire \ces_1_5_io_ins_down[14] ;
 wire \ces_1_5_io_ins_down[15] ;
 wire \ces_1_5_io_ins_down[16] ;
 wire \ces_1_5_io_ins_down[17] ;
 wire \ces_1_5_io_ins_down[18] ;
 wire \ces_1_5_io_ins_down[19] ;
 wire \ces_1_5_io_ins_down[1] ;
 wire \ces_1_5_io_ins_down[20] ;
 wire \ces_1_5_io_ins_down[21] ;
 wire \ces_1_5_io_ins_down[22] ;
 wire \ces_1_5_io_ins_down[23] ;
 wire \ces_1_5_io_ins_down[24] ;
 wire \ces_1_5_io_ins_down[25] ;
 wire \ces_1_5_io_ins_down[26] ;
 wire \ces_1_5_io_ins_down[27] ;
 wire \ces_1_5_io_ins_down[28] ;
 wire \ces_1_5_io_ins_down[29] ;
 wire \ces_1_5_io_ins_down[2] ;
 wire \ces_1_5_io_ins_down[30] ;
 wire \ces_1_5_io_ins_down[31] ;
 wire \ces_1_5_io_ins_down[32] ;
 wire \ces_1_5_io_ins_down[33] ;
 wire \ces_1_5_io_ins_down[34] ;
 wire \ces_1_5_io_ins_down[35] ;
 wire \ces_1_5_io_ins_down[36] ;
 wire \ces_1_5_io_ins_down[37] ;
 wire \ces_1_5_io_ins_down[38] ;
 wire \ces_1_5_io_ins_down[39] ;
 wire \ces_1_5_io_ins_down[3] ;
 wire \ces_1_5_io_ins_down[40] ;
 wire \ces_1_5_io_ins_down[41] ;
 wire \ces_1_5_io_ins_down[42] ;
 wire \ces_1_5_io_ins_down[43] ;
 wire \ces_1_5_io_ins_down[44] ;
 wire \ces_1_5_io_ins_down[45] ;
 wire \ces_1_5_io_ins_down[46] ;
 wire \ces_1_5_io_ins_down[47] ;
 wire \ces_1_5_io_ins_down[48] ;
 wire \ces_1_5_io_ins_down[49] ;
 wire \ces_1_5_io_ins_down[4] ;
 wire \ces_1_5_io_ins_down[50] ;
 wire \ces_1_5_io_ins_down[51] ;
 wire \ces_1_5_io_ins_down[52] ;
 wire \ces_1_5_io_ins_down[53] ;
 wire \ces_1_5_io_ins_down[54] ;
 wire \ces_1_5_io_ins_down[55] ;
 wire \ces_1_5_io_ins_down[56] ;
 wire \ces_1_5_io_ins_down[57] ;
 wire \ces_1_5_io_ins_down[58] ;
 wire \ces_1_5_io_ins_down[59] ;
 wire \ces_1_5_io_ins_down[5] ;
 wire \ces_1_5_io_ins_down[60] ;
 wire \ces_1_5_io_ins_down[61] ;
 wire \ces_1_5_io_ins_down[62] ;
 wire \ces_1_5_io_ins_down[63] ;
 wire \ces_1_5_io_ins_down[6] ;
 wire \ces_1_5_io_ins_down[7] ;
 wire \ces_1_5_io_ins_down[8] ;
 wire \ces_1_5_io_ins_down[9] ;
 wire \ces_1_5_io_ins_left[0] ;
 wire \ces_1_5_io_ins_left[10] ;
 wire \ces_1_5_io_ins_left[11] ;
 wire \ces_1_5_io_ins_left[12] ;
 wire \ces_1_5_io_ins_left[13] ;
 wire \ces_1_5_io_ins_left[14] ;
 wire \ces_1_5_io_ins_left[15] ;
 wire \ces_1_5_io_ins_left[16] ;
 wire \ces_1_5_io_ins_left[17] ;
 wire \ces_1_5_io_ins_left[18] ;
 wire \ces_1_5_io_ins_left[19] ;
 wire \ces_1_5_io_ins_left[1] ;
 wire \ces_1_5_io_ins_left[20] ;
 wire \ces_1_5_io_ins_left[21] ;
 wire \ces_1_5_io_ins_left[22] ;
 wire \ces_1_5_io_ins_left[23] ;
 wire \ces_1_5_io_ins_left[24] ;
 wire \ces_1_5_io_ins_left[25] ;
 wire \ces_1_5_io_ins_left[26] ;
 wire \ces_1_5_io_ins_left[27] ;
 wire \ces_1_5_io_ins_left[28] ;
 wire \ces_1_5_io_ins_left[29] ;
 wire \ces_1_5_io_ins_left[2] ;
 wire \ces_1_5_io_ins_left[30] ;
 wire \ces_1_5_io_ins_left[31] ;
 wire \ces_1_5_io_ins_left[32] ;
 wire \ces_1_5_io_ins_left[33] ;
 wire \ces_1_5_io_ins_left[34] ;
 wire \ces_1_5_io_ins_left[35] ;
 wire \ces_1_5_io_ins_left[36] ;
 wire \ces_1_5_io_ins_left[37] ;
 wire \ces_1_5_io_ins_left[38] ;
 wire \ces_1_5_io_ins_left[39] ;
 wire \ces_1_5_io_ins_left[3] ;
 wire \ces_1_5_io_ins_left[40] ;
 wire \ces_1_5_io_ins_left[41] ;
 wire \ces_1_5_io_ins_left[42] ;
 wire \ces_1_5_io_ins_left[43] ;
 wire \ces_1_5_io_ins_left[44] ;
 wire \ces_1_5_io_ins_left[45] ;
 wire \ces_1_5_io_ins_left[46] ;
 wire \ces_1_5_io_ins_left[47] ;
 wire \ces_1_5_io_ins_left[48] ;
 wire \ces_1_5_io_ins_left[49] ;
 wire \ces_1_5_io_ins_left[4] ;
 wire \ces_1_5_io_ins_left[50] ;
 wire \ces_1_5_io_ins_left[51] ;
 wire \ces_1_5_io_ins_left[52] ;
 wire \ces_1_5_io_ins_left[53] ;
 wire \ces_1_5_io_ins_left[54] ;
 wire \ces_1_5_io_ins_left[55] ;
 wire \ces_1_5_io_ins_left[56] ;
 wire \ces_1_5_io_ins_left[57] ;
 wire \ces_1_5_io_ins_left[58] ;
 wire \ces_1_5_io_ins_left[59] ;
 wire \ces_1_5_io_ins_left[5] ;
 wire \ces_1_5_io_ins_left[60] ;
 wire \ces_1_5_io_ins_left[61] ;
 wire \ces_1_5_io_ins_left[62] ;
 wire \ces_1_5_io_ins_left[63] ;
 wire \ces_1_5_io_ins_left[6] ;
 wire \ces_1_5_io_ins_left[7] ;
 wire \ces_1_5_io_ins_left[8] ;
 wire \ces_1_5_io_ins_left[9] ;
 wire ces_1_5_io_lsbOuts_0;
 wire ces_1_5_io_lsbOuts_1;
 wire ces_1_5_io_lsbOuts_2;
 wire ces_1_5_io_lsbOuts_3;
 wire ces_1_5_io_lsbOuts_4;
 wire ces_1_5_io_lsbOuts_5;
 wire ces_1_5_io_lsbOuts_6;
 wire ces_1_5_io_lsbOuts_7;
 wire \ces_1_5_io_outs_right[0] ;
 wire \ces_1_5_io_outs_right[10] ;
 wire \ces_1_5_io_outs_right[11] ;
 wire \ces_1_5_io_outs_right[12] ;
 wire \ces_1_5_io_outs_right[13] ;
 wire \ces_1_5_io_outs_right[14] ;
 wire \ces_1_5_io_outs_right[15] ;
 wire \ces_1_5_io_outs_right[16] ;
 wire \ces_1_5_io_outs_right[17] ;
 wire \ces_1_5_io_outs_right[18] ;
 wire \ces_1_5_io_outs_right[19] ;
 wire \ces_1_5_io_outs_right[1] ;
 wire \ces_1_5_io_outs_right[20] ;
 wire \ces_1_5_io_outs_right[21] ;
 wire \ces_1_5_io_outs_right[22] ;
 wire \ces_1_5_io_outs_right[23] ;
 wire \ces_1_5_io_outs_right[24] ;
 wire \ces_1_5_io_outs_right[25] ;
 wire \ces_1_5_io_outs_right[26] ;
 wire \ces_1_5_io_outs_right[27] ;
 wire \ces_1_5_io_outs_right[28] ;
 wire \ces_1_5_io_outs_right[29] ;
 wire \ces_1_5_io_outs_right[2] ;
 wire \ces_1_5_io_outs_right[30] ;
 wire \ces_1_5_io_outs_right[31] ;
 wire \ces_1_5_io_outs_right[32] ;
 wire \ces_1_5_io_outs_right[33] ;
 wire \ces_1_5_io_outs_right[34] ;
 wire \ces_1_5_io_outs_right[35] ;
 wire \ces_1_5_io_outs_right[36] ;
 wire \ces_1_5_io_outs_right[37] ;
 wire \ces_1_5_io_outs_right[38] ;
 wire \ces_1_5_io_outs_right[39] ;
 wire \ces_1_5_io_outs_right[3] ;
 wire \ces_1_5_io_outs_right[40] ;
 wire \ces_1_5_io_outs_right[41] ;
 wire \ces_1_5_io_outs_right[42] ;
 wire \ces_1_5_io_outs_right[43] ;
 wire \ces_1_5_io_outs_right[44] ;
 wire \ces_1_5_io_outs_right[45] ;
 wire \ces_1_5_io_outs_right[46] ;
 wire \ces_1_5_io_outs_right[47] ;
 wire \ces_1_5_io_outs_right[48] ;
 wire \ces_1_5_io_outs_right[49] ;
 wire \ces_1_5_io_outs_right[4] ;
 wire \ces_1_5_io_outs_right[50] ;
 wire \ces_1_5_io_outs_right[51] ;
 wire \ces_1_5_io_outs_right[52] ;
 wire \ces_1_5_io_outs_right[53] ;
 wire \ces_1_5_io_outs_right[54] ;
 wire \ces_1_5_io_outs_right[55] ;
 wire \ces_1_5_io_outs_right[56] ;
 wire \ces_1_5_io_outs_right[57] ;
 wire \ces_1_5_io_outs_right[58] ;
 wire \ces_1_5_io_outs_right[59] ;
 wire \ces_1_5_io_outs_right[5] ;
 wire \ces_1_5_io_outs_right[60] ;
 wire \ces_1_5_io_outs_right[61] ;
 wire \ces_1_5_io_outs_right[62] ;
 wire \ces_1_5_io_outs_right[63] ;
 wire \ces_1_5_io_outs_right[6] ;
 wire \ces_1_5_io_outs_right[7] ;
 wire \ces_1_5_io_outs_right[8] ;
 wire \ces_1_5_io_outs_right[9] ;
 wire \ces_1_5_io_outs_up[0] ;
 wire \ces_1_5_io_outs_up[10] ;
 wire \ces_1_5_io_outs_up[11] ;
 wire \ces_1_5_io_outs_up[12] ;
 wire \ces_1_5_io_outs_up[13] ;
 wire \ces_1_5_io_outs_up[14] ;
 wire \ces_1_5_io_outs_up[15] ;
 wire \ces_1_5_io_outs_up[16] ;
 wire \ces_1_5_io_outs_up[17] ;
 wire \ces_1_5_io_outs_up[18] ;
 wire \ces_1_5_io_outs_up[19] ;
 wire \ces_1_5_io_outs_up[1] ;
 wire \ces_1_5_io_outs_up[20] ;
 wire \ces_1_5_io_outs_up[21] ;
 wire \ces_1_5_io_outs_up[22] ;
 wire \ces_1_5_io_outs_up[23] ;
 wire \ces_1_5_io_outs_up[24] ;
 wire \ces_1_5_io_outs_up[25] ;
 wire \ces_1_5_io_outs_up[26] ;
 wire \ces_1_5_io_outs_up[27] ;
 wire \ces_1_5_io_outs_up[28] ;
 wire \ces_1_5_io_outs_up[29] ;
 wire \ces_1_5_io_outs_up[2] ;
 wire \ces_1_5_io_outs_up[30] ;
 wire \ces_1_5_io_outs_up[31] ;
 wire \ces_1_5_io_outs_up[32] ;
 wire \ces_1_5_io_outs_up[33] ;
 wire \ces_1_5_io_outs_up[34] ;
 wire \ces_1_5_io_outs_up[35] ;
 wire \ces_1_5_io_outs_up[36] ;
 wire \ces_1_5_io_outs_up[37] ;
 wire \ces_1_5_io_outs_up[38] ;
 wire \ces_1_5_io_outs_up[39] ;
 wire \ces_1_5_io_outs_up[3] ;
 wire \ces_1_5_io_outs_up[40] ;
 wire \ces_1_5_io_outs_up[41] ;
 wire \ces_1_5_io_outs_up[42] ;
 wire \ces_1_5_io_outs_up[43] ;
 wire \ces_1_5_io_outs_up[44] ;
 wire \ces_1_5_io_outs_up[45] ;
 wire \ces_1_5_io_outs_up[46] ;
 wire \ces_1_5_io_outs_up[47] ;
 wire \ces_1_5_io_outs_up[48] ;
 wire \ces_1_5_io_outs_up[49] ;
 wire \ces_1_5_io_outs_up[4] ;
 wire \ces_1_5_io_outs_up[50] ;
 wire \ces_1_5_io_outs_up[51] ;
 wire \ces_1_5_io_outs_up[52] ;
 wire \ces_1_5_io_outs_up[53] ;
 wire \ces_1_5_io_outs_up[54] ;
 wire \ces_1_5_io_outs_up[55] ;
 wire \ces_1_5_io_outs_up[56] ;
 wire \ces_1_5_io_outs_up[57] ;
 wire \ces_1_5_io_outs_up[58] ;
 wire \ces_1_5_io_outs_up[59] ;
 wire \ces_1_5_io_outs_up[5] ;
 wire \ces_1_5_io_outs_up[60] ;
 wire \ces_1_5_io_outs_up[61] ;
 wire \ces_1_5_io_outs_up[62] ;
 wire \ces_1_5_io_outs_up[63] ;
 wire \ces_1_5_io_outs_up[6] ;
 wire \ces_1_5_io_outs_up[7] ;
 wire \ces_1_5_io_outs_up[8] ;
 wire \ces_1_5_io_outs_up[9] ;
 wire \ces_1_6_io_ins_down[0] ;
 wire \ces_1_6_io_ins_down[10] ;
 wire \ces_1_6_io_ins_down[11] ;
 wire \ces_1_6_io_ins_down[12] ;
 wire \ces_1_6_io_ins_down[13] ;
 wire \ces_1_6_io_ins_down[14] ;
 wire \ces_1_6_io_ins_down[15] ;
 wire \ces_1_6_io_ins_down[16] ;
 wire \ces_1_6_io_ins_down[17] ;
 wire \ces_1_6_io_ins_down[18] ;
 wire \ces_1_6_io_ins_down[19] ;
 wire \ces_1_6_io_ins_down[1] ;
 wire \ces_1_6_io_ins_down[20] ;
 wire \ces_1_6_io_ins_down[21] ;
 wire \ces_1_6_io_ins_down[22] ;
 wire \ces_1_6_io_ins_down[23] ;
 wire \ces_1_6_io_ins_down[24] ;
 wire \ces_1_6_io_ins_down[25] ;
 wire \ces_1_6_io_ins_down[26] ;
 wire \ces_1_6_io_ins_down[27] ;
 wire \ces_1_6_io_ins_down[28] ;
 wire \ces_1_6_io_ins_down[29] ;
 wire \ces_1_6_io_ins_down[2] ;
 wire \ces_1_6_io_ins_down[30] ;
 wire \ces_1_6_io_ins_down[31] ;
 wire \ces_1_6_io_ins_down[32] ;
 wire \ces_1_6_io_ins_down[33] ;
 wire \ces_1_6_io_ins_down[34] ;
 wire \ces_1_6_io_ins_down[35] ;
 wire \ces_1_6_io_ins_down[36] ;
 wire \ces_1_6_io_ins_down[37] ;
 wire \ces_1_6_io_ins_down[38] ;
 wire \ces_1_6_io_ins_down[39] ;
 wire \ces_1_6_io_ins_down[3] ;
 wire \ces_1_6_io_ins_down[40] ;
 wire \ces_1_6_io_ins_down[41] ;
 wire \ces_1_6_io_ins_down[42] ;
 wire \ces_1_6_io_ins_down[43] ;
 wire \ces_1_6_io_ins_down[44] ;
 wire \ces_1_6_io_ins_down[45] ;
 wire \ces_1_6_io_ins_down[46] ;
 wire \ces_1_6_io_ins_down[47] ;
 wire \ces_1_6_io_ins_down[48] ;
 wire \ces_1_6_io_ins_down[49] ;
 wire \ces_1_6_io_ins_down[4] ;
 wire \ces_1_6_io_ins_down[50] ;
 wire \ces_1_6_io_ins_down[51] ;
 wire \ces_1_6_io_ins_down[52] ;
 wire \ces_1_6_io_ins_down[53] ;
 wire \ces_1_6_io_ins_down[54] ;
 wire \ces_1_6_io_ins_down[55] ;
 wire \ces_1_6_io_ins_down[56] ;
 wire \ces_1_6_io_ins_down[57] ;
 wire \ces_1_6_io_ins_down[58] ;
 wire \ces_1_6_io_ins_down[59] ;
 wire \ces_1_6_io_ins_down[5] ;
 wire \ces_1_6_io_ins_down[60] ;
 wire \ces_1_6_io_ins_down[61] ;
 wire \ces_1_6_io_ins_down[62] ;
 wire \ces_1_6_io_ins_down[63] ;
 wire \ces_1_6_io_ins_down[6] ;
 wire \ces_1_6_io_ins_down[7] ;
 wire \ces_1_6_io_ins_down[8] ;
 wire \ces_1_6_io_ins_down[9] ;
 wire \ces_1_6_io_ins_left[0] ;
 wire \ces_1_6_io_ins_left[10] ;
 wire \ces_1_6_io_ins_left[11] ;
 wire \ces_1_6_io_ins_left[12] ;
 wire \ces_1_6_io_ins_left[13] ;
 wire \ces_1_6_io_ins_left[14] ;
 wire \ces_1_6_io_ins_left[15] ;
 wire \ces_1_6_io_ins_left[16] ;
 wire \ces_1_6_io_ins_left[17] ;
 wire \ces_1_6_io_ins_left[18] ;
 wire \ces_1_6_io_ins_left[19] ;
 wire \ces_1_6_io_ins_left[1] ;
 wire \ces_1_6_io_ins_left[20] ;
 wire \ces_1_6_io_ins_left[21] ;
 wire \ces_1_6_io_ins_left[22] ;
 wire \ces_1_6_io_ins_left[23] ;
 wire \ces_1_6_io_ins_left[24] ;
 wire \ces_1_6_io_ins_left[25] ;
 wire \ces_1_6_io_ins_left[26] ;
 wire \ces_1_6_io_ins_left[27] ;
 wire \ces_1_6_io_ins_left[28] ;
 wire \ces_1_6_io_ins_left[29] ;
 wire \ces_1_6_io_ins_left[2] ;
 wire \ces_1_6_io_ins_left[30] ;
 wire \ces_1_6_io_ins_left[31] ;
 wire \ces_1_6_io_ins_left[32] ;
 wire \ces_1_6_io_ins_left[33] ;
 wire \ces_1_6_io_ins_left[34] ;
 wire \ces_1_6_io_ins_left[35] ;
 wire \ces_1_6_io_ins_left[36] ;
 wire \ces_1_6_io_ins_left[37] ;
 wire \ces_1_6_io_ins_left[38] ;
 wire \ces_1_6_io_ins_left[39] ;
 wire \ces_1_6_io_ins_left[3] ;
 wire \ces_1_6_io_ins_left[40] ;
 wire \ces_1_6_io_ins_left[41] ;
 wire \ces_1_6_io_ins_left[42] ;
 wire \ces_1_6_io_ins_left[43] ;
 wire \ces_1_6_io_ins_left[44] ;
 wire \ces_1_6_io_ins_left[45] ;
 wire \ces_1_6_io_ins_left[46] ;
 wire \ces_1_6_io_ins_left[47] ;
 wire \ces_1_6_io_ins_left[48] ;
 wire \ces_1_6_io_ins_left[49] ;
 wire \ces_1_6_io_ins_left[4] ;
 wire \ces_1_6_io_ins_left[50] ;
 wire \ces_1_6_io_ins_left[51] ;
 wire \ces_1_6_io_ins_left[52] ;
 wire \ces_1_6_io_ins_left[53] ;
 wire \ces_1_6_io_ins_left[54] ;
 wire \ces_1_6_io_ins_left[55] ;
 wire \ces_1_6_io_ins_left[56] ;
 wire \ces_1_6_io_ins_left[57] ;
 wire \ces_1_6_io_ins_left[58] ;
 wire \ces_1_6_io_ins_left[59] ;
 wire \ces_1_6_io_ins_left[5] ;
 wire \ces_1_6_io_ins_left[60] ;
 wire \ces_1_6_io_ins_left[61] ;
 wire \ces_1_6_io_ins_left[62] ;
 wire \ces_1_6_io_ins_left[63] ;
 wire \ces_1_6_io_ins_left[6] ;
 wire \ces_1_6_io_ins_left[7] ;
 wire \ces_1_6_io_ins_left[8] ;
 wire \ces_1_6_io_ins_left[9] ;
 wire ces_1_6_io_lsbOuts_0;
 wire ces_1_6_io_lsbOuts_1;
 wire ces_1_6_io_lsbOuts_2;
 wire ces_1_6_io_lsbOuts_3;
 wire ces_1_6_io_lsbOuts_4;
 wire ces_1_6_io_lsbOuts_5;
 wire ces_1_6_io_lsbOuts_6;
 wire ces_1_6_io_lsbOuts_7;
 wire \ces_1_6_io_outs_right[0] ;
 wire \ces_1_6_io_outs_right[10] ;
 wire \ces_1_6_io_outs_right[11] ;
 wire \ces_1_6_io_outs_right[12] ;
 wire \ces_1_6_io_outs_right[13] ;
 wire \ces_1_6_io_outs_right[14] ;
 wire \ces_1_6_io_outs_right[15] ;
 wire \ces_1_6_io_outs_right[16] ;
 wire \ces_1_6_io_outs_right[17] ;
 wire \ces_1_6_io_outs_right[18] ;
 wire \ces_1_6_io_outs_right[19] ;
 wire \ces_1_6_io_outs_right[1] ;
 wire \ces_1_6_io_outs_right[20] ;
 wire \ces_1_6_io_outs_right[21] ;
 wire \ces_1_6_io_outs_right[22] ;
 wire \ces_1_6_io_outs_right[23] ;
 wire \ces_1_6_io_outs_right[24] ;
 wire \ces_1_6_io_outs_right[25] ;
 wire \ces_1_6_io_outs_right[26] ;
 wire \ces_1_6_io_outs_right[27] ;
 wire \ces_1_6_io_outs_right[28] ;
 wire \ces_1_6_io_outs_right[29] ;
 wire \ces_1_6_io_outs_right[2] ;
 wire \ces_1_6_io_outs_right[30] ;
 wire \ces_1_6_io_outs_right[31] ;
 wire \ces_1_6_io_outs_right[32] ;
 wire \ces_1_6_io_outs_right[33] ;
 wire \ces_1_6_io_outs_right[34] ;
 wire \ces_1_6_io_outs_right[35] ;
 wire \ces_1_6_io_outs_right[36] ;
 wire \ces_1_6_io_outs_right[37] ;
 wire \ces_1_6_io_outs_right[38] ;
 wire \ces_1_6_io_outs_right[39] ;
 wire \ces_1_6_io_outs_right[3] ;
 wire \ces_1_6_io_outs_right[40] ;
 wire \ces_1_6_io_outs_right[41] ;
 wire \ces_1_6_io_outs_right[42] ;
 wire \ces_1_6_io_outs_right[43] ;
 wire \ces_1_6_io_outs_right[44] ;
 wire \ces_1_6_io_outs_right[45] ;
 wire \ces_1_6_io_outs_right[46] ;
 wire \ces_1_6_io_outs_right[47] ;
 wire \ces_1_6_io_outs_right[48] ;
 wire \ces_1_6_io_outs_right[49] ;
 wire \ces_1_6_io_outs_right[4] ;
 wire \ces_1_6_io_outs_right[50] ;
 wire \ces_1_6_io_outs_right[51] ;
 wire \ces_1_6_io_outs_right[52] ;
 wire \ces_1_6_io_outs_right[53] ;
 wire \ces_1_6_io_outs_right[54] ;
 wire \ces_1_6_io_outs_right[55] ;
 wire \ces_1_6_io_outs_right[56] ;
 wire \ces_1_6_io_outs_right[57] ;
 wire \ces_1_6_io_outs_right[58] ;
 wire \ces_1_6_io_outs_right[59] ;
 wire \ces_1_6_io_outs_right[5] ;
 wire \ces_1_6_io_outs_right[60] ;
 wire \ces_1_6_io_outs_right[61] ;
 wire \ces_1_6_io_outs_right[62] ;
 wire \ces_1_6_io_outs_right[63] ;
 wire \ces_1_6_io_outs_right[6] ;
 wire \ces_1_6_io_outs_right[7] ;
 wire \ces_1_6_io_outs_right[8] ;
 wire \ces_1_6_io_outs_right[9] ;
 wire \ces_1_6_io_outs_up[0] ;
 wire \ces_1_6_io_outs_up[10] ;
 wire \ces_1_6_io_outs_up[11] ;
 wire \ces_1_6_io_outs_up[12] ;
 wire \ces_1_6_io_outs_up[13] ;
 wire \ces_1_6_io_outs_up[14] ;
 wire \ces_1_6_io_outs_up[15] ;
 wire \ces_1_6_io_outs_up[16] ;
 wire \ces_1_6_io_outs_up[17] ;
 wire \ces_1_6_io_outs_up[18] ;
 wire \ces_1_6_io_outs_up[19] ;
 wire \ces_1_6_io_outs_up[1] ;
 wire \ces_1_6_io_outs_up[20] ;
 wire \ces_1_6_io_outs_up[21] ;
 wire \ces_1_6_io_outs_up[22] ;
 wire \ces_1_6_io_outs_up[23] ;
 wire \ces_1_6_io_outs_up[24] ;
 wire \ces_1_6_io_outs_up[25] ;
 wire \ces_1_6_io_outs_up[26] ;
 wire \ces_1_6_io_outs_up[27] ;
 wire \ces_1_6_io_outs_up[28] ;
 wire \ces_1_6_io_outs_up[29] ;
 wire \ces_1_6_io_outs_up[2] ;
 wire \ces_1_6_io_outs_up[30] ;
 wire \ces_1_6_io_outs_up[31] ;
 wire \ces_1_6_io_outs_up[32] ;
 wire \ces_1_6_io_outs_up[33] ;
 wire \ces_1_6_io_outs_up[34] ;
 wire \ces_1_6_io_outs_up[35] ;
 wire \ces_1_6_io_outs_up[36] ;
 wire \ces_1_6_io_outs_up[37] ;
 wire \ces_1_6_io_outs_up[38] ;
 wire \ces_1_6_io_outs_up[39] ;
 wire \ces_1_6_io_outs_up[3] ;
 wire \ces_1_6_io_outs_up[40] ;
 wire \ces_1_6_io_outs_up[41] ;
 wire \ces_1_6_io_outs_up[42] ;
 wire \ces_1_6_io_outs_up[43] ;
 wire \ces_1_6_io_outs_up[44] ;
 wire \ces_1_6_io_outs_up[45] ;
 wire \ces_1_6_io_outs_up[46] ;
 wire \ces_1_6_io_outs_up[47] ;
 wire \ces_1_6_io_outs_up[48] ;
 wire \ces_1_6_io_outs_up[49] ;
 wire \ces_1_6_io_outs_up[4] ;
 wire \ces_1_6_io_outs_up[50] ;
 wire \ces_1_6_io_outs_up[51] ;
 wire \ces_1_6_io_outs_up[52] ;
 wire \ces_1_6_io_outs_up[53] ;
 wire \ces_1_6_io_outs_up[54] ;
 wire \ces_1_6_io_outs_up[55] ;
 wire \ces_1_6_io_outs_up[56] ;
 wire \ces_1_6_io_outs_up[57] ;
 wire \ces_1_6_io_outs_up[58] ;
 wire \ces_1_6_io_outs_up[59] ;
 wire \ces_1_6_io_outs_up[5] ;
 wire \ces_1_6_io_outs_up[60] ;
 wire \ces_1_6_io_outs_up[61] ;
 wire \ces_1_6_io_outs_up[62] ;
 wire \ces_1_6_io_outs_up[63] ;
 wire \ces_1_6_io_outs_up[6] ;
 wire \ces_1_6_io_outs_up[7] ;
 wire \ces_1_6_io_outs_up[8] ;
 wire \ces_1_6_io_outs_up[9] ;
 wire \ces_1_7_io_ins_down[0] ;
 wire \ces_1_7_io_ins_down[10] ;
 wire \ces_1_7_io_ins_down[11] ;
 wire \ces_1_7_io_ins_down[12] ;
 wire \ces_1_7_io_ins_down[13] ;
 wire \ces_1_7_io_ins_down[14] ;
 wire \ces_1_7_io_ins_down[15] ;
 wire \ces_1_7_io_ins_down[16] ;
 wire \ces_1_7_io_ins_down[17] ;
 wire \ces_1_7_io_ins_down[18] ;
 wire \ces_1_7_io_ins_down[19] ;
 wire \ces_1_7_io_ins_down[1] ;
 wire \ces_1_7_io_ins_down[20] ;
 wire \ces_1_7_io_ins_down[21] ;
 wire \ces_1_7_io_ins_down[22] ;
 wire \ces_1_7_io_ins_down[23] ;
 wire \ces_1_7_io_ins_down[24] ;
 wire \ces_1_7_io_ins_down[25] ;
 wire \ces_1_7_io_ins_down[26] ;
 wire \ces_1_7_io_ins_down[27] ;
 wire \ces_1_7_io_ins_down[28] ;
 wire \ces_1_7_io_ins_down[29] ;
 wire \ces_1_7_io_ins_down[2] ;
 wire \ces_1_7_io_ins_down[30] ;
 wire \ces_1_7_io_ins_down[31] ;
 wire \ces_1_7_io_ins_down[32] ;
 wire \ces_1_7_io_ins_down[33] ;
 wire \ces_1_7_io_ins_down[34] ;
 wire \ces_1_7_io_ins_down[35] ;
 wire \ces_1_7_io_ins_down[36] ;
 wire \ces_1_7_io_ins_down[37] ;
 wire \ces_1_7_io_ins_down[38] ;
 wire \ces_1_7_io_ins_down[39] ;
 wire \ces_1_7_io_ins_down[3] ;
 wire \ces_1_7_io_ins_down[40] ;
 wire \ces_1_7_io_ins_down[41] ;
 wire \ces_1_7_io_ins_down[42] ;
 wire \ces_1_7_io_ins_down[43] ;
 wire \ces_1_7_io_ins_down[44] ;
 wire \ces_1_7_io_ins_down[45] ;
 wire \ces_1_7_io_ins_down[46] ;
 wire \ces_1_7_io_ins_down[47] ;
 wire \ces_1_7_io_ins_down[48] ;
 wire \ces_1_7_io_ins_down[49] ;
 wire \ces_1_7_io_ins_down[4] ;
 wire \ces_1_7_io_ins_down[50] ;
 wire \ces_1_7_io_ins_down[51] ;
 wire \ces_1_7_io_ins_down[52] ;
 wire \ces_1_7_io_ins_down[53] ;
 wire \ces_1_7_io_ins_down[54] ;
 wire \ces_1_7_io_ins_down[55] ;
 wire \ces_1_7_io_ins_down[56] ;
 wire \ces_1_7_io_ins_down[57] ;
 wire \ces_1_7_io_ins_down[58] ;
 wire \ces_1_7_io_ins_down[59] ;
 wire \ces_1_7_io_ins_down[5] ;
 wire \ces_1_7_io_ins_down[60] ;
 wire \ces_1_7_io_ins_down[61] ;
 wire \ces_1_7_io_ins_down[62] ;
 wire \ces_1_7_io_ins_down[63] ;
 wire \ces_1_7_io_ins_down[6] ;
 wire \ces_1_7_io_ins_down[7] ;
 wire \ces_1_7_io_ins_down[8] ;
 wire \ces_1_7_io_ins_down[9] ;
 wire ces_1_7_io_lsbOuts_0;
 wire ces_1_7_io_lsbOuts_1;
 wire ces_1_7_io_lsbOuts_2;
 wire ces_1_7_io_lsbOuts_3;
 wire ces_1_7_io_lsbOuts_4;
 wire ces_1_7_io_lsbOuts_5;
 wire ces_1_7_io_lsbOuts_6;
 wire ces_1_7_io_lsbOuts_7;
 wire \ces_1_7_io_outs_up[0] ;
 wire \ces_1_7_io_outs_up[10] ;
 wire \ces_1_7_io_outs_up[11] ;
 wire \ces_1_7_io_outs_up[12] ;
 wire \ces_1_7_io_outs_up[13] ;
 wire \ces_1_7_io_outs_up[14] ;
 wire \ces_1_7_io_outs_up[15] ;
 wire \ces_1_7_io_outs_up[16] ;
 wire \ces_1_7_io_outs_up[17] ;
 wire \ces_1_7_io_outs_up[18] ;
 wire \ces_1_7_io_outs_up[19] ;
 wire \ces_1_7_io_outs_up[1] ;
 wire \ces_1_7_io_outs_up[20] ;
 wire \ces_1_7_io_outs_up[21] ;
 wire \ces_1_7_io_outs_up[22] ;
 wire \ces_1_7_io_outs_up[23] ;
 wire \ces_1_7_io_outs_up[24] ;
 wire \ces_1_7_io_outs_up[25] ;
 wire \ces_1_7_io_outs_up[26] ;
 wire \ces_1_7_io_outs_up[27] ;
 wire \ces_1_7_io_outs_up[28] ;
 wire \ces_1_7_io_outs_up[29] ;
 wire \ces_1_7_io_outs_up[2] ;
 wire \ces_1_7_io_outs_up[30] ;
 wire \ces_1_7_io_outs_up[31] ;
 wire \ces_1_7_io_outs_up[32] ;
 wire \ces_1_7_io_outs_up[33] ;
 wire \ces_1_7_io_outs_up[34] ;
 wire \ces_1_7_io_outs_up[35] ;
 wire \ces_1_7_io_outs_up[36] ;
 wire \ces_1_7_io_outs_up[37] ;
 wire \ces_1_7_io_outs_up[38] ;
 wire \ces_1_7_io_outs_up[39] ;
 wire \ces_1_7_io_outs_up[3] ;
 wire \ces_1_7_io_outs_up[40] ;
 wire \ces_1_7_io_outs_up[41] ;
 wire \ces_1_7_io_outs_up[42] ;
 wire \ces_1_7_io_outs_up[43] ;
 wire \ces_1_7_io_outs_up[44] ;
 wire \ces_1_7_io_outs_up[45] ;
 wire \ces_1_7_io_outs_up[46] ;
 wire \ces_1_7_io_outs_up[47] ;
 wire \ces_1_7_io_outs_up[48] ;
 wire \ces_1_7_io_outs_up[49] ;
 wire \ces_1_7_io_outs_up[4] ;
 wire \ces_1_7_io_outs_up[50] ;
 wire \ces_1_7_io_outs_up[51] ;
 wire \ces_1_7_io_outs_up[52] ;
 wire \ces_1_7_io_outs_up[53] ;
 wire \ces_1_7_io_outs_up[54] ;
 wire \ces_1_7_io_outs_up[55] ;
 wire \ces_1_7_io_outs_up[56] ;
 wire \ces_1_7_io_outs_up[57] ;
 wire \ces_1_7_io_outs_up[58] ;
 wire \ces_1_7_io_outs_up[59] ;
 wire \ces_1_7_io_outs_up[5] ;
 wire \ces_1_7_io_outs_up[60] ;
 wire \ces_1_7_io_outs_up[61] ;
 wire \ces_1_7_io_outs_up[62] ;
 wire \ces_1_7_io_outs_up[63] ;
 wire \ces_1_7_io_outs_up[6] ;
 wire \ces_1_7_io_outs_up[7] ;
 wire \ces_1_7_io_outs_up[8] ;
 wire \ces_1_7_io_outs_up[9] ;
 wire \ces_2_0_io_ins_down[0] ;
 wire \ces_2_0_io_ins_down[10] ;
 wire \ces_2_0_io_ins_down[11] ;
 wire \ces_2_0_io_ins_down[12] ;
 wire \ces_2_0_io_ins_down[13] ;
 wire \ces_2_0_io_ins_down[14] ;
 wire \ces_2_0_io_ins_down[15] ;
 wire \ces_2_0_io_ins_down[16] ;
 wire \ces_2_0_io_ins_down[17] ;
 wire \ces_2_0_io_ins_down[18] ;
 wire \ces_2_0_io_ins_down[19] ;
 wire \ces_2_0_io_ins_down[1] ;
 wire \ces_2_0_io_ins_down[20] ;
 wire \ces_2_0_io_ins_down[21] ;
 wire \ces_2_0_io_ins_down[22] ;
 wire \ces_2_0_io_ins_down[23] ;
 wire \ces_2_0_io_ins_down[24] ;
 wire \ces_2_0_io_ins_down[25] ;
 wire \ces_2_0_io_ins_down[26] ;
 wire \ces_2_0_io_ins_down[27] ;
 wire \ces_2_0_io_ins_down[28] ;
 wire \ces_2_0_io_ins_down[29] ;
 wire \ces_2_0_io_ins_down[2] ;
 wire \ces_2_0_io_ins_down[30] ;
 wire \ces_2_0_io_ins_down[31] ;
 wire \ces_2_0_io_ins_down[32] ;
 wire \ces_2_0_io_ins_down[33] ;
 wire \ces_2_0_io_ins_down[34] ;
 wire \ces_2_0_io_ins_down[35] ;
 wire \ces_2_0_io_ins_down[36] ;
 wire \ces_2_0_io_ins_down[37] ;
 wire \ces_2_0_io_ins_down[38] ;
 wire \ces_2_0_io_ins_down[39] ;
 wire \ces_2_0_io_ins_down[3] ;
 wire \ces_2_0_io_ins_down[40] ;
 wire \ces_2_0_io_ins_down[41] ;
 wire \ces_2_0_io_ins_down[42] ;
 wire \ces_2_0_io_ins_down[43] ;
 wire \ces_2_0_io_ins_down[44] ;
 wire \ces_2_0_io_ins_down[45] ;
 wire \ces_2_0_io_ins_down[46] ;
 wire \ces_2_0_io_ins_down[47] ;
 wire \ces_2_0_io_ins_down[48] ;
 wire \ces_2_0_io_ins_down[49] ;
 wire \ces_2_0_io_ins_down[4] ;
 wire \ces_2_0_io_ins_down[50] ;
 wire \ces_2_0_io_ins_down[51] ;
 wire \ces_2_0_io_ins_down[52] ;
 wire \ces_2_0_io_ins_down[53] ;
 wire \ces_2_0_io_ins_down[54] ;
 wire \ces_2_0_io_ins_down[55] ;
 wire \ces_2_0_io_ins_down[56] ;
 wire \ces_2_0_io_ins_down[57] ;
 wire \ces_2_0_io_ins_down[58] ;
 wire \ces_2_0_io_ins_down[59] ;
 wire \ces_2_0_io_ins_down[5] ;
 wire \ces_2_0_io_ins_down[60] ;
 wire \ces_2_0_io_ins_down[61] ;
 wire \ces_2_0_io_ins_down[62] ;
 wire \ces_2_0_io_ins_down[63] ;
 wire \ces_2_0_io_ins_down[6] ;
 wire \ces_2_0_io_ins_down[7] ;
 wire \ces_2_0_io_ins_down[8] ;
 wire \ces_2_0_io_ins_down[9] ;
 wire \ces_2_0_io_ins_left[0] ;
 wire \ces_2_0_io_ins_left[10] ;
 wire \ces_2_0_io_ins_left[11] ;
 wire \ces_2_0_io_ins_left[12] ;
 wire \ces_2_0_io_ins_left[13] ;
 wire \ces_2_0_io_ins_left[14] ;
 wire \ces_2_0_io_ins_left[15] ;
 wire \ces_2_0_io_ins_left[16] ;
 wire \ces_2_0_io_ins_left[17] ;
 wire \ces_2_0_io_ins_left[18] ;
 wire \ces_2_0_io_ins_left[19] ;
 wire \ces_2_0_io_ins_left[1] ;
 wire \ces_2_0_io_ins_left[20] ;
 wire \ces_2_0_io_ins_left[21] ;
 wire \ces_2_0_io_ins_left[22] ;
 wire \ces_2_0_io_ins_left[23] ;
 wire \ces_2_0_io_ins_left[24] ;
 wire \ces_2_0_io_ins_left[25] ;
 wire \ces_2_0_io_ins_left[26] ;
 wire \ces_2_0_io_ins_left[27] ;
 wire \ces_2_0_io_ins_left[28] ;
 wire \ces_2_0_io_ins_left[29] ;
 wire \ces_2_0_io_ins_left[2] ;
 wire \ces_2_0_io_ins_left[30] ;
 wire \ces_2_0_io_ins_left[31] ;
 wire \ces_2_0_io_ins_left[32] ;
 wire \ces_2_0_io_ins_left[33] ;
 wire \ces_2_0_io_ins_left[34] ;
 wire \ces_2_0_io_ins_left[35] ;
 wire \ces_2_0_io_ins_left[36] ;
 wire \ces_2_0_io_ins_left[37] ;
 wire \ces_2_0_io_ins_left[38] ;
 wire \ces_2_0_io_ins_left[39] ;
 wire \ces_2_0_io_ins_left[3] ;
 wire \ces_2_0_io_ins_left[40] ;
 wire \ces_2_0_io_ins_left[41] ;
 wire \ces_2_0_io_ins_left[42] ;
 wire \ces_2_0_io_ins_left[43] ;
 wire \ces_2_0_io_ins_left[44] ;
 wire \ces_2_0_io_ins_left[45] ;
 wire \ces_2_0_io_ins_left[46] ;
 wire \ces_2_0_io_ins_left[47] ;
 wire \ces_2_0_io_ins_left[48] ;
 wire \ces_2_0_io_ins_left[49] ;
 wire \ces_2_0_io_ins_left[4] ;
 wire \ces_2_0_io_ins_left[50] ;
 wire \ces_2_0_io_ins_left[51] ;
 wire \ces_2_0_io_ins_left[52] ;
 wire \ces_2_0_io_ins_left[53] ;
 wire \ces_2_0_io_ins_left[54] ;
 wire \ces_2_0_io_ins_left[55] ;
 wire \ces_2_0_io_ins_left[56] ;
 wire \ces_2_0_io_ins_left[57] ;
 wire \ces_2_0_io_ins_left[58] ;
 wire \ces_2_0_io_ins_left[59] ;
 wire \ces_2_0_io_ins_left[5] ;
 wire \ces_2_0_io_ins_left[60] ;
 wire \ces_2_0_io_ins_left[61] ;
 wire \ces_2_0_io_ins_left[62] ;
 wire \ces_2_0_io_ins_left[63] ;
 wire \ces_2_0_io_ins_left[6] ;
 wire \ces_2_0_io_ins_left[7] ;
 wire \ces_2_0_io_ins_left[8] ;
 wire \ces_2_0_io_ins_left[9] ;
 wire ces_2_0_io_lsbOuts_0;
 wire ces_2_0_io_lsbOuts_1;
 wire ces_2_0_io_lsbOuts_2;
 wire ces_2_0_io_lsbOuts_3;
 wire ces_2_0_io_lsbOuts_4;
 wire ces_2_0_io_lsbOuts_5;
 wire ces_2_0_io_lsbOuts_6;
 wire ces_2_0_io_lsbOuts_7;
 wire \ces_2_0_io_outs_right[0] ;
 wire \ces_2_0_io_outs_right[10] ;
 wire \ces_2_0_io_outs_right[11] ;
 wire \ces_2_0_io_outs_right[12] ;
 wire \ces_2_0_io_outs_right[13] ;
 wire \ces_2_0_io_outs_right[14] ;
 wire \ces_2_0_io_outs_right[15] ;
 wire \ces_2_0_io_outs_right[16] ;
 wire \ces_2_0_io_outs_right[17] ;
 wire \ces_2_0_io_outs_right[18] ;
 wire \ces_2_0_io_outs_right[19] ;
 wire \ces_2_0_io_outs_right[1] ;
 wire \ces_2_0_io_outs_right[20] ;
 wire \ces_2_0_io_outs_right[21] ;
 wire \ces_2_0_io_outs_right[22] ;
 wire \ces_2_0_io_outs_right[23] ;
 wire \ces_2_0_io_outs_right[24] ;
 wire \ces_2_0_io_outs_right[25] ;
 wire \ces_2_0_io_outs_right[26] ;
 wire \ces_2_0_io_outs_right[27] ;
 wire \ces_2_0_io_outs_right[28] ;
 wire \ces_2_0_io_outs_right[29] ;
 wire \ces_2_0_io_outs_right[2] ;
 wire \ces_2_0_io_outs_right[30] ;
 wire \ces_2_0_io_outs_right[31] ;
 wire \ces_2_0_io_outs_right[32] ;
 wire \ces_2_0_io_outs_right[33] ;
 wire \ces_2_0_io_outs_right[34] ;
 wire \ces_2_0_io_outs_right[35] ;
 wire \ces_2_0_io_outs_right[36] ;
 wire \ces_2_0_io_outs_right[37] ;
 wire \ces_2_0_io_outs_right[38] ;
 wire \ces_2_0_io_outs_right[39] ;
 wire \ces_2_0_io_outs_right[3] ;
 wire \ces_2_0_io_outs_right[40] ;
 wire \ces_2_0_io_outs_right[41] ;
 wire \ces_2_0_io_outs_right[42] ;
 wire \ces_2_0_io_outs_right[43] ;
 wire \ces_2_0_io_outs_right[44] ;
 wire \ces_2_0_io_outs_right[45] ;
 wire \ces_2_0_io_outs_right[46] ;
 wire \ces_2_0_io_outs_right[47] ;
 wire \ces_2_0_io_outs_right[48] ;
 wire \ces_2_0_io_outs_right[49] ;
 wire \ces_2_0_io_outs_right[4] ;
 wire \ces_2_0_io_outs_right[50] ;
 wire \ces_2_0_io_outs_right[51] ;
 wire \ces_2_0_io_outs_right[52] ;
 wire \ces_2_0_io_outs_right[53] ;
 wire \ces_2_0_io_outs_right[54] ;
 wire \ces_2_0_io_outs_right[55] ;
 wire \ces_2_0_io_outs_right[56] ;
 wire \ces_2_0_io_outs_right[57] ;
 wire \ces_2_0_io_outs_right[58] ;
 wire \ces_2_0_io_outs_right[59] ;
 wire \ces_2_0_io_outs_right[5] ;
 wire \ces_2_0_io_outs_right[60] ;
 wire \ces_2_0_io_outs_right[61] ;
 wire \ces_2_0_io_outs_right[62] ;
 wire \ces_2_0_io_outs_right[63] ;
 wire \ces_2_0_io_outs_right[6] ;
 wire \ces_2_0_io_outs_right[7] ;
 wire \ces_2_0_io_outs_right[8] ;
 wire \ces_2_0_io_outs_right[9] ;
 wire \ces_2_0_io_outs_up[0] ;
 wire \ces_2_0_io_outs_up[10] ;
 wire \ces_2_0_io_outs_up[11] ;
 wire \ces_2_0_io_outs_up[12] ;
 wire \ces_2_0_io_outs_up[13] ;
 wire \ces_2_0_io_outs_up[14] ;
 wire \ces_2_0_io_outs_up[15] ;
 wire \ces_2_0_io_outs_up[16] ;
 wire \ces_2_0_io_outs_up[17] ;
 wire \ces_2_0_io_outs_up[18] ;
 wire \ces_2_0_io_outs_up[19] ;
 wire \ces_2_0_io_outs_up[1] ;
 wire \ces_2_0_io_outs_up[20] ;
 wire \ces_2_0_io_outs_up[21] ;
 wire \ces_2_0_io_outs_up[22] ;
 wire \ces_2_0_io_outs_up[23] ;
 wire \ces_2_0_io_outs_up[24] ;
 wire \ces_2_0_io_outs_up[25] ;
 wire \ces_2_0_io_outs_up[26] ;
 wire \ces_2_0_io_outs_up[27] ;
 wire \ces_2_0_io_outs_up[28] ;
 wire \ces_2_0_io_outs_up[29] ;
 wire \ces_2_0_io_outs_up[2] ;
 wire \ces_2_0_io_outs_up[30] ;
 wire \ces_2_0_io_outs_up[31] ;
 wire \ces_2_0_io_outs_up[32] ;
 wire \ces_2_0_io_outs_up[33] ;
 wire \ces_2_0_io_outs_up[34] ;
 wire \ces_2_0_io_outs_up[35] ;
 wire \ces_2_0_io_outs_up[36] ;
 wire \ces_2_0_io_outs_up[37] ;
 wire \ces_2_0_io_outs_up[38] ;
 wire \ces_2_0_io_outs_up[39] ;
 wire \ces_2_0_io_outs_up[3] ;
 wire \ces_2_0_io_outs_up[40] ;
 wire \ces_2_0_io_outs_up[41] ;
 wire \ces_2_0_io_outs_up[42] ;
 wire \ces_2_0_io_outs_up[43] ;
 wire \ces_2_0_io_outs_up[44] ;
 wire \ces_2_0_io_outs_up[45] ;
 wire \ces_2_0_io_outs_up[46] ;
 wire \ces_2_0_io_outs_up[47] ;
 wire \ces_2_0_io_outs_up[48] ;
 wire \ces_2_0_io_outs_up[49] ;
 wire \ces_2_0_io_outs_up[4] ;
 wire \ces_2_0_io_outs_up[50] ;
 wire \ces_2_0_io_outs_up[51] ;
 wire \ces_2_0_io_outs_up[52] ;
 wire \ces_2_0_io_outs_up[53] ;
 wire \ces_2_0_io_outs_up[54] ;
 wire \ces_2_0_io_outs_up[55] ;
 wire \ces_2_0_io_outs_up[56] ;
 wire \ces_2_0_io_outs_up[57] ;
 wire \ces_2_0_io_outs_up[58] ;
 wire \ces_2_0_io_outs_up[59] ;
 wire \ces_2_0_io_outs_up[5] ;
 wire \ces_2_0_io_outs_up[60] ;
 wire \ces_2_0_io_outs_up[61] ;
 wire \ces_2_0_io_outs_up[62] ;
 wire \ces_2_0_io_outs_up[63] ;
 wire \ces_2_0_io_outs_up[6] ;
 wire \ces_2_0_io_outs_up[7] ;
 wire \ces_2_0_io_outs_up[8] ;
 wire \ces_2_0_io_outs_up[9] ;
 wire \ces_2_1_io_ins_down[0] ;
 wire \ces_2_1_io_ins_down[10] ;
 wire \ces_2_1_io_ins_down[11] ;
 wire \ces_2_1_io_ins_down[12] ;
 wire \ces_2_1_io_ins_down[13] ;
 wire \ces_2_1_io_ins_down[14] ;
 wire \ces_2_1_io_ins_down[15] ;
 wire \ces_2_1_io_ins_down[16] ;
 wire \ces_2_1_io_ins_down[17] ;
 wire \ces_2_1_io_ins_down[18] ;
 wire \ces_2_1_io_ins_down[19] ;
 wire \ces_2_1_io_ins_down[1] ;
 wire \ces_2_1_io_ins_down[20] ;
 wire \ces_2_1_io_ins_down[21] ;
 wire \ces_2_1_io_ins_down[22] ;
 wire \ces_2_1_io_ins_down[23] ;
 wire \ces_2_1_io_ins_down[24] ;
 wire \ces_2_1_io_ins_down[25] ;
 wire \ces_2_1_io_ins_down[26] ;
 wire \ces_2_1_io_ins_down[27] ;
 wire \ces_2_1_io_ins_down[28] ;
 wire \ces_2_1_io_ins_down[29] ;
 wire \ces_2_1_io_ins_down[2] ;
 wire \ces_2_1_io_ins_down[30] ;
 wire \ces_2_1_io_ins_down[31] ;
 wire \ces_2_1_io_ins_down[32] ;
 wire \ces_2_1_io_ins_down[33] ;
 wire \ces_2_1_io_ins_down[34] ;
 wire \ces_2_1_io_ins_down[35] ;
 wire \ces_2_1_io_ins_down[36] ;
 wire \ces_2_1_io_ins_down[37] ;
 wire \ces_2_1_io_ins_down[38] ;
 wire \ces_2_1_io_ins_down[39] ;
 wire \ces_2_1_io_ins_down[3] ;
 wire \ces_2_1_io_ins_down[40] ;
 wire \ces_2_1_io_ins_down[41] ;
 wire \ces_2_1_io_ins_down[42] ;
 wire \ces_2_1_io_ins_down[43] ;
 wire \ces_2_1_io_ins_down[44] ;
 wire \ces_2_1_io_ins_down[45] ;
 wire \ces_2_1_io_ins_down[46] ;
 wire \ces_2_1_io_ins_down[47] ;
 wire \ces_2_1_io_ins_down[48] ;
 wire \ces_2_1_io_ins_down[49] ;
 wire \ces_2_1_io_ins_down[4] ;
 wire \ces_2_1_io_ins_down[50] ;
 wire \ces_2_1_io_ins_down[51] ;
 wire \ces_2_1_io_ins_down[52] ;
 wire \ces_2_1_io_ins_down[53] ;
 wire \ces_2_1_io_ins_down[54] ;
 wire \ces_2_1_io_ins_down[55] ;
 wire \ces_2_1_io_ins_down[56] ;
 wire \ces_2_1_io_ins_down[57] ;
 wire \ces_2_1_io_ins_down[58] ;
 wire \ces_2_1_io_ins_down[59] ;
 wire \ces_2_1_io_ins_down[5] ;
 wire \ces_2_1_io_ins_down[60] ;
 wire \ces_2_1_io_ins_down[61] ;
 wire \ces_2_1_io_ins_down[62] ;
 wire \ces_2_1_io_ins_down[63] ;
 wire \ces_2_1_io_ins_down[6] ;
 wire \ces_2_1_io_ins_down[7] ;
 wire \ces_2_1_io_ins_down[8] ;
 wire \ces_2_1_io_ins_down[9] ;
 wire \ces_2_1_io_ins_left[0] ;
 wire \ces_2_1_io_ins_left[10] ;
 wire \ces_2_1_io_ins_left[11] ;
 wire \ces_2_1_io_ins_left[12] ;
 wire \ces_2_1_io_ins_left[13] ;
 wire \ces_2_1_io_ins_left[14] ;
 wire \ces_2_1_io_ins_left[15] ;
 wire \ces_2_1_io_ins_left[16] ;
 wire \ces_2_1_io_ins_left[17] ;
 wire \ces_2_1_io_ins_left[18] ;
 wire \ces_2_1_io_ins_left[19] ;
 wire \ces_2_1_io_ins_left[1] ;
 wire \ces_2_1_io_ins_left[20] ;
 wire \ces_2_1_io_ins_left[21] ;
 wire \ces_2_1_io_ins_left[22] ;
 wire \ces_2_1_io_ins_left[23] ;
 wire \ces_2_1_io_ins_left[24] ;
 wire \ces_2_1_io_ins_left[25] ;
 wire \ces_2_1_io_ins_left[26] ;
 wire \ces_2_1_io_ins_left[27] ;
 wire \ces_2_1_io_ins_left[28] ;
 wire \ces_2_1_io_ins_left[29] ;
 wire \ces_2_1_io_ins_left[2] ;
 wire \ces_2_1_io_ins_left[30] ;
 wire \ces_2_1_io_ins_left[31] ;
 wire \ces_2_1_io_ins_left[32] ;
 wire \ces_2_1_io_ins_left[33] ;
 wire \ces_2_1_io_ins_left[34] ;
 wire \ces_2_1_io_ins_left[35] ;
 wire \ces_2_1_io_ins_left[36] ;
 wire \ces_2_1_io_ins_left[37] ;
 wire \ces_2_1_io_ins_left[38] ;
 wire \ces_2_1_io_ins_left[39] ;
 wire \ces_2_1_io_ins_left[3] ;
 wire \ces_2_1_io_ins_left[40] ;
 wire \ces_2_1_io_ins_left[41] ;
 wire \ces_2_1_io_ins_left[42] ;
 wire \ces_2_1_io_ins_left[43] ;
 wire \ces_2_1_io_ins_left[44] ;
 wire \ces_2_1_io_ins_left[45] ;
 wire \ces_2_1_io_ins_left[46] ;
 wire \ces_2_1_io_ins_left[47] ;
 wire \ces_2_1_io_ins_left[48] ;
 wire \ces_2_1_io_ins_left[49] ;
 wire \ces_2_1_io_ins_left[4] ;
 wire \ces_2_1_io_ins_left[50] ;
 wire \ces_2_1_io_ins_left[51] ;
 wire \ces_2_1_io_ins_left[52] ;
 wire \ces_2_1_io_ins_left[53] ;
 wire \ces_2_1_io_ins_left[54] ;
 wire \ces_2_1_io_ins_left[55] ;
 wire \ces_2_1_io_ins_left[56] ;
 wire \ces_2_1_io_ins_left[57] ;
 wire \ces_2_1_io_ins_left[58] ;
 wire \ces_2_1_io_ins_left[59] ;
 wire \ces_2_1_io_ins_left[5] ;
 wire \ces_2_1_io_ins_left[60] ;
 wire \ces_2_1_io_ins_left[61] ;
 wire \ces_2_1_io_ins_left[62] ;
 wire \ces_2_1_io_ins_left[63] ;
 wire \ces_2_1_io_ins_left[6] ;
 wire \ces_2_1_io_ins_left[7] ;
 wire \ces_2_1_io_ins_left[8] ;
 wire \ces_2_1_io_ins_left[9] ;
 wire ces_2_1_io_lsbOuts_0;
 wire ces_2_1_io_lsbOuts_1;
 wire ces_2_1_io_lsbOuts_2;
 wire ces_2_1_io_lsbOuts_3;
 wire ces_2_1_io_lsbOuts_4;
 wire ces_2_1_io_lsbOuts_5;
 wire ces_2_1_io_lsbOuts_6;
 wire ces_2_1_io_lsbOuts_7;
 wire \ces_2_1_io_outs_right[0] ;
 wire \ces_2_1_io_outs_right[10] ;
 wire \ces_2_1_io_outs_right[11] ;
 wire \ces_2_1_io_outs_right[12] ;
 wire \ces_2_1_io_outs_right[13] ;
 wire \ces_2_1_io_outs_right[14] ;
 wire \ces_2_1_io_outs_right[15] ;
 wire \ces_2_1_io_outs_right[16] ;
 wire \ces_2_1_io_outs_right[17] ;
 wire \ces_2_1_io_outs_right[18] ;
 wire \ces_2_1_io_outs_right[19] ;
 wire \ces_2_1_io_outs_right[1] ;
 wire \ces_2_1_io_outs_right[20] ;
 wire \ces_2_1_io_outs_right[21] ;
 wire \ces_2_1_io_outs_right[22] ;
 wire \ces_2_1_io_outs_right[23] ;
 wire \ces_2_1_io_outs_right[24] ;
 wire \ces_2_1_io_outs_right[25] ;
 wire \ces_2_1_io_outs_right[26] ;
 wire \ces_2_1_io_outs_right[27] ;
 wire \ces_2_1_io_outs_right[28] ;
 wire \ces_2_1_io_outs_right[29] ;
 wire \ces_2_1_io_outs_right[2] ;
 wire \ces_2_1_io_outs_right[30] ;
 wire \ces_2_1_io_outs_right[31] ;
 wire \ces_2_1_io_outs_right[32] ;
 wire \ces_2_1_io_outs_right[33] ;
 wire \ces_2_1_io_outs_right[34] ;
 wire \ces_2_1_io_outs_right[35] ;
 wire \ces_2_1_io_outs_right[36] ;
 wire \ces_2_1_io_outs_right[37] ;
 wire \ces_2_1_io_outs_right[38] ;
 wire \ces_2_1_io_outs_right[39] ;
 wire \ces_2_1_io_outs_right[3] ;
 wire \ces_2_1_io_outs_right[40] ;
 wire \ces_2_1_io_outs_right[41] ;
 wire \ces_2_1_io_outs_right[42] ;
 wire \ces_2_1_io_outs_right[43] ;
 wire \ces_2_1_io_outs_right[44] ;
 wire \ces_2_1_io_outs_right[45] ;
 wire \ces_2_1_io_outs_right[46] ;
 wire \ces_2_1_io_outs_right[47] ;
 wire \ces_2_1_io_outs_right[48] ;
 wire \ces_2_1_io_outs_right[49] ;
 wire \ces_2_1_io_outs_right[4] ;
 wire \ces_2_1_io_outs_right[50] ;
 wire \ces_2_1_io_outs_right[51] ;
 wire \ces_2_1_io_outs_right[52] ;
 wire \ces_2_1_io_outs_right[53] ;
 wire \ces_2_1_io_outs_right[54] ;
 wire \ces_2_1_io_outs_right[55] ;
 wire \ces_2_1_io_outs_right[56] ;
 wire \ces_2_1_io_outs_right[57] ;
 wire \ces_2_1_io_outs_right[58] ;
 wire \ces_2_1_io_outs_right[59] ;
 wire \ces_2_1_io_outs_right[5] ;
 wire \ces_2_1_io_outs_right[60] ;
 wire \ces_2_1_io_outs_right[61] ;
 wire \ces_2_1_io_outs_right[62] ;
 wire \ces_2_1_io_outs_right[63] ;
 wire \ces_2_1_io_outs_right[6] ;
 wire \ces_2_1_io_outs_right[7] ;
 wire \ces_2_1_io_outs_right[8] ;
 wire \ces_2_1_io_outs_right[9] ;
 wire \ces_2_1_io_outs_up[0] ;
 wire \ces_2_1_io_outs_up[10] ;
 wire \ces_2_1_io_outs_up[11] ;
 wire \ces_2_1_io_outs_up[12] ;
 wire \ces_2_1_io_outs_up[13] ;
 wire \ces_2_1_io_outs_up[14] ;
 wire \ces_2_1_io_outs_up[15] ;
 wire \ces_2_1_io_outs_up[16] ;
 wire \ces_2_1_io_outs_up[17] ;
 wire \ces_2_1_io_outs_up[18] ;
 wire \ces_2_1_io_outs_up[19] ;
 wire \ces_2_1_io_outs_up[1] ;
 wire \ces_2_1_io_outs_up[20] ;
 wire \ces_2_1_io_outs_up[21] ;
 wire \ces_2_1_io_outs_up[22] ;
 wire \ces_2_1_io_outs_up[23] ;
 wire \ces_2_1_io_outs_up[24] ;
 wire \ces_2_1_io_outs_up[25] ;
 wire \ces_2_1_io_outs_up[26] ;
 wire \ces_2_1_io_outs_up[27] ;
 wire \ces_2_1_io_outs_up[28] ;
 wire \ces_2_1_io_outs_up[29] ;
 wire \ces_2_1_io_outs_up[2] ;
 wire \ces_2_1_io_outs_up[30] ;
 wire \ces_2_1_io_outs_up[31] ;
 wire \ces_2_1_io_outs_up[32] ;
 wire \ces_2_1_io_outs_up[33] ;
 wire \ces_2_1_io_outs_up[34] ;
 wire \ces_2_1_io_outs_up[35] ;
 wire \ces_2_1_io_outs_up[36] ;
 wire \ces_2_1_io_outs_up[37] ;
 wire \ces_2_1_io_outs_up[38] ;
 wire \ces_2_1_io_outs_up[39] ;
 wire \ces_2_1_io_outs_up[3] ;
 wire \ces_2_1_io_outs_up[40] ;
 wire \ces_2_1_io_outs_up[41] ;
 wire \ces_2_1_io_outs_up[42] ;
 wire \ces_2_1_io_outs_up[43] ;
 wire \ces_2_1_io_outs_up[44] ;
 wire \ces_2_1_io_outs_up[45] ;
 wire \ces_2_1_io_outs_up[46] ;
 wire \ces_2_1_io_outs_up[47] ;
 wire \ces_2_1_io_outs_up[48] ;
 wire \ces_2_1_io_outs_up[49] ;
 wire \ces_2_1_io_outs_up[4] ;
 wire \ces_2_1_io_outs_up[50] ;
 wire \ces_2_1_io_outs_up[51] ;
 wire \ces_2_1_io_outs_up[52] ;
 wire \ces_2_1_io_outs_up[53] ;
 wire \ces_2_1_io_outs_up[54] ;
 wire \ces_2_1_io_outs_up[55] ;
 wire \ces_2_1_io_outs_up[56] ;
 wire \ces_2_1_io_outs_up[57] ;
 wire \ces_2_1_io_outs_up[58] ;
 wire \ces_2_1_io_outs_up[59] ;
 wire \ces_2_1_io_outs_up[5] ;
 wire \ces_2_1_io_outs_up[60] ;
 wire \ces_2_1_io_outs_up[61] ;
 wire \ces_2_1_io_outs_up[62] ;
 wire \ces_2_1_io_outs_up[63] ;
 wire \ces_2_1_io_outs_up[6] ;
 wire \ces_2_1_io_outs_up[7] ;
 wire \ces_2_1_io_outs_up[8] ;
 wire \ces_2_1_io_outs_up[9] ;
 wire \ces_2_2_io_ins_down[0] ;
 wire \ces_2_2_io_ins_down[10] ;
 wire \ces_2_2_io_ins_down[11] ;
 wire \ces_2_2_io_ins_down[12] ;
 wire \ces_2_2_io_ins_down[13] ;
 wire \ces_2_2_io_ins_down[14] ;
 wire \ces_2_2_io_ins_down[15] ;
 wire \ces_2_2_io_ins_down[16] ;
 wire \ces_2_2_io_ins_down[17] ;
 wire \ces_2_2_io_ins_down[18] ;
 wire \ces_2_2_io_ins_down[19] ;
 wire \ces_2_2_io_ins_down[1] ;
 wire \ces_2_2_io_ins_down[20] ;
 wire \ces_2_2_io_ins_down[21] ;
 wire \ces_2_2_io_ins_down[22] ;
 wire \ces_2_2_io_ins_down[23] ;
 wire \ces_2_2_io_ins_down[24] ;
 wire \ces_2_2_io_ins_down[25] ;
 wire \ces_2_2_io_ins_down[26] ;
 wire \ces_2_2_io_ins_down[27] ;
 wire \ces_2_2_io_ins_down[28] ;
 wire \ces_2_2_io_ins_down[29] ;
 wire \ces_2_2_io_ins_down[2] ;
 wire \ces_2_2_io_ins_down[30] ;
 wire \ces_2_2_io_ins_down[31] ;
 wire \ces_2_2_io_ins_down[32] ;
 wire \ces_2_2_io_ins_down[33] ;
 wire \ces_2_2_io_ins_down[34] ;
 wire \ces_2_2_io_ins_down[35] ;
 wire \ces_2_2_io_ins_down[36] ;
 wire \ces_2_2_io_ins_down[37] ;
 wire \ces_2_2_io_ins_down[38] ;
 wire \ces_2_2_io_ins_down[39] ;
 wire \ces_2_2_io_ins_down[3] ;
 wire \ces_2_2_io_ins_down[40] ;
 wire \ces_2_2_io_ins_down[41] ;
 wire \ces_2_2_io_ins_down[42] ;
 wire \ces_2_2_io_ins_down[43] ;
 wire \ces_2_2_io_ins_down[44] ;
 wire \ces_2_2_io_ins_down[45] ;
 wire \ces_2_2_io_ins_down[46] ;
 wire \ces_2_2_io_ins_down[47] ;
 wire \ces_2_2_io_ins_down[48] ;
 wire \ces_2_2_io_ins_down[49] ;
 wire \ces_2_2_io_ins_down[4] ;
 wire \ces_2_2_io_ins_down[50] ;
 wire \ces_2_2_io_ins_down[51] ;
 wire \ces_2_2_io_ins_down[52] ;
 wire \ces_2_2_io_ins_down[53] ;
 wire \ces_2_2_io_ins_down[54] ;
 wire \ces_2_2_io_ins_down[55] ;
 wire \ces_2_2_io_ins_down[56] ;
 wire \ces_2_2_io_ins_down[57] ;
 wire \ces_2_2_io_ins_down[58] ;
 wire \ces_2_2_io_ins_down[59] ;
 wire \ces_2_2_io_ins_down[5] ;
 wire \ces_2_2_io_ins_down[60] ;
 wire \ces_2_2_io_ins_down[61] ;
 wire \ces_2_2_io_ins_down[62] ;
 wire \ces_2_2_io_ins_down[63] ;
 wire \ces_2_2_io_ins_down[6] ;
 wire \ces_2_2_io_ins_down[7] ;
 wire \ces_2_2_io_ins_down[8] ;
 wire \ces_2_2_io_ins_down[9] ;
 wire \ces_2_2_io_ins_left[0] ;
 wire \ces_2_2_io_ins_left[10] ;
 wire \ces_2_2_io_ins_left[11] ;
 wire \ces_2_2_io_ins_left[12] ;
 wire \ces_2_2_io_ins_left[13] ;
 wire \ces_2_2_io_ins_left[14] ;
 wire \ces_2_2_io_ins_left[15] ;
 wire \ces_2_2_io_ins_left[16] ;
 wire \ces_2_2_io_ins_left[17] ;
 wire \ces_2_2_io_ins_left[18] ;
 wire \ces_2_2_io_ins_left[19] ;
 wire \ces_2_2_io_ins_left[1] ;
 wire \ces_2_2_io_ins_left[20] ;
 wire \ces_2_2_io_ins_left[21] ;
 wire \ces_2_2_io_ins_left[22] ;
 wire \ces_2_2_io_ins_left[23] ;
 wire \ces_2_2_io_ins_left[24] ;
 wire \ces_2_2_io_ins_left[25] ;
 wire \ces_2_2_io_ins_left[26] ;
 wire \ces_2_2_io_ins_left[27] ;
 wire \ces_2_2_io_ins_left[28] ;
 wire \ces_2_2_io_ins_left[29] ;
 wire \ces_2_2_io_ins_left[2] ;
 wire \ces_2_2_io_ins_left[30] ;
 wire \ces_2_2_io_ins_left[31] ;
 wire \ces_2_2_io_ins_left[32] ;
 wire \ces_2_2_io_ins_left[33] ;
 wire \ces_2_2_io_ins_left[34] ;
 wire \ces_2_2_io_ins_left[35] ;
 wire \ces_2_2_io_ins_left[36] ;
 wire \ces_2_2_io_ins_left[37] ;
 wire \ces_2_2_io_ins_left[38] ;
 wire \ces_2_2_io_ins_left[39] ;
 wire \ces_2_2_io_ins_left[3] ;
 wire \ces_2_2_io_ins_left[40] ;
 wire \ces_2_2_io_ins_left[41] ;
 wire \ces_2_2_io_ins_left[42] ;
 wire \ces_2_2_io_ins_left[43] ;
 wire \ces_2_2_io_ins_left[44] ;
 wire \ces_2_2_io_ins_left[45] ;
 wire \ces_2_2_io_ins_left[46] ;
 wire \ces_2_2_io_ins_left[47] ;
 wire \ces_2_2_io_ins_left[48] ;
 wire \ces_2_2_io_ins_left[49] ;
 wire \ces_2_2_io_ins_left[4] ;
 wire \ces_2_2_io_ins_left[50] ;
 wire \ces_2_2_io_ins_left[51] ;
 wire \ces_2_2_io_ins_left[52] ;
 wire \ces_2_2_io_ins_left[53] ;
 wire \ces_2_2_io_ins_left[54] ;
 wire \ces_2_2_io_ins_left[55] ;
 wire \ces_2_2_io_ins_left[56] ;
 wire \ces_2_2_io_ins_left[57] ;
 wire \ces_2_2_io_ins_left[58] ;
 wire \ces_2_2_io_ins_left[59] ;
 wire \ces_2_2_io_ins_left[5] ;
 wire \ces_2_2_io_ins_left[60] ;
 wire \ces_2_2_io_ins_left[61] ;
 wire \ces_2_2_io_ins_left[62] ;
 wire \ces_2_2_io_ins_left[63] ;
 wire \ces_2_2_io_ins_left[6] ;
 wire \ces_2_2_io_ins_left[7] ;
 wire \ces_2_2_io_ins_left[8] ;
 wire \ces_2_2_io_ins_left[9] ;
 wire ces_2_2_io_lsbOuts_0;
 wire ces_2_2_io_lsbOuts_1;
 wire ces_2_2_io_lsbOuts_2;
 wire ces_2_2_io_lsbOuts_3;
 wire ces_2_2_io_lsbOuts_4;
 wire ces_2_2_io_lsbOuts_5;
 wire ces_2_2_io_lsbOuts_6;
 wire ces_2_2_io_lsbOuts_7;
 wire \ces_2_2_io_outs_right[0] ;
 wire \ces_2_2_io_outs_right[10] ;
 wire \ces_2_2_io_outs_right[11] ;
 wire \ces_2_2_io_outs_right[12] ;
 wire \ces_2_2_io_outs_right[13] ;
 wire \ces_2_2_io_outs_right[14] ;
 wire \ces_2_2_io_outs_right[15] ;
 wire \ces_2_2_io_outs_right[16] ;
 wire \ces_2_2_io_outs_right[17] ;
 wire \ces_2_2_io_outs_right[18] ;
 wire \ces_2_2_io_outs_right[19] ;
 wire \ces_2_2_io_outs_right[1] ;
 wire \ces_2_2_io_outs_right[20] ;
 wire \ces_2_2_io_outs_right[21] ;
 wire \ces_2_2_io_outs_right[22] ;
 wire \ces_2_2_io_outs_right[23] ;
 wire \ces_2_2_io_outs_right[24] ;
 wire \ces_2_2_io_outs_right[25] ;
 wire \ces_2_2_io_outs_right[26] ;
 wire \ces_2_2_io_outs_right[27] ;
 wire \ces_2_2_io_outs_right[28] ;
 wire \ces_2_2_io_outs_right[29] ;
 wire \ces_2_2_io_outs_right[2] ;
 wire \ces_2_2_io_outs_right[30] ;
 wire \ces_2_2_io_outs_right[31] ;
 wire \ces_2_2_io_outs_right[32] ;
 wire \ces_2_2_io_outs_right[33] ;
 wire \ces_2_2_io_outs_right[34] ;
 wire \ces_2_2_io_outs_right[35] ;
 wire \ces_2_2_io_outs_right[36] ;
 wire \ces_2_2_io_outs_right[37] ;
 wire \ces_2_2_io_outs_right[38] ;
 wire \ces_2_2_io_outs_right[39] ;
 wire \ces_2_2_io_outs_right[3] ;
 wire \ces_2_2_io_outs_right[40] ;
 wire \ces_2_2_io_outs_right[41] ;
 wire \ces_2_2_io_outs_right[42] ;
 wire \ces_2_2_io_outs_right[43] ;
 wire \ces_2_2_io_outs_right[44] ;
 wire \ces_2_2_io_outs_right[45] ;
 wire \ces_2_2_io_outs_right[46] ;
 wire \ces_2_2_io_outs_right[47] ;
 wire \ces_2_2_io_outs_right[48] ;
 wire \ces_2_2_io_outs_right[49] ;
 wire \ces_2_2_io_outs_right[4] ;
 wire \ces_2_2_io_outs_right[50] ;
 wire \ces_2_2_io_outs_right[51] ;
 wire \ces_2_2_io_outs_right[52] ;
 wire \ces_2_2_io_outs_right[53] ;
 wire \ces_2_2_io_outs_right[54] ;
 wire \ces_2_2_io_outs_right[55] ;
 wire \ces_2_2_io_outs_right[56] ;
 wire \ces_2_2_io_outs_right[57] ;
 wire \ces_2_2_io_outs_right[58] ;
 wire \ces_2_2_io_outs_right[59] ;
 wire \ces_2_2_io_outs_right[5] ;
 wire \ces_2_2_io_outs_right[60] ;
 wire \ces_2_2_io_outs_right[61] ;
 wire \ces_2_2_io_outs_right[62] ;
 wire \ces_2_2_io_outs_right[63] ;
 wire \ces_2_2_io_outs_right[6] ;
 wire \ces_2_2_io_outs_right[7] ;
 wire \ces_2_2_io_outs_right[8] ;
 wire \ces_2_2_io_outs_right[9] ;
 wire \ces_2_2_io_outs_up[0] ;
 wire \ces_2_2_io_outs_up[10] ;
 wire \ces_2_2_io_outs_up[11] ;
 wire \ces_2_2_io_outs_up[12] ;
 wire \ces_2_2_io_outs_up[13] ;
 wire \ces_2_2_io_outs_up[14] ;
 wire \ces_2_2_io_outs_up[15] ;
 wire \ces_2_2_io_outs_up[16] ;
 wire \ces_2_2_io_outs_up[17] ;
 wire \ces_2_2_io_outs_up[18] ;
 wire \ces_2_2_io_outs_up[19] ;
 wire \ces_2_2_io_outs_up[1] ;
 wire \ces_2_2_io_outs_up[20] ;
 wire \ces_2_2_io_outs_up[21] ;
 wire \ces_2_2_io_outs_up[22] ;
 wire \ces_2_2_io_outs_up[23] ;
 wire \ces_2_2_io_outs_up[24] ;
 wire \ces_2_2_io_outs_up[25] ;
 wire \ces_2_2_io_outs_up[26] ;
 wire \ces_2_2_io_outs_up[27] ;
 wire \ces_2_2_io_outs_up[28] ;
 wire \ces_2_2_io_outs_up[29] ;
 wire \ces_2_2_io_outs_up[2] ;
 wire \ces_2_2_io_outs_up[30] ;
 wire \ces_2_2_io_outs_up[31] ;
 wire \ces_2_2_io_outs_up[32] ;
 wire \ces_2_2_io_outs_up[33] ;
 wire \ces_2_2_io_outs_up[34] ;
 wire \ces_2_2_io_outs_up[35] ;
 wire \ces_2_2_io_outs_up[36] ;
 wire \ces_2_2_io_outs_up[37] ;
 wire \ces_2_2_io_outs_up[38] ;
 wire \ces_2_2_io_outs_up[39] ;
 wire \ces_2_2_io_outs_up[3] ;
 wire \ces_2_2_io_outs_up[40] ;
 wire \ces_2_2_io_outs_up[41] ;
 wire \ces_2_2_io_outs_up[42] ;
 wire \ces_2_2_io_outs_up[43] ;
 wire \ces_2_2_io_outs_up[44] ;
 wire \ces_2_2_io_outs_up[45] ;
 wire \ces_2_2_io_outs_up[46] ;
 wire \ces_2_2_io_outs_up[47] ;
 wire \ces_2_2_io_outs_up[48] ;
 wire \ces_2_2_io_outs_up[49] ;
 wire \ces_2_2_io_outs_up[4] ;
 wire \ces_2_2_io_outs_up[50] ;
 wire \ces_2_2_io_outs_up[51] ;
 wire \ces_2_2_io_outs_up[52] ;
 wire \ces_2_2_io_outs_up[53] ;
 wire \ces_2_2_io_outs_up[54] ;
 wire \ces_2_2_io_outs_up[55] ;
 wire \ces_2_2_io_outs_up[56] ;
 wire \ces_2_2_io_outs_up[57] ;
 wire \ces_2_2_io_outs_up[58] ;
 wire \ces_2_2_io_outs_up[59] ;
 wire \ces_2_2_io_outs_up[5] ;
 wire \ces_2_2_io_outs_up[60] ;
 wire \ces_2_2_io_outs_up[61] ;
 wire \ces_2_2_io_outs_up[62] ;
 wire \ces_2_2_io_outs_up[63] ;
 wire \ces_2_2_io_outs_up[6] ;
 wire \ces_2_2_io_outs_up[7] ;
 wire \ces_2_2_io_outs_up[8] ;
 wire \ces_2_2_io_outs_up[9] ;
 wire \ces_2_3_io_ins_down[0] ;
 wire \ces_2_3_io_ins_down[10] ;
 wire \ces_2_3_io_ins_down[11] ;
 wire \ces_2_3_io_ins_down[12] ;
 wire \ces_2_3_io_ins_down[13] ;
 wire \ces_2_3_io_ins_down[14] ;
 wire \ces_2_3_io_ins_down[15] ;
 wire \ces_2_3_io_ins_down[16] ;
 wire \ces_2_3_io_ins_down[17] ;
 wire \ces_2_3_io_ins_down[18] ;
 wire \ces_2_3_io_ins_down[19] ;
 wire \ces_2_3_io_ins_down[1] ;
 wire \ces_2_3_io_ins_down[20] ;
 wire \ces_2_3_io_ins_down[21] ;
 wire \ces_2_3_io_ins_down[22] ;
 wire \ces_2_3_io_ins_down[23] ;
 wire \ces_2_3_io_ins_down[24] ;
 wire \ces_2_3_io_ins_down[25] ;
 wire \ces_2_3_io_ins_down[26] ;
 wire \ces_2_3_io_ins_down[27] ;
 wire \ces_2_3_io_ins_down[28] ;
 wire \ces_2_3_io_ins_down[29] ;
 wire \ces_2_3_io_ins_down[2] ;
 wire \ces_2_3_io_ins_down[30] ;
 wire \ces_2_3_io_ins_down[31] ;
 wire \ces_2_3_io_ins_down[32] ;
 wire \ces_2_3_io_ins_down[33] ;
 wire \ces_2_3_io_ins_down[34] ;
 wire \ces_2_3_io_ins_down[35] ;
 wire \ces_2_3_io_ins_down[36] ;
 wire \ces_2_3_io_ins_down[37] ;
 wire \ces_2_3_io_ins_down[38] ;
 wire \ces_2_3_io_ins_down[39] ;
 wire \ces_2_3_io_ins_down[3] ;
 wire \ces_2_3_io_ins_down[40] ;
 wire \ces_2_3_io_ins_down[41] ;
 wire \ces_2_3_io_ins_down[42] ;
 wire \ces_2_3_io_ins_down[43] ;
 wire \ces_2_3_io_ins_down[44] ;
 wire \ces_2_3_io_ins_down[45] ;
 wire \ces_2_3_io_ins_down[46] ;
 wire \ces_2_3_io_ins_down[47] ;
 wire \ces_2_3_io_ins_down[48] ;
 wire \ces_2_3_io_ins_down[49] ;
 wire \ces_2_3_io_ins_down[4] ;
 wire \ces_2_3_io_ins_down[50] ;
 wire \ces_2_3_io_ins_down[51] ;
 wire \ces_2_3_io_ins_down[52] ;
 wire \ces_2_3_io_ins_down[53] ;
 wire \ces_2_3_io_ins_down[54] ;
 wire \ces_2_3_io_ins_down[55] ;
 wire \ces_2_3_io_ins_down[56] ;
 wire \ces_2_3_io_ins_down[57] ;
 wire \ces_2_3_io_ins_down[58] ;
 wire \ces_2_3_io_ins_down[59] ;
 wire \ces_2_3_io_ins_down[5] ;
 wire \ces_2_3_io_ins_down[60] ;
 wire \ces_2_3_io_ins_down[61] ;
 wire \ces_2_3_io_ins_down[62] ;
 wire \ces_2_3_io_ins_down[63] ;
 wire \ces_2_3_io_ins_down[6] ;
 wire \ces_2_3_io_ins_down[7] ;
 wire \ces_2_3_io_ins_down[8] ;
 wire \ces_2_3_io_ins_down[9] ;
 wire \ces_2_3_io_ins_left[0] ;
 wire \ces_2_3_io_ins_left[10] ;
 wire \ces_2_3_io_ins_left[11] ;
 wire \ces_2_3_io_ins_left[12] ;
 wire \ces_2_3_io_ins_left[13] ;
 wire \ces_2_3_io_ins_left[14] ;
 wire \ces_2_3_io_ins_left[15] ;
 wire \ces_2_3_io_ins_left[16] ;
 wire \ces_2_3_io_ins_left[17] ;
 wire \ces_2_3_io_ins_left[18] ;
 wire \ces_2_3_io_ins_left[19] ;
 wire \ces_2_3_io_ins_left[1] ;
 wire \ces_2_3_io_ins_left[20] ;
 wire \ces_2_3_io_ins_left[21] ;
 wire \ces_2_3_io_ins_left[22] ;
 wire \ces_2_3_io_ins_left[23] ;
 wire \ces_2_3_io_ins_left[24] ;
 wire \ces_2_3_io_ins_left[25] ;
 wire \ces_2_3_io_ins_left[26] ;
 wire \ces_2_3_io_ins_left[27] ;
 wire \ces_2_3_io_ins_left[28] ;
 wire \ces_2_3_io_ins_left[29] ;
 wire \ces_2_3_io_ins_left[2] ;
 wire \ces_2_3_io_ins_left[30] ;
 wire \ces_2_3_io_ins_left[31] ;
 wire \ces_2_3_io_ins_left[32] ;
 wire \ces_2_3_io_ins_left[33] ;
 wire \ces_2_3_io_ins_left[34] ;
 wire \ces_2_3_io_ins_left[35] ;
 wire \ces_2_3_io_ins_left[36] ;
 wire \ces_2_3_io_ins_left[37] ;
 wire \ces_2_3_io_ins_left[38] ;
 wire \ces_2_3_io_ins_left[39] ;
 wire \ces_2_3_io_ins_left[3] ;
 wire \ces_2_3_io_ins_left[40] ;
 wire \ces_2_3_io_ins_left[41] ;
 wire \ces_2_3_io_ins_left[42] ;
 wire \ces_2_3_io_ins_left[43] ;
 wire \ces_2_3_io_ins_left[44] ;
 wire \ces_2_3_io_ins_left[45] ;
 wire \ces_2_3_io_ins_left[46] ;
 wire \ces_2_3_io_ins_left[47] ;
 wire \ces_2_3_io_ins_left[48] ;
 wire \ces_2_3_io_ins_left[49] ;
 wire \ces_2_3_io_ins_left[4] ;
 wire \ces_2_3_io_ins_left[50] ;
 wire \ces_2_3_io_ins_left[51] ;
 wire \ces_2_3_io_ins_left[52] ;
 wire \ces_2_3_io_ins_left[53] ;
 wire \ces_2_3_io_ins_left[54] ;
 wire \ces_2_3_io_ins_left[55] ;
 wire \ces_2_3_io_ins_left[56] ;
 wire \ces_2_3_io_ins_left[57] ;
 wire \ces_2_3_io_ins_left[58] ;
 wire \ces_2_3_io_ins_left[59] ;
 wire \ces_2_3_io_ins_left[5] ;
 wire \ces_2_3_io_ins_left[60] ;
 wire \ces_2_3_io_ins_left[61] ;
 wire \ces_2_3_io_ins_left[62] ;
 wire \ces_2_3_io_ins_left[63] ;
 wire \ces_2_3_io_ins_left[6] ;
 wire \ces_2_3_io_ins_left[7] ;
 wire \ces_2_3_io_ins_left[8] ;
 wire \ces_2_3_io_ins_left[9] ;
 wire ces_2_3_io_lsbOuts_0;
 wire ces_2_3_io_lsbOuts_1;
 wire ces_2_3_io_lsbOuts_2;
 wire ces_2_3_io_lsbOuts_3;
 wire ces_2_3_io_lsbOuts_4;
 wire ces_2_3_io_lsbOuts_5;
 wire ces_2_3_io_lsbOuts_6;
 wire ces_2_3_io_lsbOuts_7;
 wire \ces_2_3_io_outs_right[0] ;
 wire \ces_2_3_io_outs_right[10] ;
 wire \ces_2_3_io_outs_right[11] ;
 wire \ces_2_3_io_outs_right[12] ;
 wire \ces_2_3_io_outs_right[13] ;
 wire \ces_2_3_io_outs_right[14] ;
 wire \ces_2_3_io_outs_right[15] ;
 wire \ces_2_3_io_outs_right[16] ;
 wire \ces_2_3_io_outs_right[17] ;
 wire \ces_2_3_io_outs_right[18] ;
 wire \ces_2_3_io_outs_right[19] ;
 wire \ces_2_3_io_outs_right[1] ;
 wire \ces_2_3_io_outs_right[20] ;
 wire \ces_2_3_io_outs_right[21] ;
 wire \ces_2_3_io_outs_right[22] ;
 wire \ces_2_3_io_outs_right[23] ;
 wire \ces_2_3_io_outs_right[24] ;
 wire \ces_2_3_io_outs_right[25] ;
 wire \ces_2_3_io_outs_right[26] ;
 wire \ces_2_3_io_outs_right[27] ;
 wire \ces_2_3_io_outs_right[28] ;
 wire \ces_2_3_io_outs_right[29] ;
 wire \ces_2_3_io_outs_right[2] ;
 wire \ces_2_3_io_outs_right[30] ;
 wire \ces_2_3_io_outs_right[31] ;
 wire \ces_2_3_io_outs_right[32] ;
 wire \ces_2_3_io_outs_right[33] ;
 wire \ces_2_3_io_outs_right[34] ;
 wire \ces_2_3_io_outs_right[35] ;
 wire \ces_2_3_io_outs_right[36] ;
 wire \ces_2_3_io_outs_right[37] ;
 wire \ces_2_3_io_outs_right[38] ;
 wire \ces_2_3_io_outs_right[39] ;
 wire \ces_2_3_io_outs_right[3] ;
 wire \ces_2_3_io_outs_right[40] ;
 wire \ces_2_3_io_outs_right[41] ;
 wire \ces_2_3_io_outs_right[42] ;
 wire \ces_2_3_io_outs_right[43] ;
 wire \ces_2_3_io_outs_right[44] ;
 wire \ces_2_3_io_outs_right[45] ;
 wire \ces_2_3_io_outs_right[46] ;
 wire \ces_2_3_io_outs_right[47] ;
 wire \ces_2_3_io_outs_right[48] ;
 wire \ces_2_3_io_outs_right[49] ;
 wire \ces_2_3_io_outs_right[4] ;
 wire \ces_2_3_io_outs_right[50] ;
 wire \ces_2_3_io_outs_right[51] ;
 wire \ces_2_3_io_outs_right[52] ;
 wire \ces_2_3_io_outs_right[53] ;
 wire \ces_2_3_io_outs_right[54] ;
 wire \ces_2_3_io_outs_right[55] ;
 wire \ces_2_3_io_outs_right[56] ;
 wire \ces_2_3_io_outs_right[57] ;
 wire \ces_2_3_io_outs_right[58] ;
 wire \ces_2_3_io_outs_right[59] ;
 wire \ces_2_3_io_outs_right[5] ;
 wire \ces_2_3_io_outs_right[60] ;
 wire \ces_2_3_io_outs_right[61] ;
 wire \ces_2_3_io_outs_right[62] ;
 wire \ces_2_3_io_outs_right[63] ;
 wire \ces_2_3_io_outs_right[6] ;
 wire \ces_2_3_io_outs_right[7] ;
 wire \ces_2_3_io_outs_right[8] ;
 wire \ces_2_3_io_outs_right[9] ;
 wire \ces_2_3_io_outs_up[0] ;
 wire \ces_2_3_io_outs_up[10] ;
 wire \ces_2_3_io_outs_up[11] ;
 wire \ces_2_3_io_outs_up[12] ;
 wire \ces_2_3_io_outs_up[13] ;
 wire \ces_2_3_io_outs_up[14] ;
 wire \ces_2_3_io_outs_up[15] ;
 wire \ces_2_3_io_outs_up[16] ;
 wire \ces_2_3_io_outs_up[17] ;
 wire \ces_2_3_io_outs_up[18] ;
 wire \ces_2_3_io_outs_up[19] ;
 wire \ces_2_3_io_outs_up[1] ;
 wire \ces_2_3_io_outs_up[20] ;
 wire \ces_2_3_io_outs_up[21] ;
 wire \ces_2_3_io_outs_up[22] ;
 wire \ces_2_3_io_outs_up[23] ;
 wire \ces_2_3_io_outs_up[24] ;
 wire \ces_2_3_io_outs_up[25] ;
 wire \ces_2_3_io_outs_up[26] ;
 wire \ces_2_3_io_outs_up[27] ;
 wire \ces_2_3_io_outs_up[28] ;
 wire \ces_2_3_io_outs_up[29] ;
 wire \ces_2_3_io_outs_up[2] ;
 wire \ces_2_3_io_outs_up[30] ;
 wire \ces_2_3_io_outs_up[31] ;
 wire \ces_2_3_io_outs_up[32] ;
 wire \ces_2_3_io_outs_up[33] ;
 wire \ces_2_3_io_outs_up[34] ;
 wire \ces_2_3_io_outs_up[35] ;
 wire \ces_2_3_io_outs_up[36] ;
 wire \ces_2_3_io_outs_up[37] ;
 wire \ces_2_3_io_outs_up[38] ;
 wire \ces_2_3_io_outs_up[39] ;
 wire \ces_2_3_io_outs_up[3] ;
 wire \ces_2_3_io_outs_up[40] ;
 wire \ces_2_3_io_outs_up[41] ;
 wire \ces_2_3_io_outs_up[42] ;
 wire \ces_2_3_io_outs_up[43] ;
 wire \ces_2_3_io_outs_up[44] ;
 wire \ces_2_3_io_outs_up[45] ;
 wire \ces_2_3_io_outs_up[46] ;
 wire \ces_2_3_io_outs_up[47] ;
 wire \ces_2_3_io_outs_up[48] ;
 wire \ces_2_3_io_outs_up[49] ;
 wire \ces_2_3_io_outs_up[4] ;
 wire \ces_2_3_io_outs_up[50] ;
 wire \ces_2_3_io_outs_up[51] ;
 wire \ces_2_3_io_outs_up[52] ;
 wire \ces_2_3_io_outs_up[53] ;
 wire \ces_2_3_io_outs_up[54] ;
 wire \ces_2_3_io_outs_up[55] ;
 wire \ces_2_3_io_outs_up[56] ;
 wire \ces_2_3_io_outs_up[57] ;
 wire \ces_2_3_io_outs_up[58] ;
 wire \ces_2_3_io_outs_up[59] ;
 wire \ces_2_3_io_outs_up[5] ;
 wire \ces_2_3_io_outs_up[60] ;
 wire \ces_2_3_io_outs_up[61] ;
 wire \ces_2_3_io_outs_up[62] ;
 wire \ces_2_3_io_outs_up[63] ;
 wire \ces_2_3_io_outs_up[6] ;
 wire \ces_2_3_io_outs_up[7] ;
 wire \ces_2_3_io_outs_up[8] ;
 wire \ces_2_3_io_outs_up[9] ;
 wire \ces_2_4_io_ins_down[0] ;
 wire \ces_2_4_io_ins_down[10] ;
 wire \ces_2_4_io_ins_down[11] ;
 wire \ces_2_4_io_ins_down[12] ;
 wire \ces_2_4_io_ins_down[13] ;
 wire \ces_2_4_io_ins_down[14] ;
 wire \ces_2_4_io_ins_down[15] ;
 wire \ces_2_4_io_ins_down[16] ;
 wire \ces_2_4_io_ins_down[17] ;
 wire \ces_2_4_io_ins_down[18] ;
 wire \ces_2_4_io_ins_down[19] ;
 wire \ces_2_4_io_ins_down[1] ;
 wire \ces_2_4_io_ins_down[20] ;
 wire \ces_2_4_io_ins_down[21] ;
 wire \ces_2_4_io_ins_down[22] ;
 wire \ces_2_4_io_ins_down[23] ;
 wire \ces_2_4_io_ins_down[24] ;
 wire \ces_2_4_io_ins_down[25] ;
 wire \ces_2_4_io_ins_down[26] ;
 wire \ces_2_4_io_ins_down[27] ;
 wire \ces_2_4_io_ins_down[28] ;
 wire \ces_2_4_io_ins_down[29] ;
 wire \ces_2_4_io_ins_down[2] ;
 wire \ces_2_4_io_ins_down[30] ;
 wire \ces_2_4_io_ins_down[31] ;
 wire \ces_2_4_io_ins_down[32] ;
 wire \ces_2_4_io_ins_down[33] ;
 wire \ces_2_4_io_ins_down[34] ;
 wire \ces_2_4_io_ins_down[35] ;
 wire \ces_2_4_io_ins_down[36] ;
 wire \ces_2_4_io_ins_down[37] ;
 wire \ces_2_4_io_ins_down[38] ;
 wire \ces_2_4_io_ins_down[39] ;
 wire \ces_2_4_io_ins_down[3] ;
 wire \ces_2_4_io_ins_down[40] ;
 wire \ces_2_4_io_ins_down[41] ;
 wire \ces_2_4_io_ins_down[42] ;
 wire \ces_2_4_io_ins_down[43] ;
 wire \ces_2_4_io_ins_down[44] ;
 wire \ces_2_4_io_ins_down[45] ;
 wire \ces_2_4_io_ins_down[46] ;
 wire \ces_2_4_io_ins_down[47] ;
 wire \ces_2_4_io_ins_down[48] ;
 wire \ces_2_4_io_ins_down[49] ;
 wire \ces_2_4_io_ins_down[4] ;
 wire \ces_2_4_io_ins_down[50] ;
 wire \ces_2_4_io_ins_down[51] ;
 wire \ces_2_4_io_ins_down[52] ;
 wire \ces_2_4_io_ins_down[53] ;
 wire \ces_2_4_io_ins_down[54] ;
 wire \ces_2_4_io_ins_down[55] ;
 wire \ces_2_4_io_ins_down[56] ;
 wire \ces_2_4_io_ins_down[57] ;
 wire \ces_2_4_io_ins_down[58] ;
 wire \ces_2_4_io_ins_down[59] ;
 wire \ces_2_4_io_ins_down[5] ;
 wire \ces_2_4_io_ins_down[60] ;
 wire \ces_2_4_io_ins_down[61] ;
 wire \ces_2_4_io_ins_down[62] ;
 wire \ces_2_4_io_ins_down[63] ;
 wire \ces_2_4_io_ins_down[6] ;
 wire \ces_2_4_io_ins_down[7] ;
 wire \ces_2_4_io_ins_down[8] ;
 wire \ces_2_4_io_ins_down[9] ;
 wire \ces_2_4_io_ins_left[0] ;
 wire \ces_2_4_io_ins_left[10] ;
 wire \ces_2_4_io_ins_left[11] ;
 wire \ces_2_4_io_ins_left[12] ;
 wire \ces_2_4_io_ins_left[13] ;
 wire \ces_2_4_io_ins_left[14] ;
 wire \ces_2_4_io_ins_left[15] ;
 wire \ces_2_4_io_ins_left[16] ;
 wire \ces_2_4_io_ins_left[17] ;
 wire \ces_2_4_io_ins_left[18] ;
 wire \ces_2_4_io_ins_left[19] ;
 wire \ces_2_4_io_ins_left[1] ;
 wire \ces_2_4_io_ins_left[20] ;
 wire \ces_2_4_io_ins_left[21] ;
 wire \ces_2_4_io_ins_left[22] ;
 wire \ces_2_4_io_ins_left[23] ;
 wire \ces_2_4_io_ins_left[24] ;
 wire \ces_2_4_io_ins_left[25] ;
 wire \ces_2_4_io_ins_left[26] ;
 wire \ces_2_4_io_ins_left[27] ;
 wire \ces_2_4_io_ins_left[28] ;
 wire \ces_2_4_io_ins_left[29] ;
 wire \ces_2_4_io_ins_left[2] ;
 wire \ces_2_4_io_ins_left[30] ;
 wire \ces_2_4_io_ins_left[31] ;
 wire \ces_2_4_io_ins_left[32] ;
 wire \ces_2_4_io_ins_left[33] ;
 wire \ces_2_4_io_ins_left[34] ;
 wire \ces_2_4_io_ins_left[35] ;
 wire \ces_2_4_io_ins_left[36] ;
 wire \ces_2_4_io_ins_left[37] ;
 wire \ces_2_4_io_ins_left[38] ;
 wire \ces_2_4_io_ins_left[39] ;
 wire \ces_2_4_io_ins_left[3] ;
 wire \ces_2_4_io_ins_left[40] ;
 wire \ces_2_4_io_ins_left[41] ;
 wire \ces_2_4_io_ins_left[42] ;
 wire \ces_2_4_io_ins_left[43] ;
 wire \ces_2_4_io_ins_left[44] ;
 wire \ces_2_4_io_ins_left[45] ;
 wire \ces_2_4_io_ins_left[46] ;
 wire \ces_2_4_io_ins_left[47] ;
 wire \ces_2_4_io_ins_left[48] ;
 wire \ces_2_4_io_ins_left[49] ;
 wire \ces_2_4_io_ins_left[4] ;
 wire \ces_2_4_io_ins_left[50] ;
 wire \ces_2_4_io_ins_left[51] ;
 wire \ces_2_4_io_ins_left[52] ;
 wire \ces_2_4_io_ins_left[53] ;
 wire \ces_2_4_io_ins_left[54] ;
 wire \ces_2_4_io_ins_left[55] ;
 wire \ces_2_4_io_ins_left[56] ;
 wire \ces_2_4_io_ins_left[57] ;
 wire \ces_2_4_io_ins_left[58] ;
 wire \ces_2_4_io_ins_left[59] ;
 wire \ces_2_4_io_ins_left[5] ;
 wire \ces_2_4_io_ins_left[60] ;
 wire \ces_2_4_io_ins_left[61] ;
 wire \ces_2_4_io_ins_left[62] ;
 wire \ces_2_4_io_ins_left[63] ;
 wire \ces_2_4_io_ins_left[6] ;
 wire \ces_2_4_io_ins_left[7] ;
 wire \ces_2_4_io_ins_left[8] ;
 wire \ces_2_4_io_ins_left[9] ;
 wire ces_2_4_io_lsbOuts_0;
 wire ces_2_4_io_lsbOuts_1;
 wire ces_2_4_io_lsbOuts_2;
 wire ces_2_4_io_lsbOuts_3;
 wire ces_2_4_io_lsbOuts_4;
 wire ces_2_4_io_lsbOuts_5;
 wire ces_2_4_io_lsbOuts_6;
 wire ces_2_4_io_lsbOuts_7;
 wire \ces_2_4_io_outs_right[0] ;
 wire \ces_2_4_io_outs_right[10] ;
 wire \ces_2_4_io_outs_right[11] ;
 wire \ces_2_4_io_outs_right[12] ;
 wire \ces_2_4_io_outs_right[13] ;
 wire \ces_2_4_io_outs_right[14] ;
 wire \ces_2_4_io_outs_right[15] ;
 wire \ces_2_4_io_outs_right[16] ;
 wire \ces_2_4_io_outs_right[17] ;
 wire \ces_2_4_io_outs_right[18] ;
 wire \ces_2_4_io_outs_right[19] ;
 wire \ces_2_4_io_outs_right[1] ;
 wire \ces_2_4_io_outs_right[20] ;
 wire \ces_2_4_io_outs_right[21] ;
 wire \ces_2_4_io_outs_right[22] ;
 wire \ces_2_4_io_outs_right[23] ;
 wire \ces_2_4_io_outs_right[24] ;
 wire \ces_2_4_io_outs_right[25] ;
 wire \ces_2_4_io_outs_right[26] ;
 wire \ces_2_4_io_outs_right[27] ;
 wire \ces_2_4_io_outs_right[28] ;
 wire \ces_2_4_io_outs_right[29] ;
 wire \ces_2_4_io_outs_right[2] ;
 wire \ces_2_4_io_outs_right[30] ;
 wire \ces_2_4_io_outs_right[31] ;
 wire \ces_2_4_io_outs_right[32] ;
 wire \ces_2_4_io_outs_right[33] ;
 wire \ces_2_4_io_outs_right[34] ;
 wire \ces_2_4_io_outs_right[35] ;
 wire \ces_2_4_io_outs_right[36] ;
 wire \ces_2_4_io_outs_right[37] ;
 wire \ces_2_4_io_outs_right[38] ;
 wire \ces_2_4_io_outs_right[39] ;
 wire \ces_2_4_io_outs_right[3] ;
 wire \ces_2_4_io_outs_right[40] ;
 wire \ces_2_4_io_outs_right[41] ;
 wire \ces_2_4_io_outs_right[42] ;
 wire \ces_2_4_io_outs_right[43] ;
 wire \ces_2_4_io_outs_right[44] ;
 wire \ces_2_4_io_outs_right[45] ;
 wire \ces_2_4_io_outs_right[46] ;
 wire \ces_2_4_io_outs_right[47] ;
 wire \ces_2_4_io_outs_right[48] ;
 wire \ces_2_4_io_outs_right[49] ;
 wire \ces_2_4_io_outs_right[4] ;
 wire \ces_2_4_io_outs_right[50] ;
 wire \ces_2_4_io_outs_right[51] ;
 wire \ces_2_4_io_outs_right[52] ;
 wire \ces_2_4_io_outs_right[53] ;
 wire \ces_2_4_io_outs_right[54] ;
 wire \ces_2_4_io_outs_right[55] ;
 wire \ces_2_4_io_outs_right[56] ;
 wire \ces_2_4_io_outs_right[57] ;
 wire \ces_2_4_io_outs_right[58] ;
 wire \ces_2_4_io_outs_right[59] ;
 wire \ces_2_4_io_outs_right[5] ;
 wire \ces_2_4_io_outs_right[60] ;
 wire \ces_2_4_io_outs_right[61] ;
 wire \ces_2_4_io_outs_right[62] ;
 wire \ces_2_4_io_outs_right[63] ;
 wire \ces_2_4_io_outs_right[6] ;
 wire \ces_2_4_io_outs_right[7] ;
 wire \ces_2_4_io_outs_right[8] ;
 wire \ces_2_4_io_outs_right[9] ;
 wire \ces_2_4_io_outs_up[0] ;
 wire \ces_2_4_io_outs_up[10] ;
 wire \ces_2_4_io_outs_up[11] ;
 wire \ces_2_4_io_outs_up[12] ;
 wire \ces_2_4_io_outs_up[13] ;
 wire \ces_2_4_io_outs_up[14] ;
 wire \ces_2_4_io_outs_up[15] ;
 wire \ces_2_4_io_outs_up[16] ;
 wire \ces_2_4_io_outs_up[17] ;
 wire \ces_2_4_io_outs_up[18] ;
 wire \ces_2_4_io_outs_up[19] ;
 wire \ces_2_4_io_outs_up[1] ;
 wire \ces_2_4_io_outs_up[20] ;
 wire \ces_2_4_io_outs_up[21] ;
 wire \ces_2_4_io_outs_up[22] ;
 wire \ces_2_4_io_outs_up[23] ;
 wire \ces_2_4_io_outs_up[24] ;
 wire \ces_2_4_io_outs_up[25] ;
 wire \ces_2_4_io_outs_up[26] ;
 wire \ces_2_4_io_outs_up[27] ;
 wire \ces_2_4_io_outs_up[28] ;
 wire \ces_2_4_io_outs_up[29] ;
 wire \ces_2_4_io_outs_up[2] ;
 wire \ces_2_4_io_outs_up[30] ;
 wire \ces_2_4_io_outs_up[31] ;
 wire \ces_2_4_io_outs_up[32] ;
 wire \ces_2_4_io_outs_up[33] ;
 wire \ces_2_4_io_outs_up[34] ;
 wire \ces_2_4_io_outs_up[35] ;
 wire \ces_2_4_io_outs_up[36] ;
 wire \ces_2_4_io_outs_up[37] ;
 wire \ces_2_4_io_outs_up[38] ;
 wire \ces_2_4_io_outs_up[39] ;
 wire \ces_2_4_io_outs_up[3] ;
 wire \ces_2_4_io_outs_up[40] ;
 wire \ces_2_4_io_outs_up[41] ;
 wire \ces_2_4_io_outs_up[42] ;
 wire \ces_2_4_io_outs_up[43] ;
 wire \ces_2_4_io_outs_up[44] ;
 wire \ces_2_4_io_outs_up[45] ;
 wire \ces_2_4_io_outs_up[46] ;
 wire \ces_2_4_io_outs_up[47] ;
 wire \ces_2_4_io_outs_up[48] ;
 wire \ces_2_4_io_outs_up[49] ;
 wire \ces_2_4_io_outs_up[4] ;
 wire \ces_2_4_io_outs_up[50] ;
 wire \ces_2_4_io_outs_up[51] ;
 wire \ces_2_4_io_outs_up[52] ;
 wire \ces_2_4_io_outs_up[53] ;
 wire \ces_2_4_io_outs_up[54] ;
 wire \ces_2_4_io_outs_up[55] ;
 wire \ces_2_4_io_outs_up[56] ;
 wire \ces_2_4_io_outs_up[57] ;
 wire \ces_2_4_io_outs_up[58] ;
 wire \ces_2_4_io_outs_up[59] ;
 wire \ces_2_4_io_outs_up[5] ;
 wire \ces_2_4_io_outs_up[60] ;
 wire \ces_2_4_io_outs_up[61] ;
 wire \ces_2_4_io_outs_up[62] ;
 wire \ces_2_4_io_outs_up[63] ;
 wire \ces_2_4_io_outs_up[6] ;
 wire \ces_2_4_io_outs_up[7] ;
 wire \ces_2_4_io_outs_up[8] ;
 wire \ces_2_4_io_outs_up[9] ;
 wire \ces_2_5_io_ins_down[0] ;
 wire \ces_2_5_io_ins_down[10] ;
 wire \ces_2_5_io_ins_down[11] ;
 wire \ces_2_5_io_ins_down[12] ;
 wire \ces_2_5_io_ins_down[13] ;
 wire \ces_2_5_io_ins_down[14] ;
 wire \ces_2_5_io_ins_down[15] ;
 wire \ces_2_5_io_ins_down[16] ;
 wire \ces_2_5_io_ins_down[17] ;
 wire \ces_2_5_io_ins_down[18] ;
 wire \ces_2_5_io_ins_down[19] ;
 wire \ces_2_5_io_ins_down[1] ;
 wire \ces_2_5_io_ins_down[20] ;
 wire \ces_2_5_io_ins_down[21] ;
 wire \ces_2_5_io_ins_down[22] ;
 wire \ces_2_5_io_ins_down[23] ;
 wire \ces_2_5_io_ins_down[24] ;
 wire \ces_2_5_io_ins_down[25] ;
 wire \ces_2_5_io_ins_down[26] ;
 wire \ces_2_5_io_ins_down[27] ;
 wire \ces_2_5_io_ins_down[28] ;
 wire \ces_2_5_io_ins_down[29] ;
 wire \ces_2_5_io_ins_down[2] ;
 wire \ces_2_5_io_ins_down[30] ;
 wire \ces_2_5_io_ins_down[31] ;
 wire \ces_2_5_io_ins_down[32] ;
 wire \ces_2_5_io_ins_down[33] ;
 wire \ces_2_5_io_ins_down[34] ;
 wire \ces_2_5_io_ins_down[35] ;
 wire \ces_2_5_io_ins_down[36] ;
 wire \ces_2_5_io_ins_down[37] ;
 wire \ces_2_5_io_ins_down[38] ;
 wire \ces_2_5_io_ins_down[39] ;
 wire \ces_2_5_io_ins_down[3] ;
 wire \ces_2_5_io_ins_down[40] ;
 wire \ces_2_5_io_ins_down[41] ;
 wire \ces_2_5_io_ins_down[42] ;
 wire \ces_2_5_io_ins_down[43] ;
 wire \ces_2_5_io_ins_down[44] ;
 wire \ces_2_5_io_ins_down[45] ;
 wire \ces_2_5_io_ins_down[46] ;
 wire \ces_2_5_io_ins_down[47] ;
 wire \ces_2_5_io_ins_down[48] ;
 wire \ces_2_5_io_ins_down[49] ;
 wire \ces_2_5_io_ins_down[4] ;
 wire \ces_2_5_io_ins_down[50] ;
 wire \ces_2_5_io_ins_down[51] ;
 wire \ces_2_5_io_ins_down[52] ;
 wire \ces_2_5_io_ins_down[53] ;
 wire \ces_2_5_io_ins_down[54] ;
 wire \ces_2_5_io_ins_down[55] ;
 wire \ces_2_5_io_ins_down[56] ;
 wire \ces_2_5_io_ins_down[57] ;
 wire \ces_2_5_io_ins_down[58] ;
 wire \ces_2_5_io_ins_down[59] ;
 wire \ces_2_5_io_ins_down[5] ;
 wire \ces_2_5_io_ins_down[60] ;
 wire \ces_2_5_io_ins_down[61] ;
 wire \ces_2_5_io_ins_down[62] ;
 wire \ces_2_5_io_ins_down[63] ;
 wire \ces_2_5_io_ins_down[6] ;
 wire \ces_2_5_io_ins_down[7] ;
 wire \ces_2_5_io_ins_down[8] ;
 wire \ces_2_5_io_ins_down[9] ;
 wire \ces_2_5_io_ins_left[0] ;
 wire \ces_2_5_io_ins_left[10] ;
 wire \ces_2_5_io_ins_left[11] ;
 wire \ces_2_5_io_ins_left[12] ;
 wire \ces_2_5_io_ins_left[13] ;
 wire \ces_2_5_io_ins_left[14] ;
 wire \ces_2_5_io_ins_left[15] ;
 wire \ces_2_5_io_ins_left[16] ;
 wire \ces_2_5_io_ins_left[17] ;
 wire \ces_2_5_io_ins_left[18] ;
 wire \ces_2_5_io_ins_left[19] ;
 wire \ces_2_5_io_ins_left[1] ;
 wire \ces_2_5_io_ins_left[20] ;
 wire \ces_2_5_io_ins_left[21] ;
 wire \ces_2_5_io_ins_left[22] ;
 wire \ces_2_5_io_ins_left[23] ;
 wire \ces_2_5_io_ins_left[24] ;
 wire \ces_2_5_io_ins_left[25] ;
 wire \ces_2_5_io_ins_left[26] ;
 wire \ces_2_5_io_ins_left[27] ;
 wire \ces_2_5_io_ins_left[28] ;
 wire \ces_2_5_io_ins_left[29] ;
 wire \ces_2_5_io_ins_left[2] ;
 wire \ces_2_5_io_ins_left[30] ;
 wire \ces_2_5_io_ins_left[31] ;
 wire \ces_2_5_io_ins_left[32] ;
 wire \ces_2_5_io_ins_left[33] ;
 wire \ces_2_5_io_ins_left[34] ;
 wire \ces_2_5_io_ins_left[35] ;
 wire \ces_2_5_io_ins_left[36] ;
 wire \ces_2_5_io_ins_left[37] ;
 wire \ces_2_5_io_ins_left[38] ;
 wire \ces_2_5_io_ins_left[39] ;
 wire \ces_2_5_io_ins_left[3] ;
 wire \ces_2_5_io_ins_left[40] ;
 wire \ces_2_5_io_ins_left[41] ;
 wire \ces_2_5_io_ins_left[42] ;
 wire \ces_2_5_io_ins_left[43] ;
 wire \ces_2_5_io_ins_left[44] ;
 wire \ces_2_5_io_ins_left[45] ;
 wire \ces_2_5_io_ins_left[46] ;
 wire \ces_2_5_io_ins_left[47] ;
 wire \ces_2_5_io_ins_left[48] ;
 wire \ces_2_5_io_ins_left[49] ;
 wire \ces_2_5_io_ins_left[4] ;
 wire \ces_2_5_io_ins_left[50] ;
 wire \ces_2_5_io_ins_left[51] ;
 wire \ces_2_5_io_ins_left[52] ;
 wire \ces_2_5_io_ins_left[53] ;
 wire \ces_2_5_io_ins_left[54] ;
 wire \ces_2_5_io_ins_left[55] ;
 wire \ces_2_5_io_ins_left[56] ;
 wire \ces_2_5_io_ins_left[57] ;
 wire \ces_2_5_io_ins_left[58] ;
 wire \ces_2_5_io_ins_left[59] ;
 wire \ces_2_5_io_ins_left[5] ;
 wire \ces_2_5_io_ins_left[60] ;
 wire \ces_2_5_io_ins_left[61] ;
 wire \ces_2_5_io_ins_left[62] ;
 wire \ces_2_5_io_ins_left[63] ;
 wire \ces_2_5_io_ins_left[6] ;
 wire \ces_2_5_io_ins_left[7] ;
 wire \ces_2_5_io_ins_left[8] ;
 wire \ces_2_5_io_ins_left[9] ;
 wire ces_2_5_io_lsbOuts_0;
 wire ces_2_5_io_lsbOuts_1;
 wire ces_2_5_io_lsbOuts_2;
 wire ces_2_5_io_lsbOuts_3;
 wire ces_2_5_io_lsbOuts_4;
 wire ces_2_5_io_lsbOuts_5;
 wire ces_2_5_io_lsbOuts_6;
 wire ces_2_5_io_lsbOuts_7;
 wire \ces_2_5_io_outs_right[0] ;
 wire \ces_2_5_io_outs_right[10] ;
 wire \ces_2_5_io_outs_right[11] ;
 wire \ces_2_5_io_outs_right[12] ;
 wire \ces_2_5_io_outs_right[13] ;
 wire \ces_2_5_io_outs_right[14] ;
 wire \ces_2_5_io_outs_right[15] ;
 wire \ces_2_5_io_outs_right[16] ;
 wire \ces_2_5_io_outs_right[17] ;
 wire \ces_2_5_io_outs_right[18] ;
 wire \ces_2_5_io_outs_right[19] ;
 wire \ces_2_5_io_outs_right[1] ;
 wire \ces_2_5_io_outs_right[20] ;
 wire \ces_2_5_io_outs_right[21] ;
 wire \ces_2_5_io_outs_right[22] ;
 wire \ces_2_5_io_outs_right[23] ;
 wire \ces_2_5_io_outs_right[24] ;
 wire \ces_2_5_io_outs_right[25] ;
 wire \ces_2_5_io_outs_right[26] ;
 wire \ces_2_5_io_outs_right[27] ;
 wire \ces_2_5_io_outs_right[28] ;
 wire \ces_2_5_io_outs_right[29] ;
 wire \ces_2_5_io_outs_right[2] ;
 wire \ces_2_5_io_outs_right[30] ;
 wire \ces_2_5_io_outs_right[31] ;
 wire \ces_2_5_io_outs_right[32] ;
 wire \ces_2_5_io_outs_right[33] ;
 wire \ces_2_5_io_outs_right[34] ;
 wire \ces_2_5_io_outs_right[35] ;
 wire \ces_2_5_io_outs_right[36] ;
 wire \ces_2_5_io_outs_right[37] ;
 wire \ces_2_5_io_outs_right[38] ;
 wire \ces_2_5_io_outs_right[39] ;
 wire \ces_2_5_io_outs_right[3] ;
 wire \ces_2_5_io_outs_right[40] ;
 wire \ces_2_5_io_outs_right[41] ;
 wire \ces_2_5_io_outs_right[42] ;
 wire \ces_2_5_io_outs_right[43] ;
 wire \ces_2_5_io_outs_right[44] ;
 wire \ces_2_5_io_outs_right[45] ;
 wire \ces_2_5_io_outs_right[46] ;
 wire \ces_2_5_io_outs_right[47] ;
 wire \ces_2_5_io_outs_right[48] ;
 wire \ces_2_5_io_outs_right[49] ;
 wire \ces_2_5_io_outs_right[4] ;
 wire \ces_2_5_io_outs_right[50] ;
 wire \ces_2_5_io_outs_right[51] ;
 wire \ces_2_5_io_outs_right[52] ;
 wire \ces_2_5_io_outs_right[53] ;
 wire \ces_2_5_io_outs_right[54] ;
 wire \ces_2_5_io_outs_right[55] ;
 wire \ces_2_5_io_outs_right[56] ;
 wire \ces_2_5_io_outs_right[57] ;
 wire \ces_2_5_io_outs_right[58] ;
 wire \ces_2_5_io_outs_right[59] ;
 wire \ces_2_5_io_outs_right[5] ;
 wire \ces_2_5_io_outs_right[60] ;
 wire \ces_2_5_io_outs_right[61] ;
 wire \ces_2_5_io_outs_right[62] ;
 wire \ces_2_5_io_outs_right[63] ;
 wire \ces_2_5_io_outs_right[6] ;
 wire \ces_2_5_io_outs_right[7] ;
 wire \ces_2_5_io_outs_right[8] ;
 wire \ces_2_5_io_outs_right[9] ;
 wire \ces_2_5_io_outs_up[0] ;
 wire \ces_2_5_io_outs_up[10] ;
 wire \ces_2_5_io_outs_up[11] ;
 wire \ces_2_5_io_outs_up[12] ;
 wire \ces_2_5_io_outs_up[13] ;
 wire \ces_2_5_io_outs_up[14] ;
 wire \ces_2_5_io_outs_up[15] ;
 wire \ces_2_5_io_outs_up[16] ;
 wire \ces_2_5_io_outs_up[17] ;
 wire \ces_2_5_io_outs_up[18] ;
 wire \ces_2_5_io_outs_up[19] ;
 wire \ces_2_5_io_outs_up[1] ;
 wire \ces_2_5_io_outs_up[20] ;
 wire \ces_2_5_io_outs_up[21] ;
 wire \ces_2_5_io_outs_up[22] ;
 wire \ces_2_5_io_outs_up[23] ;
 wire \ces_2_5_io_outs_up[24] ;
 wire \ces_2_5_io_outs_up[25] ;
 wire \ces_2_5_io_outs_up[26] ;
 wire \ces_2_5_io_outs_up[27] ;
 wire \ces_2_5_io_outs_up[28] ;
 wire \ces_2_5_io_outs_up[29] ;
 wire \ces_2_5_io_outs_up[2] ;
 wire \ces_2_5_io_outs_up[30] ;
 wire \ces_2_5_io_outs_up[31] ;
 wire \ces_2_5_io_outs_up[32] ;
 wire \ces_2_5_io_outs_up[33] ;
 wire \ces_2_5_io_outs_up[34] ;
 wire \ces_2_5_io_outs_up[35] ;
 wire \ces_2_5_io_outs_up[36] ;
 wire \ces_2_5_io_outs_up[37] ;
 wire \ces_2_5_io_outs_up[38] ;
 wire \ces_2_5_io_outs_up[39] ;
 wire \ces_2_5_io_outs_up[3] ;
 wire \ces_2_5_io_outs_up[40] ;
 wire \ces_2_5_io_outs_up[41] ;
 wire \ces_2_5_io_outs_up[42] ;
 wire \ces_2_5_io_outs_up[43] ;
 wire \ces_2_5_io_outs_up[44] ;
 wire \ces_2_5_io_outs_up[45] ;
 wire \ces_2_5_io_outs_up[46] ;
 wire \ces_2_5_io_outs_up[47] ;
 wire \ces_2_5_io_outs_up[48] ;
 wire \ces_2_5_io_outs_up[49] ;
 wire \ces_2_5_io_outs_up[4] ;
 wire \ces_2_5_io_outs_up[50] ;
 wire \ces_2_5_io_outs_up[51] ;
 wire \ces_2_5_io_outs_up[52] ;
 wire \ces_2_5_io_outs_up[53] ;
 wire \ces_2_5_io_outs_up[54] ;
 wire \ces_2_5_io_outs_up[55] ;
 wire \ces_2_5_io_outs_up[56] ;
 wire \ces_2_5_io_outs_up[57] ;
 wire \ces_2_5_io_outs_up[58] ;
 wire \ces_2_5_io_outs_up[59] ;
 wire \ces_2_5_io_outs_up[5] ;
 wire \ces_2_5_io_outs_up[60] ;
 wire \ces_2_5_io_outs_up[61] ;
 wire \ces_2_5_io_outs_up[62] ;
 wire \ces_2_5_io_outs_up[63] ;
 wire \ces_2_5_io_outs_up[6] ;
 wire \ces_2_5_io_outs_up[7] ;
 wire \ces_2_5_io_outs_up[8] ;
 wire \ces_2_5_io_outs_up[9] ;
 wire \ces_2_6_io_ins_down[0] ;
 wire \ces_2_6_io_ins_down[10] ;
 wire \ces_2_6_io_ins_down[11] ;
 wire \ces_2_6_io_ins_down[12] ;
 wire \ces_2_6_io_ins_down[13] ;
 wire \ces_2_6_io_ins_down[14] ;
 wire \ces_2_6_io_ins_down[15] ;
 wire \ces_2_6_io_ins_down[16] ;
 wire \ces_2_6_io_ins_down[17] ;
 wire \ces_2_6_io_ins_down[18] ;
 wire \ces_2_6_io_ins_down[19] ;
 wire \ces_2_6_io_ins_down[1] ;
 wire \ces_2_6_io_ins_down[20] ;
 wire \ces_2_6_io_ins_down[21] ;
 wire \ces_2_6_io_ins_down[22] ;
 wire \ces_2_6_io_ins_down[23] ;
 wire \ces_2_6_io_ins_down[24] ;
 wire \ces_2_6_io_ins_down[25] ;
 wire \ces_2_6_io_ins_down[26] ;
 wire \ces_2_6_io_ins_down[27] ;
 wire \ces_2_6_io_ins_down[28] ;
 wire \ces_2_6_io_ins_down[29] ;
 wire \ces_2_6_io_ins_down[2] ;
 wire \ces_2_6_io_ins_down[30] ;
 wire \ces_2_6_io_ins_down[31] ;
 wire \ces_2_6_io_ins_down[32] ;
 wire \ces_2_6_io_ins_down[33] ;
 wire \ces_2_6_io_ins_down[34] ;
 wire \ces_2_6_io_ins_down[35] ;
 wire \ces_2_6_io_ins_down[36] ;
 wire \ces_2_6_io_ins_down[37] ;
 wire \ces_2_6_io_ins_down[38] ;
 wire \ces_2_6_io_ins_down[39] ;
 wire \ces_2_6_io_ins_down[3] ;
 wire \ces_2_6_io_ins_down[40] ;
 wire \ces_2_6_io_ins_down[41] ;
 wire \ces_2_6_io_ins_down[42] ;
 wire \ces_2_6_io_ins_down[43] ;
 wire \ces_2_6_io_ins_down[44] ;
 wire \ces_2_6_io_ins_down[45] ;
 wire \ces_2_6_io_ins_down[46] ;
 wire \ces_2_6_io_ins_down[47] ;
 wire \ces_2_6_io_ins_down[48] ;
 wire \ces_2_6_io_ins_down[49] ;
 wire \ces_2_6_io_ins_down[4] ;
 wire \ces_2_6_io_ins_down[50] ;
 wire \ces_2_6_io_ins_down[51] ;
 wire \ces_2_6_io_ins_down[52] ;
 wire \ces_2_6_io_ins_down[53] ;
 wire \ces_2_6_io_ins_down[54] ;
 wire \ces_2_6_io_ins_down[55] ;
 wire \ces_2_6_io_ins_down[56] ;
 wire \ces_2_6_io_ins_down[57] ;
 wire \ces_2_6_io_ins_down[58] ;
 wire \ces_2_6_io_ins_down[59] ;
 wire \ces_2_6_io_ins_down[5] ;
 wire \ces_2_6_io_ins_down[60] ;
 wire \ces_2_6_io_ins_down[61] ;
 wire \ces_2_6_io_ins_down[62] ;
 wire \ces_2_6_io_ins_down[63] ;
 wire \ces_2_6_io_ins_down[6] ;
 wire \ces_2_6_io_ins_down[7] ;
 wire \ces_2_6_io_ins_down[8] ;
 wire \ces_2_6_io_ins_down[9] ;
 wire \ces_2_6_io_ins_left[0] ;
 wire \ces_2_6_io_ins_left[10] ;
 wire \ces_2_6_io_ins_left[11] ;
 wire \ces_2_6_io_ins_left[12] ;
 wire \ces_2_6_io_ins_left[13] ;
 wire \ces_2_6_io_ins_left[14] ;
 wire \ces_2_6_io_ins_left[15] ;
 wire \ces_2_6_io_ins_left[16] ;
 wire \ces_2_6_io_ins_left[17] ;
 wire \ces_2_6_io_ins_left[18] ;
 wire \ces_2_6_io_ins_left[19] ;
 wire \ces_2_6_io_ins_left[1] ;
 wire \ces_2_6_io_ins_left[20] ;
 wire \ces_2_6_io_ins_left[21] ;
 wire \ces_2_6_io_ins_left[22] ;
 wire \ces_2_6_io_ins_left[23] ;
 wire \ces_2_6_io_ins_left[24] ;
 wire \ces_2_6_io_ins_left[25] ;
 wire \ces_2_6_io_ins_left[26] ;
 wire \ces_2_6_io_ins_left[27] ;
 wire \ces_2_6_io_ins_left[28] ;
 wire \ces_2_6_io_ins_left[29] ;
 wire \ces_2_6_io_ins_left[2] ;
 wire \ces_2_6_io_ins_left[30] ;
 wire \ces_2_6_io_ins_left[31] ;
 wire \ces_2_6_io_ins_left[32] ;
 wire \ces_2_6_io_ins_left[33] ;
 wire \ces_2_6_io_ins_left[34] ;
 wire \ces_2_6_io_ins_left[35] ;
 wire \ces_2_6_io_ins_left[36] ;
 wire \ces_2_6_io_ins_left[37] ;
 wire \ces_2_6_io_ins_left[38] ;
 wire \ces_2_6_io_ins_left[39] ;
 wire \ces_2_6_io_ins_left[3] ;
 wire \ces_2_6_io_ins_left[40] ;
 wire \ces_2_6_io_ins_left[41] ;
 wire \ces_2_6_io_ins_left[42] ;
 wire \ces_2_6_io_ins_left[43] ;
 wire \ces_2_6_io_ins_left[44] ;
 wire \ces_2_6_io_ins_left[45] ;
 wire \ces_2_6_io_ins_left[46] ;
 wire \ces_2_6_io_ins_left[47] ;
 wire \ces_2_6_io_ins_left[48] ;
 wire \ces_2_6_io_ins_left[49] ;
 wire \ces_2_6_io_ins_left[4] ;
 wire \ces_2_6_io_ins_left[50] ;
 wire \ces_2_6_io_ins_left[51] ;
 wire \ces_2_6_io_ins_left[52] ;
 wire \ces_2_6_io_ins_left[53] ;
 wire \ces_2_6_io_ins_left[54] ;
 wire \ces_2_6_io_ins_left[55] ;
 wire \ces_2_6_io_ins_left[56] ;
 wire \ces_2_6_io_ins_left[57] ;
 wire \ces_2_6_io_ins_left[58] ;
 wire \ces_2_6_io_ins_left[59] ;
 wire \ces_2_6_io_ins_left[5] ;
 wire \ces_2_6_io_ins_left[60] ;
 wire \ces_2_6_io_ins_left[61] ;
 wire \ces_2_6_io_ins_left[62] ;
 wire \ces_2_6_io_ins_left[63] ;
 wire \ces_2_6_io_ins_left[6] ;
 wire \ces_2_6_io_ins_left[7] ;
 wire \ces_2_6_io_ins_left[8] ;
 wire \ces_2_6_io_ins_left[9] ;
 wire ces_2_6_io_lsbOuts_0;
 wire ces_2_6_io_lsbOuts_1;
 wire ces_2_6_io_lsbOuts_2;
 wire ces_2_6_io_lsbOuts_3;
 wire ces_2_6_io_lsbOuts_4;
 wire ces_2_6_io_lsbOuts_5;
 wire ces_2_6_io_lsbOuts_6;
 wire ces_2_6_io_lsbOuts_7;
 wire \ces_2_6_io_outs_right[0] ;
 wire \ces_2_6_io_outs_right[10] ;
 wire \ces_2_6_io_outs_right[11] ;
 wire \ces_2_6_io_outs_right[12] ;
 wire \ces_2_6_io_outs_right[13] ;
 wire \ces_2_6_io_outs_right[14] ;
 wire \ces_2_6_io_outs_right[15] ;
 wire \ces_2_6_io_outs_right[16] ;
 wire \ces_2_6_io_outs_right[17] ;
 wire \ces_2_6_io_outs_right[18] ;
 wire \ces_2_6_io_outs_right[19] ;
 wire \ces_2_6_io_outs_right[1] ;
 wire \ces_2_6_io_outs_right[20] ;
 wire \ces_2_6_io_outs_right[21] ;
 wire \ces_2_6_io_outs_right[22] ;
 wire \ces_2_6_io_outs_right[23] ;
 wire \ces_2_6_io_outs_right[24] ;
 wire \ces_2_6_io_outs_right[25] ;
 wire \ces_2_6_io_outs_right[26] ;
 wire \ces_2_6_io_outs_right[27] ;
 wire \ces_2_6_io_outs_right[28] ;
 wire \ces_2_6_io_outs_right[29] ;
 wire \ces_2_6_io_outs_right[2] ;
 wire \ces_2_6_io_outs_right[30] ;
 wire \ces_2_6_io_outs_right[31] ;
 wire \ces_2_6_io_outs_right[32] ;
 wire \ces_2_6_io_outs_right[33] ;
 wire \ces_2_6_io_outs_right[34] ;
 wire \ces_2_6_io_outs_right[35] ;
 wire \ces_2_6_io_outs_right[36] ;
 wire \ces_2_6_io_outs_right[37] ;
 wire \ces_2_6_io_outs_right[38] ;
 wire \ces_2_6_io_outs_right[39] ;
 wire \ces_2_6_io_outs_right[3] ;
 wire \ces_2_6_io_outs_right[40] ;
 wire \ces_2_6_io_outs_right[41] ;
 wire \ces_2_6_io_outs_right[42] ;
 wire \ces_2_6_io_outs_right[43] ;
 wire \ces_2_6_io_outs_right[44] ;
 wire \ces_2_6_io_outs_right[45] ;
 wire \ces_2_6_io_outs_right[46] ;
 wire \ces_2_6_io_outs_right[47] ;
 wire \ces_2_6_io_outs_right[48] ;
 wire \ces_2_6_io_outs_right[49] ;
 wire \ces_2_6_io_outs_right[4] ;
 wire \ces_2_6_io_outs_right[50] ;
 wire \ces_2_6_io_outs_right[51] ;
 wire \ces_2_6_io_outs_right[52] ;
 wire \ces_2_6_io_outs_right[53] ;
 wire \ces_2_6_io_outs_right[54] ;
 wire \ces_2_6_io_outs_right[55] ;
 wire \ces_2_6_io_outs_right[56] ;
 wire \ces_2_6_io_outs_right[57] ;
 wire \ces_2_6_io_outs_right[58] ;
 wire \ces_2_6_io_outs_right[59] ;
 wire \ces_2_6_io_outs_right[5] ;
 wire \ces_2_6_io_outs_right[60] ;
 wire \ces_2_6_io_outs_right[61] ;
 wire \ces_2_6_io_outs_right[62] ;
 wire \ces_2_6_io_outs_right[63] ;
 wire \ces_2_6_io_outs_right[6] ;
 wire \ces_2_6_io_outs_right[7] ;
 wire \ces_2_6_io_outs_right[8] ;
 wire \ces_2_6_io_outs_right[9] ;
 wire \ces_2_6_io_outs_up[0] ;
 wire \ces_2_6_io_outs_up[10] ;
 wire \ces_2_6_io_outs_up[11] ;
 wire \ces_2_6_io_outs_up[12] ;
 wire \ces_2_6_io_outs_up[13] ;
 wire \ces_2_6_io_outs_up[14] ;
 wire \ces_2_6_io_outs_up[15] ;
 wire \ces_2_6_io_outs_up[16] ;
 wire \ces_2_6_io_outs_up[17] ;
 wire \ces_2_6_io_outs_up[18] ;
 wire \ces_2_6_io_outs_up[19] ;
 wire \ces_2_6_io_outs_up[1] ;
 wire \ces_2_6_io_outs_up[20] ;
 wire \ces_2_6_io_outs_up[21] ;
 wire \ces_2_6_io_outs_up[22] ;
 wire \ces_2_6_io_outs_up[23] ;
 wire \ces_2_6_io_outs_up[24] ;
 wire \ces_2_6_io_outs_up[25] ;
 wire \ces_2_6_io_outs_up[26] ;
 wire \ces_2_6_io_outs_up[27] ;
 wire \ces_2_6_io_outs_up[28] ;
 wire \ces_2_6_io_outs_up[29] ;
 wire \ces_2_6_io_outs_up[2] ;
 wire \ces_2_6_io_outs_up[30] ;
 wire \ces_2_6_io_outs_up[31] ;
 wire \ces_2_6_io_outs_up[32] ;
 wire \ces_2_6_io_outs_up[33] ;
 wire \ces_2_6_io_outs_up[34] ;
 wire \ces_2_6_io_outs_up[35] ;
 wire \ces_2_6_io_outs_up[36] ;
 wire \ces_2_6_io_outs_up[37] ;
 wire \ces_2_6_io_outs_up[38] ;
 wire \ces_2_6_io_outs_up[39] ;
 wire \ces_2_6_io_outs_up[3] ;
 wire \ces_2_6_io_outs_up[40] ;
 wire \ces_2_6_io_outs_up[41] ;
 wire \ces_2_6_io_outs_up[42] ;
 wire \ces_2_6_io_outs_up[43] ;
 wire \ces_2_6_io_outs_up[44] ;
 wire \ces_2_6_io_outs_up[45] ;
 wire \ces_2_6_io_outs_up[46] ;
 wire \ces_2_6_io_outs_up[47] ;
 wire \ces_2_6_io_outs_up[48] ;
 wire \ces_2_6_io_outs_up[49] ;
 wire \ces_2_6_io_outs_up[4] ;
 wire \ces_2_6_io_outs_up[50] ;
 wire \ces_2_6_io_outs_up[51] ;
 wire \ces_2_6_io_outs_up[52] ;
 wire \ces_2_6_io_outs_up[53] ;
 wire \ces_2_6_io_outs_up[54] ;
 wire \ces_2_6_io_outs_up[55] ;
 wire \ces_2_6_io_outs_up[56] ;
 wire \ces_2_6_io_outs_up[57] ;
 wire \ces_2_6_io_outs_up[58] ;
 wire \ces_2_6_io_outs_up[59] ;
 wire \ces_2_6_io_outs_up[5] ;
 wire \ces_2_6_io_outs_up[60] ;
 wire \ces_2_6_io_outs_up[61] ;
 wire \ces_2_6_io_outs_up[62] ;
 wire \ces_2_6_io_outs_up[63] ;
 wire \ces_2_6_io_outs_up[6] ;
 wire \ces_2_6_io_outs_up[7] ;
 wire \ces_2_6_io_outs_up[8] ;
 wire \ces_2_6_io_outs_up[9] ;
 wire \ces_2_7_io_ins_down[0] ;
 wire \ces_2_7_io_ins_down[10] ;
 wire \ces_2_7_io_ins_down[11] ;
 wire \ces_2_7_io_ins_down[12] ;
 wire \ces_2_7_io_ins_down[13] ;
 wire \ces_2_7_io_ins_down[14] ;
 wire \ces_2_7_io_ins_down[15] ;
 wire \ces_2_7_io_ins_down[16] ;
 wire \ces_2_7_io_ins_down[17] ;
 wire \ces_2_7_io_ins_down[18] ;
 wire \ces_2_7_io_ins_down[19] ;
 wire \ces_2_7_io_ins_down[1] ;
 wire \ces_2_7_io_ins_down[20] ;
 wire \ces_2_7_io_ins_down[21] ;
 wire \ces_2_7_io_ins_down[22] ;
 wire \ces_2_7_io_ins_down[23] ;
 wire \ces_2_7_io_ins_down[24] ;
 wire \ces_2_7_io_ins_down[25] ;
 wire \ces_2_7_io_ins_down[26] ;
 wire \ces_2_7_io_ins_down[27] ;
 wire \ces_2_7_io_ins_down[28] ;
 wire \ces_2_7_io_ins_down[29] ;
 wire \ces_2_7_io_ins_down[2] ;
 wire \ces_2_7_io_ins_down[30] ;
 wire \ces_2_7_io_ins_down[31] ;
 wire \ces_2_7_io_ins_down[32] ;
 wire \ces_2_7_io_ins_down[33] ;
 wire \ces_2_7_io_ins_down[34] ;
 wire \ces_2_7_io_ins_down[35] ;
 wire \ces_2_7_io_ins_down[36] ;
 wire \ces_2_7_io_ins_down[37] ;
 wire \ces_2_7_io_ins_down[38] ;
 wire \ces_2_7_io_ins_down[39] ;
 wire \ces_2_7_io_ins_down[3] ;
 wire \ces_2_7_io_ins_down[40] ;
 wire \ces_2_7_io_ins_down[41] ;
 wire \ces_2_7_io_ins_down[42] ;
 wire \ces_2_7_io_ins_down[43] ;
 wire \ces_2_7_io_ins_down[44] ;
 wire \ces_2_7_io_ins_down[45] ;
 wire \ces_2_7_io_ins_down[46] ;
 wire \ces_2_7_io_ins_down[47] ;
 wire \ces_2_7_io_ins_down[48] ;
 wire \ces_2_7_io_ins_down[49] ;
 wire \ces_2_7_io_ins_down[4] ;
 wire \ces_2_7_io_ins_down[50] ;
 wire \ces_2_7_io_ins_down[51] ;
 wire \ces_2_7_io_ins_down[52] ;
 wire \ces_2_7_io_ins_down[53] ;
 wire \ces_2_7_io_ins_down[54] ;
 wire \ces_2_7_io_ins_down[55] ;
 wire \ces_2_7_io_ins_down[56] ;
 wire \ces_2_7_io_ins_down[57] ;
 wire \ces_2_7_io_ins_down[58] ;
 wire \ces_2_7_io_ins_down[59] ;
 wire \ces_2_7_io_ins_down[5] ;
 wire \ces_2_7_io_ins_down[60] ;
 wire \ces_2_7_io_ins_down[61] ;
 wire \ces_2_7_io_ins_down[62] ;
 wire \ces_2_7_io_ins_down[63] ;
 wire \ces_2_7_io_ins_down[6] ;
 wire \ces_2_7_io_ins_down[7] ;
 wire \ces_2_7_io_ins_down[8] ;
 wire \ces_2_7_io_ins_down[9] ;
 wire ces_2_7_io_lsbOuts_0;
 wire ces_2_7_io_lsbOuts_1;
 wire ces_2_7_io_lsbOuts_2;
 wire ces_2_7_io_lsbOuts_3;
 wire ces_2_7_io_lsbOuts_4;
 wire ces_2_7_io_lsbOuts_5;
 wire ces_2_7_io_lsbOuts_6;
 wire ces_2_7_io_lsbOuts_7;
 wire \ces_2_7_io_outs_up[0] ;
 wire \ces_2_7_io_outs_up[10] ;
 wire \ces_2_7_io_outs_up[11] ;
 wire \ces_2_7_io_outs_up[12] ;
 wire \ces_2_7_io_outs_up[13] ;
 wire \ces_2_7_io_outs_up[14] ;
 wire \ces_2_7_io_outs_up[15] ;
 wire \ces_2_7_io_outs_up[16] ;
 wire \ces_2_7_io_outs_up[17] ;
 wire \ces_2_7_io_outs_up[18] ;
 wire \ces_2_7_io_outs_up[19] ;
 wire \ces_2_7_io_outs_up[1] ;
 wire \ces_2_7_io_outs_up[20] ;
 wire \ces_2_7_io_outs_up[21] ;
 wire \ces_2_7_io_outs_up[22] ;
 wire \ces_2_7_io_outs_up[23] ;
 wire \ces_2_7_io_outs_up[24] ;
 wire \ces_2_7_io_outs_up[25] ;
 wire \ces_2_7_io_outs_up[26] ;
 wire \ces_2_7_io_outs_up[27] ;
 wire \ces_2_7_io_outs_up[28] ;
 wire \ces_2_7_io_outs_up[29] ;
 wire \ces_2_7_io_outs_up[2] ;
 wire \ces_2_7_io_outs_up[30] ;
 wire \ces_2_7_io_outs_up[31] ;
 wire \ces_2_7_io_outs_up[32] ;
 wire \ces_2_7_io_outs_up[33] ;
 wire \ces_2_7_io_outs_up[34] ;
 wire \ces_2_7_io_outs_up[35] ;
 wire \ces_2_7_io_outs_up[36] ;
 wire \ces_2_7_io_outs_up[37] ;
 wire \ces_2_7_io_outs_up[38] ;
 wire \ces_2_7_io_outs_up[39] ;
 wire \ces_2_7_io_outs_up[3] ;
 wire \ces_2_7_io_outs_up[40] ;
 wire \ces_2_7_io_outs_up[41] ;
 wire \ces_2_7_io_outs_up[42] ;
 wire \ces_2_7_io_outs_up[43] ;
 wire \ces_2_7_io_outs_up[44] ;
 wire \ces_2_7_io_outs_up[45] ;
 wire \ces_2_7_io_outs_up[46] ;
 wire \ces_2_7_io_outs_up[47] ;
 wire \ces_2_7_io_outs_up[48] ;
 wire \ces_2_7_io_outs_up[49] ;
 wire \ces_2_7_io_outs_up[4] ;
 wire \ces_2_7_io_outs_up[50] ;
 wire \ces_2_7_io_outs_up[51] ;
 wire \ces_2_7_io_outs_up[52] ;
 wire \ces_2_7_io_outs_up[53] ;
 wire \ces_2_7_io_outs_up[54] ;
 wire \ces_2_7_io_outs_up[55] ;
 wire \ces_2_7_io_outs_up[56] ;
 wire \ces_2_7_io_outs_up[57] ;
 wire \ces_2_7_io_outs_up[58] ;
 wire \ces_2_7_io_outs_up[59] ;
 wire \ces_2_7_io_outs_up[5] ;
 wire \ces_2_7_io_outs_up[60] ;
 wire \ces_2_7_io_outs_up[61] ;
 wire \ces_2_7_io_outs_up[62] ;
 wire \ces_2_7_io_outs_up[63] ;
 wire \ces_2_7_io_outs_up[6] ;
 wire \ces_2_7_io_outs_up[7] ;
 wire \ces_2_7_io_outs_up[8] ;
 wire \ces_2_7_io_outs_up[9] ;
 wire \ces_3_0_io_ins_down[0] ;
 wire \ces_3_0_io_ins_down[10] ;
 wire \ces_3_0_io_ins_down[11] ;
 wire \ces_3_0_io_ins_down[12] ;
 wire \ces_3_0_io_ins_down[13] ;
 wire \ces_3_0_io_ins_down[14] ;
 wire \ces_3_0_io_ins_down[15] ;
 wire \ces_3_0_io_ins_down[16] ;
 wire \ces_3_0_io_ins_down[17] ;
 wire \ces_3_0_io_ins_down[18] ;
 wire \ces_3_0_io_ins_down[19] ;
 wire \ces_3_0_io_ins_down[1] ;
 wire \ces_3_0_io_ins_down[20] ;
 wire \ces_3_0_io_ins_down[21] ;
 wire \ces_3_0_io_ins_down[22] ;
 wire \ces_3_0_io_ins_down[23] ;
 wire \ces_3_0_io_ins_down[24] ;
 wire \ces_3_0_io_ins_down[25] ;
 wire \ces_3_0_io_ins_down[26] ;
 wire \ces_3_0_io_ins_down[27] ;
 wire \ces_3_0_io_ins_down[28] ;
 wire \ces_3_0_io_ins_down[29] ;
 wire \ces_3_0_io_ins_down[2] ;
 wire \ces_3_0_io_ins_down[30] ;
 wire \ces_3_0_io_ins_down[31] ;
 wire \ces_3_0_io_ins_down[32] ;
 wire \ces_3_0_io_ins_down[33] ;
 wire \ces_3_0_io_ins_down[34] ;
 wire \ces_3_0_io_ins_down[35] ;
 wire \ces_3_0_io_ins_down[36] ;
 wire \ces_3_0_io_ins_down[37] ;
 wire \ces_3_0_io_ins_down[38] ;
 wire \ces_3_0_io_ins_down[39] ;
 wire \ces_3_0_io_ins_down[3] ;
 wire \ces_3_0_io_ins_down[40] ;
 wire \ces_3_0_io_ins_down[41] ;
 wire \ces_3_0_io_ins_down[42] ;
 wire \ces_3_0_io_ins_down[43] ;
 wire \ces_3_0_io_ins_down[44] ;
 wire \ces_3_0_io_ins_down[45] ;
 wire \ces_3_0_io_ins_down[46] ;
 wire \ces_3_0_io_ins_down[47] ;
 wire \ces_3_0_io_ins_down[48] ;
 wire \ces_3_0_io_ins_down[49] ;
 wire \ces_3_0_io_ins_down[4] ;
 wire \ces_3_0_io_ins_down[50] ;
 wire \ces_3_0_io_ins_down[51] ;
 wire \ces_3_0_io_ins_down[52] ;
 wire \ces_3_0_io_ins_down[53] ;
 wire \ces_3_0_io_ins_down[54] ;
 wire \ces_3_0_io_ins_down[55] ;
 wire \ces_3_0_io_ins_down[56] ;
 wire \ces_3_0_io_ins_down[57] ;
 wire \ces_3_0_io_ins_down[58] ;
 wire \ces_3_0_io_ins_down[59] ;
 wire \ces_3_0_io_ins_down[5] ;
 wire \ces_3_0_io_ins_down[60] ;
 wire \ces_3_0_io_ins_down[61] ;
 wire \ces_3_0_io_ins_down[62] ;
 wire \ces_3_0_io_ins_down[63] ;
 wire \ces_3_0_io_ins_down[6] ;
 wire \ces_3_0_io_ins_down[7] ;
 wire \ces_3_0_io_ins_down[8] ;
 wire \ces_3_0_io_ins_down[9] ;
 wire \ces_3_0_io_ins_left[0] ;
 wire \ces_3_0_io_ins_left[10] ;
 wire \ces_3_0_io_ins_left[11] ;
 wire \ces_3_0_io_ins_left[12] ;
 wire \ces_3_0_io_ins_left[13] ;
 wire \ces_3_0_io_ins_left[14] ;
 wire \ces_3_0_io_ins_left[15] ;
 wire \ces_3_0_io_ins_left[16] ;
 wire \ces_3_0_io_ins_left[17] ;
 wire \ces_3_0_io_ins_left[18] ;
 wire \ces_3_0_io_ins_left[19] ;
 wire \ces_3_0_io_ins_left[1] ;
 wire \ces_3_0_io_ins_left[20] ;
 wire \ces_3_0_io_ins_left[21] ;
 wire \ces_3_0_io_ins_left[22] ;
 wire \ces_3_0_io_ins_left[23] ;
 wire \ces_3_0_io_ins_left[24] ;
 wire \ces_3_0_io_ins_left[25] ;
 wire \ces_3_0_io_ins_left[26] ;
 wire \ces_3_0_io_ins_left[27] ;
 wire \ces_3_0_io_ins_left[28] ;
 wire \ces_3_0_io_ins_left[29] ;
 wire \ces_3_0_io_ins_left[2] ;
 wire \ces_3_0_io_ins_left[30] ;
 wire \ces_3_0_io_ins_left[31] ;
 wire \ces_3_0_io_ins_left[32] ;
 wire \ces_3_0_io_ins_left[33] ;
 wire \ces_3_0_io_ins_left[34] ;
 wire \ces_3_0_io_ins_left[35] ;
 wire \ces_3_0_io_ins_left[36] ;
 wire \ces_3_0_io_ins_left[37] ;
 wire \ces_3_0_io_ins_left[38] ;
 wire \ces_3_0_io_ins_left[39] ;
 wire \ces_3_0_io_ins_left[3] ;
 wire \ces_3_0_io_ins_left[40] ;
 wire \ces_3_0_io_ins_left[41] ;
 wire \ces_3_0_io_ins_left[42] ;
 wire \ces_3_0_io_ins_left[43] ;
 wire \ces_3_0_io_ins_left[44] ;
 wire \ces_3_0_io_ins_left[45] ;
 wire \ces_3_0_io_ins_left[46] ;
 wire \ces_3_0_io_ins_left[47] ;
 wire \ces_3_0_io_ins_left[48] ;
 wire \ces_3_0_io_ins_left[49] ;
 wire \ces_3_0_io_ins_left[4] ;
 wire \ces_3_0_io_ins_left[50] ;
 wire \ces_3_0_io_ins_left[51] ;
 wire \ces_3_0_io_ins_left[52] ;
 wire \ces_3_0_io_ins_left[53] ;
 wire \ces_3_0_io_ins_left[54] ;
 wire \ces_3_0_io_ins_left[55] ;
 wire \ces_3_0_io_ins_left[56] ;
 wire \ces_3_0_io_ins_left[57] ;
 wire \ces_3_0_io_ins_left[58] ;
 wire \ces_3_0_io_ins_left[59] ;
 wire \ces_3_0_io_ins_left[5] ;
 wire \ces_3_0_io_ins_left[60] ;
 wire \ces_3_0_io_ins_left[61] ;
 wire \ces_3_0_io_ins_left[62] ;
 wire \ces_3_0_io_ins_left[63] ;
 wire \ces_3_0_io_ins_left[6] ;
 wire \ces_3_0_io_ins_left[7] ;
 wire \ces_3_0_io_ins_left[8] ;
 wire \ces_3_0_io_ins_left[9] ;
 wire ces_3_0_io_lsbOuts_0;
 wire ces_3_0_io_lsbOuts_1;
 wire ces_3_0_io_lsbOuts_2;
 wire ces_3_0_io_lsbOuts_3;
 wire ces_3_0_io_lsbOuts_4;
 wire ces_3_0_io_lsbOuts_5;
 wire ces_3_0_io_lsbOuts_6;
 wire ces_3_0_io_lsbOuts_7;
 wire \ces_3_0_io_outs_right[0] ;
 wire \ces_3_0_io_outs_right[10] ;
 wire \ces_3_0_io_outs_right[11] ;
 wire \ces_3_0_io_outs_right[12] ;
 wire \ces_3_0_io_outs_right[13] ;
 wire \ces_3_0_io_outs_right[14] ;
 wire \ces_3_0_io_outs_right[15] ;
 wire \ces_3_0_io_outs_right[16] ;
 wire \ces_3_0_io_outs_right[17] ;
 wire \ces_3_0_io_outs_right[18] ;
 wire \ces_3_0_io_outs_right[19] ;
 wire \ces_3_0_io_outs_right[1] ;
 wire \ces_3_0_io_outs_right[20] ;
 wire \ces_3_0_io_outs_right[21] ;
 wire \ces_3_0_io_outs_right[22] ;
 wire \ces_3_0_io_outs_right[23] ;
 wire \ces_3_0_io_outs_right[24] ;
 wire \ces_3_0_io_outs_right[25] ;
 wire \ces_3_0_io_outs_right[26] ;
 wire \ces_3_0_io_outs_right[27] ;
 wire \ces_3_0_io_outs_right[28] ;
 wire \ces_3_0_io_outs_right[29] ;
 wire \ces_3_0_io_outs_right[2] ;
 wire \ces_3_0_io_outs_right[30] ;
 wire \ces_3_0_io_outs_right[31] ;
 wire \ces_3_0_io_outs_right[32] ;
 wire \ces_3_0_io_outs_right[33] ;
 wire \ces_3_0_io_outs_right[34] ;
 wire \ces_3_0_io_outs_right[35] ;
 wire \ces_3_0_io_outs_right[36] ;
 wire \ces_3_0_io_outs_right[37] ;
 wire \ces_3_0_io_outs_right[38] ;
 wire \ces_3_0_io_outs_right[39] ;
 wire \ces_3_0_io_outs_right[3] ;
 wire \ces_3_0_io_outs_right[40] ;
 wire \ces_3_0_io_outs_right[41] ;
 wire \ces_3_0_io_outs_right[42] ;
 wire \ces_3_0_io_outs_right[43] ;
 wire \ces_3_0_io_outs_right[44] ;
 wire \ces_3_0_io_outs_right[45] ;
 wire \ces_3_0_io_outs_right[46] ;
 wire \ces_3_0_io_outs_right[47] ;
 wire \ces_3_0_io_outs_right[48] ;
 wire \ces_3_0_io_outs_right[49] ;
 wire \ces_3_0_io_outs_right[4] ;
 wire \ces_3_0_io_outs_right[50] ;
 wire \ces_3_0_io_outs_right[51] ;
 wire \ces_3_0_io_outs_right[52] ;
 wire \ces_3_0_io_outs_right[53] ;
 wire \ces_3_0_io_outs_right[54] ;
 wire \ces_3_0_io_outs_right[55] ;
 wire \ces_3_0_io_outs_right[56] ;
 wire \ces_3_0_io_outs_right[57] ;
 wire \ces_3_0_io_outs_right[58] ;
 wire \ces_3_0_io_outs_right[59] ;
 wire \ces_3_0_io_outs_right[5] ;
 wire \ces_3_0_io_outs_right[60] ;
 wire \ces_3_0_io_outs_right[61] ;
 wire \ces_3_0_io_outs_right[62] ;
 wire \ces_3_0_io_outs_right[63] ;
 wire \ces_3_0_io_outs_right[6] ;
 wire \ces_3_0_io_outs_right[7] ;
 wire \ces_3_0_io_outs_right[8] ;
 wire \ces_3_0_io_outs_right[9] ;
 wire \ces_3_0_io_outs_up[0] ;
 wire \ces_3_0_io_outs_up[10] ;
 wire \ces_3_0_io_outs_up[11] ;
 wire \ces_3_0_io_outs_up[12] ;
 wire \ces_3_0_io_outs_up[13] ;
 wire \ces_3_0_io_outs_up[14] ;
 wire \ces_3_0_io_outs_up[15] ;
 wire \ces_3_0_io_outs_up[16] ;
 wire \ces_3_0_io_outs_up[17] ;
 wire \ces_3_0_io_outs_up[18] ;
 wire \ces_3_0_io_outs_up[19] ;
 wire \ces_3_0_io_outs_up[1] ;
 wire \ces_3_0_io_outs_up[20] ;
 wire \ces_3_0_io_outs_up[21] ;
 wire \ces_3_0_io_outs_up[22] ;
 wire \ces_3_0_io_outs_up[23] ;
 wire \ces_3_0_io_outs_up[24] ;
 wire \ces_3_0_io_outs_up[25] ;
 wire \ces_3_0_io_outs_up[26] ;
 wire \ces_3_0_io_outs_up[27] ;
 wire \ces_3_0_io_outs_up[28] ;
 wire \ces_3_0_io_outs_up[29] ;
 wire \ces_3_0_io_outs_up[2] ;
 wire \ces_3_0_io_outs_up[30] ;
 wire \ces_3_0_io_outs_up[31] ;
 wire \ces_3_0_io_outs_up[32] ;
 wire \ces_3_0_io_outs_up[33] ;
 wire \ces_3_0_io_outs_up[34] ;
 wire \ces_3_0_io_outs_up[35] ;
 wire \ces_3_0_io_outs_up[36] ;
 wire \ces_3_0_io_outs_up[37] ;
 wire \ces_3_0_io_outs_up[38] ;
 wire \ces_3_0_io_outs_up[39] ;
 wire \ces_3_0_io_outs_up[3] ;
 wire \ces_3_0_io_outs_up[40] ;
 wire \ces_3_0_io_outs_up[41] ;
 wire \ces_3_0_io_outs_up[42] ;
 wire \ces_3_0_io_outs_up[43] ;
 wire \ces_3_0_io_outs_up[44] ;
 wire \ces_3_0_io_outs_up[45] ;
 wire \ces_3_0_io_outs_up[46] ;
 wire \ces_3_0_io_outs_up[47] ;
 wire \ces_3_0_io_outs_up[48] ;
 wire \ces_3_0_io_outs_up[49] ;
 wire \ces_3_0_io_outs_up[4] ;
 wire \ces_3_0_io_outs_up[50] ;
 wire \ces_3_0_io_outs_up[51] ;
 wire \ces_3_0_io_outs_up[52] ;
 wire \ces_3_0_io_outs_up[53] ;
 wire \ces_3_0_io_outs_up[54] ;
 wire \ces_3_0_io_outs_up[55] ;
 wire \ces_3_0_io_outs_up[56] ;
 wire \ces_3_0_io_outs_up[57] ;
 wire \ces_3_0_io_outs_up[58] ;
 wire \ces_3_0_io_outs_up[59] ;
 wire \ces_3_0_io_outs_up[5] ;
 wire \ces_3_0_io_outs_up[60] ;
 wire \ces_3_0_io_outs_up[61] ;
 wire \ces_3_0_io_outs_up[62] ;
 wire \ces_3_0_io_outs_up[63] ;
 wire \ces_3_0_io_outs_up[6] ;
 wire \ces_3_0_io_outs_up[7] ;
 wire \ces_3_0_io_outs_up[8] ;
 wire \ces_3_0_io_outs_up[9] ;
 wire \ces_3_1_io_ins_down[0] ;
 wire \ces_3_1_io_ins_down[10] ;
 wire \ces_3_1_io_ins_down[11] ;
 wire \ces_3_1_io_ins_down[12] ;
 wire \ces_3_1_io_ins_down[13] ;
 wire \ces_3_1_io_ins_down[14] ;
 wire \ces_3_1_io_ins_down[15] ;
 wire \ces_3_1_io_ins_down[16] ;
 wire \ces_3_1_io_ins_down[17] ;
 wire \ces_3_1_io_ins_down[18] ;
 wire \ces_3_1_io_ins_down[19] ;
 wire \ces_3_1_io_ins_down[1] ;
 wire \ces_3_1_io_ins_down[20] ;
 wire \ces_3_1_io_ins_down[21] ;
 wire \ces_3_1_io_ins_down[22] ;
 wire \ces_3_1_io_ins_down[23] ;
 wire \ces_3_1_io_ins_down[24] ;
 wire \ces_3_1_io_ins_down[25] ;
 wire \ces_3_1_io_ins_down[26] ;
 wire \ces_3_1_io_ins_down[27] ;
 wire \ces_3_1_io_ins_down[28] ;
 wire \ces_3_1_io_ins_down[29] ;
 wire \ces_3_1_io_ins_down[2] ;
 wire \ces_3_1_io_ins_down[30] ;
 wire \ces_3_1_io_ins_down[31] ;
 wire \ces_3_1_io_ins_down[32] ;
 wire \ces_3_1_io_ins_down[33] ;
 wire \ces_3_1_io_ins_down[34] ;
 wire \ces_3_1_io_ins_down[35] ;
 wire \ces_3_1_io_ins_down[36] ;
 wire \ces_3_1_io_ins_down[37] ;
 wire \ces_3_1_io_ins_down[38] ;
 wire \ces_3_1_io_ins_down[39] ;
 wire \ces_3_1_io_ins_down[3] ;
 wire \ces_3_1_io_ins_down[40] ;
 wire \ces_3_1_io_ins_down[41] ;
 wire \ces_3_1_io_ins_down[42] ;
 wire \ces_3_1_io_ins_down[43] ;
 wire \ces_3_1_io_ins_down[44] ;
 wire \ces_3_1_io_ins_down[45] ;
 wire \ces_3_1_io_ins_down[46] ;
 wire \ces_3_1_io_ins_down[47] ;
 wire \ces_3_1_io_ins_down[48] ;
 wire \ces_3_1_io_ins_down[49] ;
 wire \ces_3_1_io_ins_down[4] ;
 wire \ces_3_1_io_ins_down[50] ;
 wire \ces_3_1_io_ins_down[51] ;
 wire \ces_3_1_io_ins_down[52] ;
 wire \ces_3_1_io_ins_down[53] ;
 wire \ces_3_1_io_ins_down[54] ;
 wire \ces_3_1_io_ins_down[55] ;
 wire \ces_3_1_io_ins_down[56] ;
 wire \ces_3_1_io_ins_down[57] ;
 wire \ces_3_1_io_ins_down[58] ;
 wire \ces_3_1_io_ins_down[59] ;
 wire \ces_3_1_io_ins_down[5] ;
 wire \ces_3_1_io_ins_down[60] ;
 wire \ces_3_1_io_ins_down[61] ;
 wire \ces_3_1_io_ins_down[62] ;
 wire \ces_3_1_io_ins_down[63] ;
 wire \ces_3_1_io_ins_down[6] ;
 wire \ces_3_1_io_ins_down[7] ;
 wire \ces_3_1_io_ins_down[8] ;
 wire \ces_3_1_io_ins_down[9] ;
 wire \ces_3_1_io_ins_left[0] ;
 wire \ces_3_1_io_ins_left[10] ;
 wire \ces_3_1_io_ins_left[11] ;
 wire \ces_3_1_io_ins_left[12] ;
 wire \ces_3_1_io_ins_left[13] ;
 wire \ces_3_1_io_ins_left[14] ;
 wire \ces_3_1_io_ins_left[15] ;
 wire \ces_3_1_io_ins_left[16] ;
 wire \ces_3_1_io_ins_left[17] ;
 wire \ces_3_1_io_ins_left[18] ;
 wire \ces_3_1_io_ins_left[19] ;
 wire \ces_3_1_io_ins_left[1] ;
 wire \ces_3_1_io_ins_left[20] ;
 wire \ces_3_1_io_ins_left[21] ;
 wire \ces_3_1_io_ins_left[22] ;
 wire \ces_3_1_io_ins_left[23] ;
 wire \ces_3_1_io_ins_left[24] ;
 wire \ces_3_1_io_ins_left[25] ;
 wire \ces_3_1_io_ins_left[26] ;
 wire \ces_3_1_io_ins_left[27] ;
 wire \ces_3_1_io_ins_left[28] ;
 wire \ces_3_1_io_ins_left[29] ;
 wire \ces_3_1_io_ins_left[2] ;
 wire \ces_3_1_io_ins_left[30] ;
 wire \ces_3_1_io_ins_left[31] ;
 wire \ces_3_1_io_ins_left[32] ;
 wire \ces_3_1_io_ins_left[33] ;
 wire \ces_3_1_io_ins_left[34] ;
 wire \ces_3_1_io_ins_left[35] ;
 wire \ces_3_1_io_ins_left[36] ;
 wire \ces_3_1_io_ins_left[37] ;
 wire \ces_3_1_io_ins_left[38] ;
 wire \ces_3_1_io_ins_left[39] ;
 wire \ces_3_1_io_ins_left[3] ;
 wire \ces_3_1_io_ins_left[40] ;
 wire \ces_3_1_io_ins_left[41] ;
 wire \ces_3_1_io_ins_left[42] ;
 wire \ces_3_1_io_ins_left[43] ;
 wire \ces_3_1_io_ins_left[44] ;
 wire \ces_3_1_io_ins_left[45] ;
 wire \ces_3_1_io_ins_left[46] ;
 wire \ces_3_1_io_ins_left[47] ;
 wire \ces_3_1_io_ins_left[48] ;
 wire \ces_3_1_io_ins_left[49] ;
 wire \ces_3_1_io_ins_left[4] ;
 wire \ces_3_1_io_ins_left[50] ;
 wire \ces_3_1_io_ins_left[51] ;
 wire \ces_3_1_io_ins_left[52] ;
 wire \ces_3_1_io_ins_left[53] ;
 wire \ces_3_1_io_ins_left[54] ;
 wire \ces_3_1_io_ins_left[55] ;
 wire \ces_3_1_io_ins_left[56] ;
 wire \ces_3_1_io_ins_left[57] ;
 wire \ces_3_1_io_ins_left[58] ;
 wire \ces_3_1_io_ins_left[59] ;
 wire \ces_3_1_io_ins_left[5] ;
 wire \ces_3_1_io_ins_left[60] ;
 wire \ces_3_1_io_ins_left[61] ;
 wire \ces_3_1_io_ins_left[62] ;
 wire \ces_3_1_io_ins_left[63] ;
 wire \ces_3_1_io_ins_left[6] ;
 wire \ces_3_1_io_ins_left[7] ;
 wire \ces_3_1_io_ins_left[8] ;
 wire \ces_3_1_io_ins_left[9] ;
 wire ces_3_1_io_lsbOuts_0;
 wire ces_3_1_io_lsbOuts_1;
 wire ces_3_1_io_lsbOuts_2;
 wire ces_3_1_io_lsbOuts_3;
 wire ces_3_1_io_lsbOuts_4;
 wire ces_3_1_io_lsbOuts_5;
 wire ces_3_1_io_lsbOuts_6;
 wire ces_3_1_io_lsbOuts_7;
 wire \ces_3_1_io_outs_right[0] ;
 wire \ces_3_1_io_outs_right[10] ;
 wire \ces_3_1_io_outs_right[11] ;
 wire \ces_3_1_io_outs_right[12] ;
 wire \ces_3_1_io_outs_right[13] ;
 wire \ces_3_1_io_outs_right[14] ;
 wire \ces_3_1_io_outs_right[15] ;
 wire \ces_3_1_io_outs_right[16] ;
 wire \ces_3_1_io_outs_right[17] ;
 wire \ces_3_1_io_outs_right[18] ;
 wire \ces_3_1_io_outs_right[19] ;
 wire \ces_3_1_io_outs_right[1] ;
 wire \ces_3_1_io_outs_right[20] ;
 wire \ces_3_1_io_outs_right[21] ;
 wire \ces_3_1_io_outs_right[22] ;
 wire \ces_3_1_io_outs_right[23] ;
 wire \ces_3_1_io_outs_right[24] ;
 wire \ces_3_1_io_outs_right[25] ;
 wire \ces_3_1_io_outs_right[26] ;
 wire \ces_3_1_io_outs_right[27] ;
 wire \ces_3_1_io_outs_right[28] ;
 wire \ces_3_1_io_outs_right[29] ;
 wire \ces_3_1_io_outs_right[2] ;
 wire \ces_3_1_io_outs_right[30] ;
 wire \ces_3_1_io_outs_right[31] ;
 wire \ces_3_1_io_outs_right[32] ;
 wire \ces_3_1_io_outs_right[33] ;
 wire \ces_3_1_io_outs_right[34] ;
 wire \ces_3_1_io_outs_right[35] ;
 wire \ces_3_1_io_outs_right[36] ;
 wire \ces_3_1_io_outs_right[37] ;
 wire \ces_3_1_io_outs_right[38] ;
 wire \ces_3_1_io_outs_right[39] ;
 wire \ces_3_1_io_outs_right[3] ;
 wire \ces_3_1_io_outs_right[40] ;
 wire \ces_3_1_io_outs_right[41] ;
 wire \ces_3_1_io_outs_right[42] ;
 wire \ces_3_1_io_outs_right[43] ;
 wire \ces_3_1_io_outs_right[44] ;
 wire \ces_3_1_io_outs_right[45] ;
 wire \ces_3_1_io_outs_right[46] ;
 wire \ces_3_1_io_outs_right[47] ;
 wire \ces_3_1_io_outs_right[48] ;
 wire \ces_3_1_io_outs_right[49] ;
 wire \ces_3_1_io_outs_right[4] ;
 wire \ces_3_1_io_outs_right[50] ;
 wire \ces_3_1_io_outs_right[51] ;
 wire \ces_3_1_io_outs_right[52] ;
 wire \ces_3_1_io_outs_right[53] ;
 wire \ces_3_1_io_outs_right[54] ;
 wire \ces_3_1_io_outs_right[55] ;
 wire \ces_3_1_io_outs_right[56] ;
 wire \ces_3_1_io_outs_right[57] ;
 wire \ces_3_1_io_outs_right[58] ;
 wire \ces_3_1_io_outs_right[59] ;
 wire \ces_3_1_io_outs_right[5] ;
 wire \ces_3_1_io_outs_right[60] ;
 wire \ces_3_1_io_outs_right[61] ;
 wire \ces_3_1_io_outs_right[62] ;
 wire \ces_3_1_io_outs_right[63] ;
 wire \ces_3_1_io_outs_right[6] ;
 wire \ces_3_1_io_outs_right[7] ;
 wire \ces_3_1_io_outs_right[8] ;
 wire \ces_3_1_io_outs_right[9] ;
 wire \ces_3_1_io_outs_up[0] ;
 wire \ces_3_1_io_outs_up[10] ;
 wire \ces_3_1_io_outs_up[11] ;
 wire \ces_3_1_io_outs_up[12] ;
 wire \ces_3_1_io_outs_up[13] ;
 wire \ces_3_1_io_outs_up[14] ;
 wire \ces_3_1_io_outs_up[15] ;
 wire \ces_3_1_io_outs_up[16] ;
 wire \ces_3_1_io_outs_up[17] ;
 wire \ces_3_1_io_outs_up[18] ;
 wire \ces_3_1_io_outs_up[19] ;
 wire \ces_3_1_io_outs_up[1] ;
 wire \ces_3_1_io_outs_up[20] ;
 wire \ces_3_1_io_outs_up[21] ;
 wire \ces_3_1_io_outs_up[22] ;
 wire \ces_3_1_io_outs_up[23] ;
 wire \ces_3_1_io_outs_up[24] ;
 wire \ces_3_1_io_outs_up[25] ;
 wire \ces_3_1_io_outs_up[26] ;
 wire \ces_3_1_io_outs_up[27] ;
 wire \ces_3_1_io_outs_up[28] ;
 wire \ces_3_1_io_outs_up[29] ;
 wire \ces_3_1_io_outs_up[2] ;
 wire \ces_3_1_io_outs_up[30] ;
 wire \ces_3_1_io_outs_up[31] ;
 wire \ces_3_1_io_outs_up[32] ;
 wire \ces_3_1_io_outs_up[33] ;
 wire \ces_3_1_io_outs_up[34] ;
 wire \ces_3_1_io_outs_up[35] ;
 wire \ces_3_1_io_outs_up[36] ;
 wire \ces_3_1_io_outs_up[37] ;
 wire \ces_3_1_io_outs_up[38] ;
 wire \ces_3_1_io_outs_up[39] ;
 wire \ces_3_1_io_outs_up[3] ;
 wire \ces_3_1_io_outs_up[40] ;
 wire \ces_3_1_io_outs_up[41] ;
 wire \ces_3_1_io_outs_up[42] ;
 wire \ces_3_1_io_outs_up[43] ;
 wire \ces_3_1_io_outs_up[44] ;
 wire \ces_3_1_io_outs_up[45] ;
 wire \ces_3_1_io_outs_up[46] ;
 wire \ces_3_1_io_outs_up[47] ;
 wire \ces_3_1_io_outs_up[48] ;
 wire \ces_3_1_io_outs_up[49] ;
 wire \ces_3_1_io_outs_up[4] ;
 wire \ces_3_1_io_outs_up[50] ;
 wire \ces_3_1_io_outs_up[51] ;
 wire \ces_3_1_io_outs_up[52] ;
 wire \ces_3_1_io_outs_up[53] ;
 wire \ces_3_1_io_outs_up[54] ;
 wire \ces_3_1_io_outs_up[55] ;
 wire \ces_3_1_io_outs_up[56] ;
 wire \ces_3_1_io_outs_up[57] ;
 wire \ces_3_1_io_outs_up[58] ;
 wire \ces_3_1_io_outs_up[59] ;
 wire \ces_3_1_io_outs_up[5] ;
 wire \ces_3_1_io_outs_up[60] ;
 wire \ces_3_1_io_outs_up[61] ;
 wire \ces_3_1_io_outs_up[62] ;
 wire \ces_3_1_io_outs_up[63] ;
 wire \ces_3_1_io_outs_up[6] ;
 wire \ces_3_1_io_outs_up[7] ;
 wire \ces_3_1_io_outs_up[8] ;
 wire \ces_3_1_io_outs_up[9] ;
 wire \ces_3_2_io_ins_down[0] ;
 wire \ces_3_2_io_ins_down[10] ;
 wire \ces_3_2_io_ins_down[11] ;
 wire \ces_3_2_io_ins_down[12] ;
 wire \ces_3_2_io_ins_down[13] ;
 wire \ces_3_2_io_ins_down[14] ;
 wire \ces_3_2_io_ins_down[15] ;
 wire \ces_3_2_io_ins_down[16] ;
 wire \ces_3_2_io_ins_down[17] ;
 wire \ces_3_2_io_ins_down[18] ;
 wire \ces_3_2_io_ins_down[19] ;
 wire \ces_3_2_io_ins_down[1] ;
 wire \ces_3_2_io_ins_down[20] ;
 wire \ces_3_2_io_ins_down[21] ;
 wire \ces_3_2_io_ins_down[22] ;
 wire \ces_3_2_io_ins_down[23] ;
 wire \ces_3_2_io_ins_down[24] ;
 wire \ces_3_2_io_ins_down[25] ;
 wire \ces_3_2_io_ins_down[26] ;
 wire \ces_3_2_io_ins_down[27] ;
 wire \ces_3_2_io_ins_down[28] ;
 wire \ces_3_2_io_ins_down[29] ;
 wire \ces_3_2_io_ins_down[2] ;
 wire \ces_3_2_io_ins_down[30] ;
 wire \ces_3_2_io_ins_down[31] ;
 wire \ces_3_2_io_ins_down[32] ;
 wire \ces_3_2_io_ins_down[33] ;
 wire \ces_3_2_io_ins_down[34] ;
 wire \ces_3_2_io_ins_down[35] ;
 wire \ces_3_2_io_ins_down[36] ;
 wire \ces_3_2_io_ins_down[37] ;
 wire \ces_3_2_io_ins_down[38] ;
 wire \ces_3_2_io_ins_down[39] ;
 wire \ces_3_2_io_ins_down[3] ;
 wire \ces_3_2_io_ins_down[40] ;
 wire \ces_3_2_io_ins_down[41] ;
 wire \ces_3_2_io_ins_down[42] ;
 wire \ces_3_2_io_ins_down[43] ;
 wire \ces_3_2_io_ins_down[44] ;
 wire \ces_3_2_io_ins_down[45] ;
 wire \ces_3_2_io_ins_down[46] ;
 wire \ces_3_2_io_ins_down[47] ;
 wire \ces_3_2_io_ins_down[48] ;
 wire \ces_3_2_io_ins_down[49] ;
 wire \ces_3_2_io_ins_down[4] ;
 wire \ces_3_2_io_ins_down[50] ;
 wire \ces_3_2_io_ins_down[51] ;
 wire \ces_3_2_io_ins_down[52] ;
 wire \ces_3_2_io_ins_down[53] ;
 wire \ces_3_2_io_ins_down[54] ;
 wire \ces_3_2_io_ins_down[55] ;
 wire \ces_3_2_io_ins_down[56] ;
 wire \ces_3_2_io_ins_down[57] ;
 wire \ces_3_2_io_ins_down[58] ;
 wire \ces_3_2_io_ins_down[59] ;
 wire \ces_3_2_io_ins_down[5] ;
 wire \ces_3_2_io_ins_down[60] ;
 wire \ces_3_2_io_ins_down[61] ;
 wire \ces_3_2_io_ins_down[62] ;
 wire \ces_3_2_io_ins_down[63] ;
 wire \ces_3_2_io_ins_down[6] ;
 wire \ces_3_2_io_ins_down[7] ;
 wire \ces_3_2_io_ins_down[8] ;
 wire \ces_3_2_io_ins_down[9] ;
 wire \ces_3_2_io_ins_left[0] ;
 wire \ces_3_2_io_ins_left[10] ;
 wire \ces_3_2_io_ins_left[11] ;
 wire \ces_3_2_io_ins_left[12] ;
 wire \ces_3_2_io_ins_left[13] ;
 wire \ces_3_2_io_ins_left[14] ;
 wire \ces_3_2_io_ins_left[15] ;
 wire \ces_3_2_io_ins_left[16] ;
 wire \ces_3_2_io_ins_left[17] ;
 wire \ces_3_2_io_ins_left[18] ;
 wire \ces_3_2_io_ins_left[19] ;
 wire \ces_3_2_io_ins_left[1] ;
 wire \ces_3_2_io_ins_left[20] ;
 wire \ces_3_2_io_ins_left[21] ;
 wire \ces_3_2_io_ins_left[22] ;
 wire \ces_3_2_io_ins_left[23] ;
 wire \ces_3_2_io_ins_left[24] ;
 wire \ces_3_2_io_ins_left[25] ;
 wire \ces_3_2_io_ins_left[26] ;
 wire \ces_3_2_io_ins_left[27] ;
 wire \ces_3_2_io_ins_left[28] ;
 wire \ces_3_2_io_ins_left[29] ;
 wire \ces_3_2_io_ins_left[2] ;
 wire \ces_3_2_io_ins_left[30] ;
 wire \ces_3_2_io_ins_left[31] ;
 wire \ces_3_2_io_ins_left[32] ;
 wire \ces_3_2_io_ins_left[33] ;
 wire \ces_3_2_io_ins_left[34] ;
 wire \ces_3_2_io_ins_left[35] ;
 wire \ces_3_2_io_ins_left[36] ;
 wire \ces_3_2_io_ins_left[37] ;
 wire \ces_3_2_io_ins_left[38] ;
 wire \ces_3_2_io_ins_left[39] ;
 wire \ces_3_2_io_ins_left[3] ;
 wire \ces_3_2_io_ins_left[40] ;
 wire \ces_3_2_io_ins_left[41] ;
 wire \ces_3_2_io_ins_left[42] ;
 wire \ces_3_2_io_ins_left[43] ;
 wire \ces_3_2_io_ins_left[44] ;
 wire \ces_3_2_io_ins_left[45] ;
 wire \ces_3_2_io_ins_left[46] ;
 wire \ces_3_2_io_ins_left[47] ;
 wire \ces_3_2_io_ins_left[48] ;
 wire \ces_3_2_io_ins_left[49] ;
 wire \ces_3_2_io_ins_left[4] ;
 wire \ces_3_2_io_ins_left[50] ;
 wire \ces_3_2_io_ins_left[51] ;
 wire \ces_3_2_io_ins_left[52] ;
 wire \ces_3_2_io_ins_left[53] ;
 wire \ces_3_2_io_ins_left[54] ;
 wire \ces_3_2_io_ins_left[55] ;
 wire \ces_3_2_io_ins_left[56] ;
 wire \ces_3_2_io_ins_left[57] ;
 wire \ces_3_2_io_ins_left[58] ;
 wire \ces_3_2_io_ins_left[59] ;
 wire \ces_3_2_io_ins_left[5] ;
 wire \ces_3_2_io_ins_left[60] ;
 wire \ces_3_2_io_ins_left[61] ;
 wire \ces_3_2_io_ins_left[62] ;
 wire \ces_3_2_io_ins_left[63] ;
 wire \ces_3_2_io_ins_left[6] ;
 wire \ces_3_2_io_ins_left[7] ;
 wire \ces_3_2_io_ins_left[8] ;
 wire \ces_3_2_io_ins_left[9] ;
 wire ces_3_2_io_lsbOuts_0;
 wire ces_3_2_io_lsbOuts_1;
 wire ces_3_2_io_lsbOuts_2;
 wire ces_3_2_io_lsbOuts_3;
 wire ces_3_2_io_lsbOuts_4;
 wire ces_3_2_io_lsbOuts_5;
 wire ces_3_2_io_lsbOuts_6;
 wire ces_3_2_io_lsbOuts_7;
 wire \ces_3_2_io_outs_right[0] ;
 wire \ces_3_2_io_outs_right[10] ;
 wire \ces_3_2_io_outs_right[11] ;
 wire \ces_3_2_io_outs_right[12] ;
 wire \ces_3_2_io_outs_right[13] ;
 wire \ces_3_2_io_outs_right[14] ;
 wire \ces_3_2_io_outs_right[15] ;
 wire \ces_3_2_io_outs_right[16] ;
 wire \ces_3_2_io_outs_right[17] ;
 wire \ces_3_2_io_outs_right[18] ;
 wire \ces_3_2_io_outs_right[19] ;
 wire \ces_3_2_io_outs_right[1] ;
 wire \ces_3_2_io_outs_right[20] ;
 wire \ces_3_2_io_outs_right[21] ;
 wire \ces_3_2_io_outs_right[22] ;
 wire \ces_3_2_io_outs_right[23] ;
 wire \ces_3_2_io_outs_right[24] ;
 wire \ces_3_2_io_outs_right[25] ;
 wire \ces_3_2_io_outs_right[26] ;
 wire \ces_3_2_io_outs_right[27] ;
 wire \ces_3_2_io_outs_right[28] ;
 wire \ces_3_2_io_outs_right[29] ;
 wire \ces_3_2_io_outs_right[2] ;
 wire \ces_3_2_io_outs_right[30] ;
 wire \ces_3_2_io_outs_right[31] ;
 wire \ces_3_2_io_outs_right[32] ;
 wire \ces_3_2_io_outs_right[33] ;
 wire \ces_3_2_io_outs_right[34] ;
 wire \ces_3_2_io_outs_right[35] ;
 wire \ces_3_2_io_outs_right[36] ;
 wire \ces_3_2_io_outs_right[37] ;
 wire \ces_3_2_io_outs_right[38] ;
 wire \ces_3_2_io_outs_right[39] ;
 wire \ces_3_2_io_outs_right[3] ;
 wire \ces_3_2_io_outs_right[40] ;
 wire \ces_3_2_io_outs_right[41] ;
 wire \ces_3_2_io_outs_right[42] ;
 wire \ces_3_2_io_outs_right[43] ;
 wire \ces_3_2_io_outs_right[44] ;
 wire \ces_3_2_io_outs_right[45] ;
 wire \ces_3_2_io_outs_right[46] ;
 wire \ces_3_2_io_outs_right[47] ;
 wire \ces_3_2_io_outs_right[48] ;
 wire \ces_3_2_io_outs_right[49] ;
 wire \ces_3_2_io_outs_right[4] ;
 wire \ces_3_2_io_outs_right[50] ;
 wire \ces_3_2_io_outs_right[51] ;
 wire \ces_3_2_io_outs_right[52] ;
 wire \ces_3_2_io_outs_right[53] ;
 wire \ces_3_2_io_outs_right[54] ;
 wire \ces_3_2_io_outs_right[55] ;
 wire \ces_3_2_io_outs_right[56] ;
 wire \ces_3_2_io_outs_right[57] ;
 wire \ces_3_2_io_outs_right[58] ;
 wire \ces_3_2_io_outs_right[59] ;
 wire \ces_3_2_io_outs_right[5] ;
 wire \ces_3_2_io_outs_right[60] ;
 wire \ces_3_2_io_outs_right[61] ;
 wire \ces_3_2_io_outs_right[62] ;
 wire \ces_3_2_io_outs_right[63] ;
 wire \ces_3_2_io_outs_right[6] ;
 wire \ces_3_2_io_outs_right[7] ;
 wire \ces_3_2_io_outs_right[8] ;
 wire \ces_3_2_io_outs_right[9] ;
 wire \ces_3_2_io_outs_up[0] ;
 wire \ces_3_2_io_outs_up[10] ;
 wire \ces_3_2_io_outs_up[11] ;
 wire \ces_3_2_io_outs_up[12] ;
 wire \ces_3_2_io_outs_up[13] ;
 wire \ces_3_2_io_outs_up[14] ;
 wire \ces_3_2_io_outs_up[15] ;
 wire \ces_3_2_io_outs_up[16] ;
 wire \ces_3_2_io_outs_up[17] ;
 wire \ces_3_2_io_outs_up[18] ;
 wire \ces_3_2_io_outs_up[19] ;
 wire \ces_3_2_io_outs_up[1] ;
 wire \ces_3_2_io_outs_up[20] ;
 wire \ces_3_2_io_outs_up[21] ;
 wire \ces_3_2_io_outs_up[22] ;
 wire \ces_3_2_io_outs_up[23] ;
 wire \ces_3_2_io_outs_up[24] ;
 wire \ces_3_2_io_outs_up[25] ;
 wire \ces_3_2_io_outs_up[26] ;
 wire \ces_3_2_io_outs_up[27] ;
 wire \ces_3_2_io_outs_up[28] ;
 wire \ces_3_2_io_outs_up[29] ;
 wire \ces_3_2_io_outs_up[2] ;
 wire \ces_3_2_io_outs_up[30] ;
 wire \ces_3_2_io_outs_up[31] ;
 wire \ces_3_2_io_outs_up[32] ;
 wire \ces_3_2_io_outs_up[33] ;
 wire \ces_3_2_io_outs_up[34] ;
 wire \ces_3_2_io_outs_up[35] ;
 wire \ces_3_2_io_outs_up[36] ;
 wire \ces_3_2_io_outs_up[37] ;
 wire \ces_3_2_io_outs_up[38] ;
 wire \ces_3_2_io_outs_up[39] ;
 wire \ces_3_2_io_outs_up[3] ;
 wire \ces_3_2_io_outs_up[40] ;
 wire \ces_3_2_io_outs_up[41] ;
 wire \ces_3_2_io_outs_up[42] ;
 wire \ces_3_2_io_outs_up[43] ;
 wire \ces_3_2_io_outs_up[44] ;
 wire \ces_3_2_io_outs_up[45] ;
 wire \ces_3_2_io_outs_up[46] ;
 wire \ces_3_2_io_outs_up[47] ;
 wire \ces_3_2_io_outs_up[48] ;
 wire \ces_3_2_io_outs_up[49] ;
 wire \ces_3_2_io_outs_up[4] ;
 wire \ces_3_2_io_outs_up[50] ;
 wire \ces_3_2_io_outs_up[51] ;
 wire \ces_3_2_io_outs_up[52] ;
 wire \ces_3_2_io_outs_up[53] ;
 wire \ces_3_2_io_outs_up[54] ;
 wire \ces_3_2_io_outs_up[55] ;
 wire \ces_3_2_io_outs_up[56] ;
 wire \ces_3_2_io_outs_up[57] ;
 wire \ces_3_2_io_outs_up[58] ;
 wire \ces_3_2_io_outs_up[59] ;
 wire \ces_3_2_io_outs_up[5] ;
 wire \ces_3_2_io_outs_up[60] ;
 wire \ces_3_2_io_outs_up[61] ;
 wire \ces_3_2_io_outs_up[62] ;
 wire \ces_3_2_io_outs_up[63] ;
 wire \ces_3_2_io_outs_up[6] ;
 wire \ces_3_2_io_outs_up[7] ;
 wire \ces_3_2_io_outs_up[8] ;
 wire \ces_3_2_io_outs_up[9] ;
 wire \ces_3_3_io_ins_down[0] ;
 wire \ces_3_3_io_ins_down[10] ;
 wire \ces_3_3_io_ins_down[11] ;
 wire \ces_3_3_io_ins_down[12] ;
 wire \ces_3_3_io_ins_down[13] ;
 wire \ces_3_3_io_ins_down[14] ;
 wire \ces_3_3_io_ins_down[15] ;
 wire \ces_3_3_io_ins_down[16] ;
 wire \ces_3_3_io_ins_down[17] ;
 wire \ces_3_3_io_ins_down[18] ;
 wire \ces_3_3_io_ins_down[19] ;
 wire \ces_3_3_io_ins_down[1] ;
 wire \ces_3_3_io_ins_down[20] ;
 wire \ces_3_3_io_ins_down[21] ;
 wire \ces_3_3_io_ins_down[22] ;
 wire \ces_3_3_io_ins_down[23] ;
 wire \ces_3_3_io_ins_down[24] ;
 wire \ces_3_3_io_ins_down[25] ;
 wire \ces_3_3_io_ins_down[26] ;
 wire \ces_3_3_io_ins_down[27] ;
 wire \ces_3_3_io_ins_down[28] ;
 wire \ces_3_3_io_ins_down[29] ;
 wire \ces_3_3_io_ins_down[2] ;
 wire \ces_3_3_io_ins_down[30] ;
 wire \ces_3_3_io_ins_down[31] ;
 wire \ces_3_3_io_ins_down[32] ;
 wire \ces_3_3_io_ins_down[33] ;
 wire \ces_3_3_io_ins_down[34] ;
 wire \ces_3_3_io_ins_down[35] ;
 wire \ces_3_3_io_ins_down[36] ;
 wire \ces_3_3_io_ins_down[37] ;
 wire \ces_3_3_io_ins_down[38] ;
 wire \ces_3_3_io_ins_down[39] ;
 wire \ces_3_3_io_ins_down[3] ;
 wire \ces_3_3_io_ins_down[40] ;
 wire \ces_3_3_io_ins_down[41] ;
 wire \ces_3_3_io_ins_down[42] ;
 wire \ces_3_3_io_ins_down[43] ;
 wire \ces_3_3_io_ins_down[44] ;
 wire \ces_3_3_io_ins_down[45] ;
 wire \ces_3_3_io_ins_down[46] ;
 wire \ces_3_3_io_ins_down[47] ;
 wire \ces_3_3_io_ins_down[48] ;
 wire \ces_3_3_io_ins_down[49] ;
 wire \ces_3_3_io_ins_down[4] ;
 wire \ces_3_3_io_ins_down[50] ;
 wire \ces_3_3_io_ins_down[51] ;
 wire \ces_3_3_io_ins_down[52] ;
 wire \ces_3_3_io_ins_down[53] ;
 wire \ces_3_3_io_ins_down[54] ;
 wire \ces_3_3_io_ins_down[55] ;
 wire \ces_3_3_io_ins_down[56] ;
 wire \ces_3_3_io_ins_down[57] ;
 wire \ces_3_3_io_ins_down[58] ;
 wire \ces_3_3_io_ins_down[59] ;
 wire \ces_3_3_io_ins_down[5] ;
 wire \ces_3_3_io_ins_down[60] ;
 wire \ces_3_3_io_ins_down[61] ;
 wire \ces_3_3_io_ins_down[62] ;
 wire \ces_3_3_io_ins_down[63] ;
 wire \ces_3_3_io_ins_down[6] ;
 wire \ces_3_3_io_ins_down[7] ;
 wire \ces_3_3_io_ins_down[8] ;
 wire \ces_3_3_io_ins_down[9] ;
 wire \ces_3_3_io_ins_left[0] ;
 wire \ces_3_3_io_ins_left[10] ;
 wire \ces_3_3_io_ins_left[11] ;
 wire \ces_3_3_io_ins_left[12] ;
 wire \ces_3_3_io_ins_left[13] ;
 wire \ces_3_3_io_ins_left[14] ;
 wire \ces_3_3_io_ins_left[15] ;
 wire \ces_3_3_io_ins_left[16] ;
 wire \ces_3_3_io_ins_left[17] ;
 wire \ces_3_3_io_ins_left[18] ;
 wire \ces_3_3_io_ins_left[19] ;
 wire \ces_3_3_io_ins_left[1] ;
 wire \ces_3_3_io_ins_left[20] ;
 wire \ces_3_3_io_ins_left[21] ;
 wire \ces_3_3_io_ins_left[22] ;
 wire \ces_3_3_io_ins_left[23] ;
 wire \ces_3_3_io_ins_left[24] ;
 wire \ces_3_3_io_ins_left[25] ;
 wire \ces_3_3_io_ins_left[26] ;
 wire \ces_3_3_io_ins_left[27] ;
 wire \ces_3_3_io_ins_left[28] ;
 wire \ces_3_3_io_ins_left[29] ;
 wire \ces_3_3_io_ins_left[2] ;
 wire \ces_3_3_io_ins_left[30] ;
 wire \ces_3_3_io_ins_left[31] ;
 wire \ces_3_3_io_ins_left[32] ;
 wire \ces_3_3_io_ins_left[33] ;
 wire \ces_3_3_io_ins_left[34] ;
 wire \ces_3_3_io_ins_left[35] ;
 wire \ces_3_3_io_ins_left[36] ;
 wire \ces_3_3_io_ins_left[37] ;
 wire \ces_3_3_io_ins_left[38] ;
 wire \ces_3_3_io_ins_left[39] ;
 wire \ces_3_3_io_ins_left[3] ;
 wire \ces_3_3_io_ins_left[40] ;
 wire \ces_3_3_io_ins_left[41] ;
 wire \ces_3_3_io_ins_left[42] ;
 wire \ces_3_3_io_ins_left[43] ;
 wire \ces_3_3_io_ins_left[44] ;
 wire \ces_3_3_io_ins_left[45] ;
 wire \ces_3_3_io_ins_left[46] ;
 wire \ces_3_3_io_ins_left[47] ;
 wire \ces_3_3_io_ins_left[48] ;
 wire \ces_3_3_io_ins_left[49] ;
 wire \ces_3_3_io_ins_left[4] ;
 wire \ces_3_3_io_ins_left[50] ;
 wire \ces_3_3_io_ins_left[51] ;
 wire \ces_3_3_io_ins_left[52] ;
 wire \ces_3_3_io_ins_left[53] ;
 wire \ces_3_3_io_ins_left[54] ;
 wire \ces_3_3_io_ins_left[55] ;
 wire \ces_3_3_io_ins_left[56] ;
 wire \ces_3_3_io_ins_left[57] ;
 wire \ces_3_3_io_ins_left[58] ;
 wire \ces_3_3_io_ins_left[59] ;
 wire \ces_3_3_io_ins_left[5] ;
 wire \ces_3_3_io_ins_left[60] ;
 wire \ces_3_3_io_ins_left[61] ;
 wire \ces_3_3_io_ins_left[62] ;
 wire \ces_3_3_io_ins_left[63] ;
 wire \ces_3_3_io_ins_left[6] ;
 wire \ces_3_3_io_ins_left[7] ;
 wire \ces_3_3_io_ins_left[8] ;
 wire \ces_3_3_io_ins_left[9] ;
 wire ces_3_3_io_lsbOuts_0;
 wire ces_3_3_io_lsbOuts_1;
 wire ces_3_3_io_lsbOuts_2;
 wire ces_3_3_io_lsbOuts_3;
 wire ces_3_3_io_lsbOuts_4;
 wire ces_3_3_io_lsbOuts_5;
 wire ces_3_3_io_lsbOuts_6;
 wire ces_3_3_io_lsbOuts_7;
 wire \ces_3_3_io_outs_right[0] ;
 wire \ces_3_3_io_outs_right[10] ;
 wire \ces_3_3_io_outs_right[11] ;
 wire \ces_3_3_io_outs_right[12] ;
 wire \ces_3_3_io_outs_right[13] ;
 wire \ces_3_3_io_outs_right[14] ;
 wire \ces_3_3_io_outs_right[15] ;
 wire \ces_3_3_io_outs_right[16] ;
 wire \ces_3_3_io_outs_right[17] ;
 wire \ces_3_3_io_outs_right[18] ;
 wire \ces_3_3_io_outs_right[19] ;
 wire \ces_3_3_io_outs_right[1] ;
 wire \ces_3_3_io_outs_right[20] ;
 wire \ces_3_3_io_outs_right[21] ;
 wire \ces_3_3_io_outs_right[22] ;
 wire \ces_3_3_io_outs_right[23] ;
 wire \ces_3_3_io_outs_right[24] ;
 wire \ces_3_3_io_outs_right[25] ;
 wire \ces_3_3_io_outs_right[26] ;
 wire \ces_3_3_io_outs_right[27] ;
 wire \ces_3_3_io_outs_right[28] ;
 wire \ces_3_3_io_outs_right[29] ;
 wire \ces_3_3_io_outs_right[2] ;
 wire \ces_3_3_io_outs_right[30] ;
 wire \ces_3_3_io_outs_right[31] ;
 wire \ces_3_3_io_outs_right[32] ;
 wire \ces_3_3_io_outs_right[33] ;
 wire \ces_3_3_io_outs_right[34] ;
 wire \ces_3_3_io_outs_right[35] ;
 wire \ces_3_3_io_outs_right[36] ;
 wire \ces_3_3_io_outs_right[37] ;
 wire \ces_3_3_io_outs_right[38] ;
 wire \ces_3_3_io_outs_right[39] ;
 wire \ces_3_3_io_outs_right[3] ;
 wire \ces_3_3_io_outs_right[40] ;
 wire \ces_3_3_io_outs_right[41] ;
 wire \ces_3_3_io_outs_right[42] ;
 wire \ces_3_3_io_outs_right[43] ;
 wire \ces_3_3_io_outs_right[44] ;
 wire \ces_3_3_io_outs_right[45] ;
 wire \ces_3_3_io_outs_right[46] ;
 wire \ces_3_3_io_outs_right[47] ;
 wire \ces_3_3_io_outs_right[48] ;
 wire \ces_3_3_io_outs_right[49] ;
 wire \ces_3_3_io_outs_right[4] ;
 wire \ces_3_3_io_outs_right[50] ;
 wire \ces_3_3_io_outs_right[51] ;
 wire \ces_3_3_io_outs_right[52] ;
 wire \ces_3_3_io_outs_right[53] ;
 wire \ces_3_3_io_outs_right[54] ;
 wire \ces_3_3_io_outs_right[55] ;
 wire \ces_3_3_io_outs_right[56] ;
 wire \ces_3_3_io_outs_right[57] ;
 wire \ces_3_3_io_outs_right[58] ;
 wire \ces_3_3_io_outs_right[59] ;
 wire \ces_3_3_io_outs_right[5] ;
 wire \ces_3_3_io_outs_right[60] ;
 wire \ces_3_3_io_outs_right[61] ;
 wire \ces_3_3_io_outs_right[62] ;
 wire \ces_3_3_io_outs_right[63] ;
 wire \ces_3_3_io_outs_right[6] ;
 wire \ces_3_3_io_outs_right[7] ;
 wire \ces_3_3_io_outs_right[8] ;
 wire \ces_3_3_io_outs_right[9] ;
 wire \ces_3_3_io_outs_up[0] ;
 wire \ces_3_3_io_outs_up[10] ;
 wire \ces_3_3_io_outs_up[11] ;
 wire \ces_3_3_io_outs_up[12] ;
 wire \ces_3_3_io_outs_up[13] ;
 wire \ces_3_3_io_outs_up[14] ;
 wire \ces_3_3_io_outs_up[15] ;
 wire \ces_3_3_io_outs_up[16] ;
 wire \ces_3_3_io_outs_up[17] ;
 wire \ces_3_3_io_outs_up[18] ;
 wire \ces_3_3_io_outs_up[19] ;
 wire \ces_3_3_io_outs_up[1] ;
 wire \ces_3_3_io_outs_up[20] ;
 wire \ces_3_3_io_outs_up[21] ;
 wire \ces_3_3_io_outs_up[22] ;
 wire \ces_3_3_io_outs_up[23] ;
 wire \ces_3_3_io_outs_up[24] ;
 wire \ces_3_3_io_outs_up[25] ;
 wire \ces_3_3_io_outs_up[26] ;
 wire \ces_3_3_io_outs_up[27] ;
 wire \ces_3_3_io_outs_up[28] ;
 wire \ces_3_3_io_outs_up[29] ;
 wire \ces_3_3_io_outs_up[2] ;
 wire \ces_3_3_io_outs_up[30] ;
 wire \ces_3_3_io_outs_up[31] ;
 wire \ces_3_3_io_outs_up[32] ;
 wire \ces_3_3_io_outs_up[33] ;
 wire \ces_3_3_io_outs_up[34] ;
 wire \ces_3_3_io_outs_up[35] ;
 wire \ces_3_3_io_outs_up[36] ;
 wire \ces_3_3_io_outs_up[37] ;
 wire \ces_3_3_io_outs_up[38] ;
 wire \ces_3_3_io_outs_up[39] ;
 wire \ces_3_3_io_outs_up[3] ;
 wire \ces_3_3_io_outs_up[40] ;
 wire \ces_3_3_io_outs_up[41] ;
 wire \ces_3_3_io_outs_up[42] ;
 wire \ces_3_3_io_outs_up[43] ;
 wire \ces_3_3_io_outs_up[44] ;
 wire \ces_3_3_io_outs_up[45] ;
 wire \ces_3_3_io_outs_up[46] ;
 wire \ces_3_3_io_outs_up[47] ;
 wire \ces_3_3_io_outs_up[48] ;
 wire \ces_3_3_io_outs_up[49] ;
 wire \ces_3_3_io_outs_up[4] ;
 wire \ces_3_3_io_outs_up[50] ;
 wire \ces_3_3_io_outs_up[51] ;
 wire \ces_3_3_io_outs_up[52] ;
 wire \ces_3_3_io_outs_up[53] ;
 wire \ces_3_3_io_outs_up[54] ;
 wire \ces_3_3_io_outs_up[55] ;
 wire \ces_3_3_io_outs_up[56] ;
 wire \ces_3_3_io_outs_up[57] ;
 wire \ces_3_3_io_outs_up[58] ;
 wire \ces_3_3_io_outs_up[59] ;
 wire \ces_3_3_io_outs_up[5] ;
 wire \ces_3_3_io_outs_up[60] ;
 wire \ces_3_3_io_outs_up[61] ;
 wire \ces_3_3_io_outs_up[62] ;
 wire \ces_3_3_io_outs_up[63] ;
 wire \ces_3_3_io_outs_up[6] ;
 wire \ces_3_3_io_outs_up[7] ;
 wire \ces_3_3_io_outs_up[8] ;
 wire \ces_3_3_io_outs_up[9] ;
 wire \ces_3_4_io_ins_down[0] ;
 wire \ces_3_4_io_ins_down[10] ;
 wire \ces_3_4_io_ins_down[11] ;
 wire \ces_3_4_io_ins_down[12] ;
 wire \ces_3_4_io_ins_down[13] ;
 wire \ces_3_4_io_ins_down[14] ;
 wire \ces_3_4_io_ins_down[15] ;
 wire \ces_3_4_io_ins_down[16] ;
 wire \ces_3_4_io_ins_down[17] ;
 wire \ces_3_4_io_ins_down[18] ;
 wire \ces_3_4_io_ins_down[19] ;
 wire \ces_3_4_io_ins_down[1] ;
 wire \ces_3_4_io_ins_down[20] ;
 wire \ces_3_4_io_ins_down[21] ;
 wire \ces_3_4_io_ins_down[22] ;
 wire \ces_3_4_io_ins_down[23] ;
 wire \ces_3_4_io_ins_down[24] ;
 wire \ces_3_4_io_ins_down[25] ;
 wire \ces_3_4_io_ins_down[26] ;
 wire \ces_3_4_io_ins_down[27] ;
 wire \ces_3_4_io_ins_down[28] ;
 wire \ces_3_4_io_ins_down[29] ;
 wire \ces_3_4_io_ins_down[2] ;
 wire \ces_3_4_io_ins_down[30] ;
 wire \ces_3_4_io_ins_down[31] ;
 wire \ces_3_4_io_ins_down[32] ;
 wire \ces_3_4_io_ins_down[33] ;
 wire \ces_3_4_io_ins_down[34] ;
 wire \ces_3_4_io_ins_down[35] ;
 wire \ces_3_4_io_ins_down[36] ;
 wire \ces_3_4_io_ins_down[37] ;
 wire \ces_3_4_io_ins_down[38] ;
 wire \ces_3_4_io_ins_down[39] ;
 wire \ces_3_4_io_ins_down[3] ;
 wire \ces_3_4_io_ins_down[40] ;
 wire \ces_3_4_io_ins_down[41] ;
 wire \ces_3_4_io_ins_down[42] ;
 wire \ces_3_4_io_ins_down[43] ;
 wire \ces_3_4_io_ins_down[44] ;
 wire \ces_3_4_io_ins_down[45] ;
 wire \ces_3_4_io_ins_down[46] ;
 wire \ces_3_4_io_ins_down[47] ;
 wire \ces_3_4_io_ins_down[48] ;
 wire \ces_3_4_io_ins_down[49] ;
 wire \ces_3_4_io_ins_down[4] ;
 wire \ces_3_4_io_ins_down[50] ;
 wire \ces_3_4_io_ins_down[51] ;
 wire \ces_3_4_io_ins_down[52] ;
 wire \ces_3_4_io_ins_down[53] ;
 wire \ces_3_4_io_ins_down[54] ;
 wire \ces_3_4_io_ins_down[55] ;
 wire \ces_3_4_io_ins_down[56] ;
 wire \ces_3_4_io_ins_down[57] ;
 wire \ces_3_4_io_ins_down[58] ;
 wire \ces_3_4_io_ins_down[59] ;
 wire \ces_3_4_io_ins_down[5] ;
 wire \ces_3_4_io_ins_down[60] ;
 wire \ces_3_4_io_ins_down[61] ;
 wire \ces_3_4_io_ins_down[62] ;
 wire \ces_3_4_io_ins_down[63] ;
 wire \ces_3_4_io_ins_down[6] ;
 wire \ces_3_4_io_ins_down[7] ;
 wire \ces_3_4_io_ins_down[8] ;
 wire \ces_3_4_io_ins_down[9] ;
 wire \ces_3_4_io_ins_left[0] ;
 wire \ces_3_4_io_ins_left[10] ;
 wire \ces_3_4_io_ins_left[11] ;
 wire \ces_3_4_io_ins_left[12] ;
 wire \ces_3_4_io_ins_left[13] ;
 wire \ces_3_4_io_ins_left[14] ;
 wire \ces_3_4_io_ins_left[15] ;
 wire \ces_3_4_io_ins_left[16] ;
 wire \ces_3_4_io_ins_left[17] ;
 wire \ces_3_4_io_ins_left[18] ;
 wire \ces_3_4_io_ins_left[19] ;
 wire \ces_3_4_io_ins_left[1] ;
 wire \ces_3_4_io_ins_left[20] ;
 wire \ces_3_4_io_ins_left[21] ;
 wire \ces_3_4_io_ins_left[22] ;
 wire \ces_3_4_io_ins_left[23] ;
 wire \ces_3_4_io_ins_left[24] ;
 wire \ces_3_4_io_ins_left[25] ;
 wire \ces_3_4_io_ins_left[26] ;
 wire \ces_3_4_io_ins_left[27] ;
 wire \ces_3_4_io_ins_left[28] ;
 wire \ces_3_4_io_ins_left[29] ;
 wire \ces_3_4_io_ins_left[2] ;
 wire \ces_3_4_io_ins_left[30] ;
 wire \ces_3_4_io_ins_left[31] ;
 wire \ces_3_4_io_ins_left[32] ;
 wire \ces_3_4_io_ins_left[33] ;
 wire \ces_3_4_io_ins_left[34] ;
 wire \ces_3_4_io_ins_left[35] ;
 wire \ces_3_4_io_ins_left[36] ;
 wire \ces_3_4_io_ins_left[37] ;
 wire \ces_3_4_io_ins_left[38] ;
 wire \ces_3_4_io_ins_left[39] ;
 wire \ces_3_4_io_ins_left[3] ;
 wire \ces_3_4_io_ins_left[40] ;
 wire \ces_3_4_io_ins_left[41] ;
 wire \ces_3_4_io_ins_left[42] ;
 wire \ces_3_4_io_ins_left[43] ;
 wire \ces_3_4_io_ins_left[44] ;
 wire \ces_3_4_io_ins_left[45] ;
 wire \ces_3_4_io_ins_left[46] ;
 wire \ces_3_4_io_ins_left[47] ;
 wire \ces_3_4_io_ins_left[48] ;
 wire \ces_3_4_io_ins_left[49] ;
 wire \ces_3_4_io_ins_left[4] ;
 wire \ces_3_4_io_ins_left[50] ;
 wire \ces_3_4_io_ins_left[51] ;
 wire \ces_3_4_io_ins_left[52] ;
 wire \ces_3_4_io_ins_left[53] ;
 wire \ces_3_4_io_ins_left[54] ;
 wire \ces_3_4_io_ins_left[55] ;
 wire \ces_3_4_io_ins_left[56] ;
 wire \ces_3_4_io_ins_left[57] ;
 wire \ces_3_4_io_ins_left[58] ;
 wire \ces_3_4_io_ins_left[59] ;
 wire \ces_3_4_io_ins_left[5] ;
 wire \ces_3_4_io_ins_left[60] ;
 wire \ces_3_4_io_ins_left[61] ;
 wire \ces_3_4_io_ins_left[62] ;
 wire \ces_3_4_io_ins_left[63] ;
 wire \ces_3_4_io_ins_left[6] ;
 wire \ces_3_4_io_ins_left[7] ;
 wire \ces_3_4_io_ins_left[8] ;
 wire \ces_3_4_io_ins_left[9] ;
 wire ces_3_4_io_lsbOuts_0;
 wire ces_3_4_io_lsbOuts_1;
 wire ces_3_4_io_lsbOuts_2;
 wire ces_3_4_io_lsbOuts_3;
 wire ces_3_4_io_lsbOuts_4;
 wire ces_3_4_io_lsbOuts_5;
 wire ces_3_4_io_lsbOuts_6;
 wire ces_3_4_io_lsbOuts_7;
 wire \ces_3_4_io_outs_right[0] ;
 wire \ces_3_4_io_outs_right[10] ;
 wire \ces_3_4_io_outs_right[11] ;
 wire \ces_3_4_io_outs_right[12] ;
 wire \ces_3_4_io_outs_right[13] ;
 wire \ces_3_4_io_outs_right[14] ;
 wire \ces_3_4_io_outs_right[15] ;
 wire \ces_3_4_io_outs_right[16] ;
 wire \ces_3_4_io_outs_right[17] ;
 wire \ces_3_4_io_outs_right[18] ;
 wire \ces_3_4_io_outs_right[19] ;
 wire \ces_3_4_io_outs_right[1] ;
 wire \ces_3_4_io_outs_right[20] ;
 wire \ces_3_4_io_outs_right[21] ;
 wire \ces_3_4_io_outs_right[22] ;
 wire \ces_3_4_io_outs_right[23] ;
 wire \ces_3_4_io_outs_right[24] ;
 wire \ces_3_4_io_outs_right[25] ;
 wire \ces_3_4_io_outs_right[26] ;
 wire \ces_3_4_io_outs_right[27] ;
 wire \ces_3_4_io_outs_right[28] ;
 wire \ces_3_4_io_outs_right[29] ;
 wire \ces_3_4_io_outs_right[2] ;
 wire \ces_3_4_io_outs_right[30] ;
 wire \ces_3_4_io_outs_right[31] ;
 wire \ces_3_4_io_outs_right[32] ;
 wire \ces_3_4_io_outs_right[33] ;
 wire \ces_3_4_io_outs_right[34] ;
 wire \ces_3_4_io_outs_right[35] ;
 wire \ces_3_4_io_outs_right[36] ;
 wire \ces_3_4_io_outs_right[37] ;
 wire \ces_3_4_io_outs_right[38] ;
 wire \ces_3_4_io_outs_right[39] ;
 wire \ces_3_4_io_outs_right[3] ;
 wire \ces_3_4_io_outs_right[40] ;
 wire \ces_3_4_io_outs_right[41] ;
 wire \ces_3_4_io_outs_right[42] ;
 wire \ces_3_4_io_outs_right[43] ;
 wire \ces_3_4_io_outs_right[44] ;
 wire \ces_3_4_io_outs_right[45] ;
 wire \ces_3_4_io_outs_right[46] ;
 wire \ces_3_4_io_outs_right[47] ;
 wire \ces_3_4_io_outs_right[48] ;
 wire \ces_3_4_io_outs_right[49] ;
 wire \ces_3_4_io_outs_right[4] ;
 wire \ces_3_4_io_outs_right[50] ;
 wire \ces_3_4_io_outs_right[51] ;
 wire \ces_3_4_io_outs_right[52] ;
 wire \ces_3_4_io_outs_right[53] ;
 wire \ces_3_4_io_outs_right[54] ;
 wire \ces_3_4_io_outs_right[55] ;
 wire \ces_3_4_io_outs_right[56] ;
 wire \ces_3_4_io_outs_right[57] ;
 wire \ces_3_4_io_outs_right[58] ;
 wire \ces_3_4_io_outs_right[59] ;
 wire \ces_3_4_io_outs_right[5] ;
 wire \ces_3_4_io_outs_right[60] ;
 wire \ces_3_4_io_outs_right[61] ;
 wire \ces_3_4_io_outs_right[62] ;
 wire \ces_3_4_io_outs_right[63] ;
 wire \ces_3_4_io_outs_right[6] ;
 wire \ces_3_4_io_outs_right[7] ;
 wire \ces_3_4_io_outs_right[8] ;
 wire \ces_3_4_io_outs_right[9] ;
 wire \ces_3_4_io_outs_up[0] ;
 wire \ces_3_4_io_outs_up[10] ;
 wire \ces_3_4_io_outs_up[11] ;
 wire \ces_3_4_io_outs_up[12] ;
 wire \ces_3_4_io_outs_up[13] ;
 wire \ces_3_4_io_outs_up[14] ;
 wire \ces_3_4_io_outs_up[15] ;
 wire \ces_3_4_io_outs_up[16] ;
 wire \ces_3_4_io_outs_up[17] ;
 wire \ces_3_4_io_outs_up[18] ;
 wire \ces_3_4_io_outs_up[19] ;
 wire \ces_3_4_io_outs_up[1] ;
 wire \ces_3_4_io_outs_up[20] ;
 wire \ces_3_4_io_outs_up[21] ;
 wire \ces_3_4_io_outs_up[22] ;
 wire \ces_3_4_io_outs_up[23] ;
 wire \ces_3_4_io_outs_up[24] ;
 wire \ces_3_4_io_outs_up[25] ;
 wire \ces_3_4_io_outs_up[26] ;
 wire \ces_3_4_io_outs_up[27] ;
 wire \ces_3_4_io_outs_up[28] ;
 wire \ces_3_4_io_outs_up[29] ;
 wire \ces_3_4_io_outs_up[2] ;
 wire \ces_3_4_io_outs_up[30] ;
 wire \ces_3_4_io_outs_up[31] ;
 wire \ces_3_4_io_outs_up[32] ;
 wire \ces_3_4_io_outs_up[33] ;
 wire \ces_3_4_io_outs_up[34] ;
 wire \ces_3_4_io_outs_up[35] ;
 wire \ces_3_4_io_outs_up[36] ;
 wire \ces_3_4_io_outs_up[37] ;
 wire \ces_3_4_io_outs_up[38] ;
 wire \ces_3_4_io_outs_up[39] ;
 wire \ces_3_4_io_outs_up[3] ;
 wire \ces_3_4_io_outs_up[40] ;
 wire \ces_3_4_io_outs_up[41] ;
 wire \ces_3_4_io_outs_up[42] ;
 wire \ces_3_4_io_outs_up[43] ;
 wire \ces_3_4_io_outs_up[44] ;
 wire \ces_3_4_io_outs_up[45] ;
 wire \ces_3_4_io_outs_up[46] ;
 wire \ces_3_4_io_outs_up[47] ;
 wire \ces_3_4_io_outs_up[48] ;
 wire \ces_3_4_io_outs_up[49] ;
 wire \ces_3_4_io_outs_up[4] ;
 wire \ces_3_4_io_outs_up[50] ;
 wire \ces_3_4_io_outs_up[51] ;
 wire \ces_3_4_io_outs_up[52] ;
 wire \ces_3_4_io_outs_up[53] ;
 wire \ces_3_4_io_outs_up[54] ;
 wire \ces_3_4_io_outs_up[55] ;
 wire \ces_3_4_io_outs_up[56] ;
 wire \ces_3_4_io_outs_up[57] ;
 wire \ces_3_4_io_outs_up[58] ;
 wire \ces_3_4_io_outs_up[59] ;
 wire \ces_3_4_io_outs_up[5] ;
 wire \ces_3_4_io_outs_up[60] ;
 wire \ces_3_4_io_outs_up[61] ;
 wire \ces_3_4_io_outs_up[62] ;
 wire \ces_3_4_io_outs_up[63] ;
 wire \ces_3_4_io_outs_up[6] ;
 wire \ces_3_4_io_outs_up[7] ;
 wire \ces_3_4_io_outs_up[8] ;
 wire \ces_3_4_io_outs_up[9] ;
 wire \ces_3_5_io_ins_down[0] ;
 wire \ces_3_5_io_ins_down[10] ;
 wire \ces_3_5_io_ins_down[11] ;
 wire \ces_3_5_io_ins_down[12] ;
 wire \ces_3_5_io_ins_down[13] ;
 wire \ces_3_5_io_ins_down[14] ;
 wire \ces_3_5_io_ins_down[15] ;
 wire \ces_3_5_io_ins_down[16] ;
 wire \ces_3_5_io_ins_down[17] ;
 wire \ces_3_5_io_ins_down[18] ;
 wire \ces_3_5_io_ins_down[19] ;
 wire \ces_3_5_io_ins_down[1] ;
 wire \ces_3_5_io_ins_down[20] ;
 wire \ces_3_5_io_ins_down[21] ;
 wire \ces_3_5_io_ins_down[22] ;
 wire \ces_3_5_io_ins_down[23] ;
 wire \ces_3_5_io_ins_down[24] ;
 wire \ces_3_5_io_ins_down[25] ;
 wire \ces_3_5_io_ins_down[26] ;
 wire \ces_3_5_io_ins_down[27] ;
 wire \ces_3_5_io_ins_down[28] ;
 wire \ces_3_5_io_ins_down[29] ;
 wire \ces_3_5_io_ins_down[2] ;
 wire \ces_3_5_io_ins_down[30] ;
 wire \ces_3_5_io_ins_down[31] ;
 wire \ces_3_5_io_ins_down[32] ;
 wire \ces_3_5_io_ins_down[33] ;
 wire \ces_3_5_io_ins_down[34] ;
 wire \ces_3_5_io_ins_down[35] ;
 wire \ces_3_5_io_ins_down[36] ;
 wire \ces_3_5_io_ins_down[37] ;
 wire \ces_3_5_io_ins_down[38] ;
 wire \ces_3_5_io_ins_down[39] ;
 wire \ces_3_5_io_ins_down[3] ;
 wire \ces_3_5_io_ins_down[40] ;
 wire \ces_3_5_io_ins_down[41] ;
 wire \ces_3_5_io_ins_down[42] ;
 wire \ces_3_5_io_ins_down[43] ;
 wire \ces_3_5_io_ins_down[44] ;
 wire \ces_3_5_io_ins_down[45] ;
 wire \ces_3_5_io_ins_down[46] ;
 wire \ces_3_5_io_ins_down[47] ;
 wire \ces_3_5_io_ins_down[48] ;
 wire \ces_3_5_io_ins_down[49] ;
 wire \ces_3_5_io_ins_down[4] ;
 wire \ces_3_5_io_ins_down[50] ;
 wire \ces_3_5_io_ins_down[51] ;
 wire \ces_3_5_io_ins_down[52] ;
 wire \ces_3_5_io_ins_down[53] ;
 wire \ces_3_5_io_ins_down[54] ;
 wire \ces_3_5_io_ins_down[55] ;
 wire \ces_3_5_io_ins_down[56] ;
 wire \ces_3_5_io_ins_down[57] ;
 wire \ces_3_5_io_ins_down[58] ;
 wire \ces_3_5_io_ins_down[59] ;
 wire \ces_3_5_io_ins_down[5] ;
 wire \ces_3_5_io_ins_down[60] ;
 wire \ces_3_5_io_ins_down[61] ;
 wire \ces_3_5_io_ins_down[62] ;
 wire \ces_3_5_io_ins_down[63] ;
 wire \ces_3_5_io_ins_down[6] ;
 wire \ces_3_5_io_ins_down[7] ;
 wire \ces_3_5_io_ins_down[8] ;
 wire \ces_3_5_io_ins_down[9] ;
 wire \ces_3_5_io_ins_left[0] ;
 wire \ces_3_5_io_ins_left[10] ;
 wire \ces_3_5_io_ins_left[11] ;
 wire \ces_3_5_io_ins_left[12] ;
 wire \ces_3_5_io_ins_left[13] ;
 wire \ces_3_5_io_ins_left[14] ;
 wire \ces_3_5_io_ins_left[15] ;
 wire \ces_3_5_io_ins_left[16] ;
 wire \ces_3_5_io_ins_left[17] ;
 wire \ces_3_5_io_ins_left[18] ;
 wire \ces_3_5_io_ins_left[19] ;
 wire \ces_3_5_io_ins_left[1] ;
 wire \ces_3_5_io_ins_left[20] ;
 wire \ces_3_5_io_ins_left[21] ;
 wire \ces_3_5_io_ins_left[22] ;
 wire \ces_3_5_io_ins_left[23] ;
 wire \ces_3_5_io_ins_left[24] ;
 wire \ces_3_5_io_ins_left[25] ;
 wire \ces_3_5_io_ins_left[26] ;
 wire \ces_3_5_io_ins_left[27] ;
 wire \ces_3_5_io_ins_left[28] ;
 wire \ces_3_5_io_ins_left[29] ;
 wire \ces_3_5_io_ins_left[2] ;
 wire \ces_3_5_io_ins_left[30] ;
 wire \ces_3_5_io_ins_left[31] ;
 wire \ces_3_5_io_ins_left[32] ;
 wire \ces_3_5_io_ins_left[33] ;
 wire \ces_3_5_io_ins_left[34] ;
 wire \ces_3_5_io_ins_left[35] ;
 wire \ces_3_5_io_ins_left[36] ;
 wire \ces_3_5_io_ins_left[37] ;
 wire \ces_3_5_io_ins_left[38] ;
 wire \ces_3_5_io_ins_left[39] ;
 wire \ces_3_5_io_ins_left[3] ;
 wire \ces_3_5_io_ins_left[40] ;
 wire \ces_3_5_io_ins_left[41] ;
 wire \ces_3_5_io_ins_left[42] ;
 wire \ces_3_5_io_ins_left[43] ;
 wire \ces_3_5_io_ins_left[44] ;
 wire \ces_3_5_io_ins_left[45] ;
 wire \ces_3_5_io_ins_left[46] ;
 wire \ces_3_5_io_ins_left[47] ;
 wire \ces_3_5_io_ins_left[48] ;
 wire \ces_3_5_io_ins_left[49] ;
 wire \ces_3_5_io_ins_left[4] ;
 wire \ces_3_5_io_ins_left[50] ;
 wire \ces_3_5_io_ins_left[51] ;
 wire \ces_3_5_io_ins_left[52] ;
 wire \ces_3_5_io_ins_left[53] ;
 wire \ces_3_5_io_ins_left[54] ;
 wire \ces_3_5_io_ins_left[55] ;
 wire \ces_3_5_io_ins_left[56] ;
 wire \ces_3_5_io_ins_left[57] ;
 wire \ces_3_5_io_ins_left[58] ;
 wire \ces_3_5_io_ins_left[59] ;
 wire \ces_3_5_io_ins_left[5] ;
 wire \ces_3_5_io_ins_left[60] ;
 wire \ces_3_5_io_ins_left[61] ;
 wire \ces_3_5_io_ins_left[62] ;
 wire \ces_3_5_io_ins_left[63] ;
 wire \ces_3_5_io_ins_left[6] ;
 wire \ces_3_5_io_ins_left[7] ;
 wire \ces_3_5_io_ins_left[8] ;
 wire \ces_3_5_io_ins_left[9] ;
 wire ces_3_5_io_lsbOuts_0;
 wire ces_3_5_io_lsbOuts_1;
 wire ces_3_5_io_lsbOuts_2;
 wire ces_3_5_io_lsbOuts_3;
 wire ces_3_5_io_lsbOuts_4;
 wire ces_3_5_io_lsbOuts_5;
 wire ces_3_5_io_lsbOuts_6;
 wire ces_3_5_io_lsbOuts_7;
 wire \ces_3_5_io_outs_right[0] ;
 wire \ces_3_5_io_outs_right[10] ;
 wire \ces_3_5_io_outs_right[11] ;
 wire \ces_3_5_io_outs_right[12] ;
 wire \ces_3_5_io_outs_right[13] ;
 wire \ces_3_5_io_outs_right[14] ;
 wire \ces_3_5_io_outs_right[15] ;
 wire \ces_3_5_io_outs_right[16] ;
 wire \ces_3_5_io_outs_right[17] ;
 wire \ces_3_5_io_outs_right[18] ;
 wire \ces_3_5_io_outs_right[19] ;
 wire \ces_3_5_io_outs_right[1] ;
 wire \ces_3_5_io_outs_right[20] ;
 wire \ces_3_5_io_outs_right[21] ;
 wire \ces_3_5_io_outs_right[22] ;
 wire \ces_3_5_io_outs_right[23] ;
 wire \ces_3_5_io_outs_right[24] ;
 wire \ces_3_5_io_outs_right[25] ;
 wire \ces_3_5_io_outs_right[26] ;
 wire \ces_3_5_io_outs_right[27] ;
 wire \ces_3_5_io_outs_right[28] ;
 wire \ces_3_5_io_outs_right[29] ;
 wire \ces_3_5_io_outs_right[2] ;
 wire \ces_3_5_io_outs_right[30] ;
 wire \ces_3_5_io_outs_right[31] ;
 wire \ces_3_5_io_outs_right[32] ;
 wire \ces_3_5_io_outs_right[33] ;
 wire \ces_3_5_io_outs_right[34] ;
 wire \ces_3_5_io_outs_right[35] ;
 wire \ces_3_5_io_outs_right[36] ;
 wire \ces_3_5_io_outs_right[37] ;
 wire \ces_3_5_io_outs_right[38] ;
 wire \ces_3_5_io_outs_right[39] ;
 wire \ces_3_5_io_outs_right[3] ;
 wire \ces_3_5_io_outs_right[40] ;
 wire \ces_3_5_io_outs_right[41] ;
 wire \ces_3_5_io_outs_right[42] ;
 wire \ces_3_5_io_outs_right[43] ;
 wire \ces_3_5_io_outs_right[44] ;
 wire \ces_3_5_io_outs_right[45] ;
 wire \ces_3_5_io_outs_right[46] ;
 wire \ces_3_5_io_outs_right[47] ;
 wire \ces_3_5_io_outs_right[48] ;
 wire \ces_3_5_io_outs_right[49] ;
 wire \ces_3_5_io_outs_right[4] ;
 wire \ces_3_5_io_outs_right[50] ;
 wire \ces_3_5_io_outs_right[51] ;
 wire \ces_3_5_io_outs_right[52] ;
 wire \ces_3_5_io_outs_right[53] ;
 wire \ces_3_5_io_outs_right[54] ;
 wire \ces_3_5_io_outs_right[55] ;
 wire \ces_3_5_io_outs_right[56] ;
 wire \ces_3_5_io_outs_right[57] ;
 wire \ces_3_5_io_outs_right[58] ;
 wire \ces_3_5_io_outs_right[59] ;
 wire \ces_3_5_io_outs_right[5] ;
 wire \ces_3_5_io_outs_right[60] ;
 wire \ces_3_5_io_outs_right[61] ;
 wire \ces_3_5_io_outs_right[62] ;
 wire \ces_3_5_io_outs_right[63] ;
 wire \ces_3_5_io_outs_right[6] ;
 wire \ces_3_5_io_outs_right[7] ;
 wire \ces_3_5_io_outs_right[8] ;
 wire \ces_3_5_io_outs_right[9] ;
 wire \ces_3_5_io_outs_up[0] ;
 wire \ces_3_5_io_outs_up[10] ;
 wire \ces_3_5_io_outs_up[11] ;
 wire \ces_3_5_io_outs_up[12] ;
 wire \ces_3_5_io_outs_up[13] ;
 wire \ces_3_5_io_outs_up[14] ;
 wire \ces_3_5_io_outs_up[15] ;
 wire \ces_3_5_io_outs_up[16] ;
 wire \ces_3_5_io_outs_up[17] ;
 wire \ces_3_5_io_outs_up[18] ;
 wire \ces_3_5_io_outs_up[19] ;
 wire \ces_3_5_io_outs_up[1] ;
 wire \ces_3_5_io_outs_up[20] ;
 wire \ces_3_5_io_outs_up[21] ;
 wire \ces_3_5_io_outs_up[22] ;
 wire \ces_3_5_io_outs_up[23] ;
 wire \ces_3_5_io_outs_up[24] ;
 wire \ces_3_5_io_outs_up[25] ;
 wire \ces_3_5_io_outs_up[26] ;
 wire \ces_3_5_io_outs_up[27] ;
 wire \ces_3_5_io_outs_up[28] ;
 wire \ces_3_5_io_outs_up[29] ;
 wire \ces_3_5_io_outs_up[2] ;
 wire \ces_3_5_io_outs_up[30] ;
 wire \ces_3_5_io_outs_up[31] ;
 wire \ces_3_5_io_outs_up[32] ;
 wire \ces_3_5_io_outs_up[33] ;
 wire \ces_3_5_io_outs_up[34] ;
 wire \ces_3_5_io_outs_up[35] ;
 wire \ces_3_5_io_outs_up[36] ;
 wire \ces_3_5_io_outs_up[37] ;
 wire \ces_3_5_io_outs_up[38] ;
 wire \ces_3_5_io_outs_up[39] ;
 wire \ces_3_5_io_outs_up[3] ;
 wire \ces_3_5_io_outs_up[40] ;
 wire \ces_3_5_io_outs_up[41] ;
 wire \ces_3_5_io_outs_up[42] ;
 wire \ces_3_5_io_outs_up[43] ;
 wire \ces_3_5_io_outs_up[44] ;
 wire \ces_3_5_io_outs_up[45] ;
 wire \ces_3_5_io_outs_up[46] ;
 wire \ces_3_5_io_outs_up[47] ;
 wire \ces_3_5_io_outs_up[48] ;
 wire \ces_3_5_io_outs_up[49] ;
 wire \ces_3_5_io_outs_up[4] ;
 wire \ces_3_5_io_outs_up[50] ;
 wire \ces_3_5_io_outs_up[51] ;
 wire \ces_3_5_io_outs_up[52] ;
 wire \ces_3_5_io_outs_up[53] ;
 wire \ces_3_5_io_outs_up[54] ;
 wire \ces_3_5_io_outs_up[55] ;
 wire \ces_3_5_io_outs_up[56] ;
 wire \ces_3_5_io_outs_up[57] ;
 wire \ces_3_5_io_outs_up[58] ;
 wire \ces_3_5_io_outs_up[59] ;
 wire \ces_3_5_io_outs_up[5] ;
 wire \ces_3_5_io_outs_up[60] ;
 wire \ces_3_5_io_outs_up[61] ;
 wire \ces_3_5_io_outs_up[62] ;
 wire \ces_3_5_io_outs_up[63] ;
 wire \ces_3_5_io_outs_up[6] ;
 wire \ces_3_5_io_outs_up[7] ;
 wire \ces_3_5_io_outs_up[8] ;
 wire \ces_3_5_io_outs_up[9] ;
 wire \ces_3_6_io_ins_down[0] ;
 wire \ces_3_6_io_ins_down[10] ;
 wire \ces_3_6_io_ins_down[11] ;
 wire \ces_3_6_io_ins_down[12] ;
 wire \ces_3_6_io_ins_down[13] ;
 wire \ces_3_6_io_ins_down[14] ;
 wire \ces_3_6_io_ins_down[15] ;
 wire \ces_3_6_io_ins_down[16] ;
 wire \ces_3_6_io_ins_down[17] ;
 wire \ces_3_6_io_ins_down[18] ;
 wire \ces_3_6_io_ins_down[19] ;
 wire \ces_3_6_io_ins_down[1] ;
 wire \ces_3_6_io_ins_down[20] ;
 wire \ces_3_6_io_ins_down[21] ;
 wire \ces_3_6_io_ins_down[22] ;
 wire \ces_3_6_io_ins_down[23] ;
 wire \ces_3_6_io_ins_down[24] ;
 wire \ces_3_6_io_ins_down[25] ;
 wire \ces_3_6_io_ins_down[26] ;
 wire \ces_3_6_io_ins_down[27] ;
 wire \ces_3_6_io_ins_down[28] ;
 wire \ces_3_6_io_ins_down[29] ;
 wire \ces_3_6_io_ins_down[2] ;
 wire \ces_3_6_io_ins_down[30] ;
 wire \ces_3_6_io_ins_down[31] ;
 wire \ces_3_6_io_ins_down[32] ;
 wire \ces_3_6_io_ins_down[33] ;
 wire \ces_3_6_io_ins_down[34] ;
 wire \ces_3_6_io_ins_down[35] ;
 wire \ces_3_6_io_ins_down[36] ;
 wire \ces_3_6_io_ins_down[37] ;
 wire \ces_3_6_io_ins_down[38] ;
 wire \ces_3_6_io_ins_down[39] ;
 wire \ces_3_6_io_ins_down[3] ;
 wire \ces_3_6_io_ins_down[40] ;
 wire \ces_3_6_io_ins_down[41] ;
 wire \ces_3_6_io_ins_down[42] ;
 wire \ces_3_6_io_ins_down[43] ;
 wire \ces_3_6_io_ins_down[44] ;
 wire \ces_3_6_io_ins_down[45] ;
 wire \ces_3_6_io_ins_down[46] ;
 wire \ces_3_6_io_ins_down[47] ;
 wire \ces_3_6_io_ins_down[48] ;
 wire \ces_3_6_io_ins_down[49] ;
 wire \ces_3_6_io_ins_down[4] ;
 wire \ces_3_6_io_ins_down[50] ;
 wire \ces_3_6_io_ins_down[51] ;
 wire \ces_3_6_io_ins_down[52] ;
 wire \ces_3_6_io_ins_down[53] ;
 wire \ces_3_6_io_ins_down[54] ;
 wire \ces_3_6_io_ins_down[55] ;
 wire \ces_3_6_io_ins_down[56] ;
 wire \ces_3_6_io_ins_down[57] ;
 wire \ces_3_6_io_ins_down[58] ;
 wire \ces_3_6_io_ins_down[59] ;
 wire \ces_3_6_io_ins_down[5] ;
 wire \ces_3_6_io_ins_down[60] ;
 wire \ces_3_6_io_ins_down[61] ;
 wire \ces_3_6_io_ins_down[62] ;
 wire \ces_3_6_io_ins_down[63] ;
 wire \ces_3_6_io_ins_down[6] ;
 wire \ces_3_6_io_ins_down[7] ;
 wire \ces_3_6_io_ins_down[8] ;
 wire \ces_3_6_io_ins_down[9] ;
 wire \ces_3_6_io_ins_left[0] ;
 wire \ces_3_6_io_ins_left[10] ;
 wire \ces_3_6_io_ins_left[11] ;
 wire \ces_3_6_io_ins_left[12] ;
 wire \ces_3_6_io_ins_left[13] ;
 wire \ces_3_6_io_ins_left[14] ;
 wire \ces_3_6_io_ins_left[15] ;
 wire \ces_3_6_io_ins_left[16] ;
 wire \ces_3_6_io_ins_left[17] ;
 wire \ces_3_6_io_ins_left[18] ;
 wire \ces_3_6_io_ins_left[19] ;
 wire \ces_3_6_io_ins_left[1] ;
 wire \ces_3_6_io_ins_left[20] ;
 wire \ces_3_6_io_ins_left[21] ;
 wire \ces_3_6_io_ins_left[22] ;
 wire \ces_3_6_io_ins_left[23] ;
 wire \ces_3_6_io_ins_left[24] ;
 wire \ces_3_6_io_ins_left[25] ;
 wire \ces_3_6_io_ins_left[26] ;
 wire \ces_3_6_io_ins_left[27] ;
 wire \ces_3_6_io_ins_left[28] ;
 wire \ces_3_6_io_ins_left[29] ;
 wire \ces_3_6_io_ins_left[2] ;
 wire \ces_3_6_io_ins_left[30] ;
 wire \ces_3_6_io_ins_left[31] ;
 wire \ces_3_6_io_ins_left[32] ;
 wire \ces_3_6_io_ins_left[33] ;
 wire \ces_3_6_io_ins_left[34] ;
 wire \ces_3_6_io_ins_left[35] ;
 wire \ces_3_6_io_ins_left[36] ;
 wire \ces_3_6_io_ins_left[37] ;
 wire \ces_3_6_io_ins_left[38] ;
 wire \ces_3_6_io_ins_left[39] ;
 wire \ces_3_6_io_ins_left[3] ;
 wire \ces_3_6_io_ins_left[40] ;
 wire \ces_3_6_io_ins_left[41] ;
 wire \ces_3_6_io_ins_left[42] ;
 wire \ces_3_6_io_ins_left[43] ;
 wire \ces_3_6_io_ins_left[44] ;
 wire \ces_3_6_io_ins_left[45] ;
 wire \ces_3_6_io_ins_left[46] ;
 wire \ces_3_6_io_ins_left[47] ;
 wire \ces_3_6_io_ins_left[48] ;
 wire \ces_3_6_io_ins_left[49] ;
 wire \ces_3_6_io_ins_left[4] ;
 wire \ces_3_6_io_ins_left[50] ;
 wire \ces_3_6_io_ins_left[51] ;
 wire \ces_3_6_io_ins_left[52] ;
 wire \ces_3_6_io_ins_left[53] ;
 wire \ces_3_6_io_ins_left[54] ;
 wire \ces_3_6_io_ins_left[55] ;
 wire \ces_3_6_io_ins_left[56] ;
 wire \ces_3_6_io_ins_left[57] ;
 wire \ces_3_6_io_ins_left[58] ;
 wire \ces_3_6_io_ins_left[59] ;
 wire \ces_3_6_io_ins_left[5] ;
 wire \ces_3_6_io_ins_left[60] ;
 wire \ces_3_6_io_ins_left[61] ;
 wire \ces_3_6_io_ins_left[62] ;
 wire \ces_3_6_io_ins_left[63] ;
 wire \ces_3_6_io_ins_left[6] ;
 wire \ces_3_6_io_ins_left[7] ;
 wire \ces_3_6_io_ins_left[8] ;
 wire \ces_3_6_io_ins_left[9] ;
 wire ces_3_6_io_lsbOuts_0;
 wire ces_3_6_io_lsbOuts_1;
 wire ces_3_6_io_lsbOuts_2;
 wire ces_3_6_io_lsbOuts_3;
 wire ces_3_6_io_lsbOuts_4;
 wire ces_3_6_io_lsbOuts_5;
 wire ces_3_6_io_lsbOuts_6;
 wire ces_3_6_io_lsbOuts_7;
 wire \ces_3_6_io_outs_right[0] ;
 wire \ces_3_6_io_outs_right[10] ;
 wire \ces_3_6_io_outs_right[11] ;
 wire \ces_3_6_io_outs_right[12] ;
 wire \ces_3_6_io_outs_right[13] ;
 wire \ces_3_6_io_outs_right[14] ;
 wire \ces_3_6_io_outs_right[15] ;
 wire \ces_3_6_io_outs_right[16] ;
 wire \ces_3_6_io_outs_right[17] ;
 wire \ces_3_6_io_outs_right[18] ;
 wire \ces_3_6_io_outs_right[19] ;
 wire \ces_3_6_io_outs_right[1] ;
 wire \ces_3_6_io_outs_right[20] ;
 wire \ces_3_6_io_outs_right[21] ;
 wire \ces_3_6_io_outs_right[22] ;
 wire \ces_3_6_io_outs_right[23] ;
 wire \ces_3_6_io_outs_right[24] ;
 wire \ces_3_6_io_outs_right[25] ;
 wire \ces_3_6_io_outs_right[26] ;
 wire \ces_3_6_io_outs_right[27] ;
 wire \ces_3_6_io_outs_right[28] ;
 wire \ces_3_6_io_outs_right[29] ;
 wire \ces_3_6_io_outs_right[2] ;
 wire \ces_3_6_io_outs_right[30] ;
 wire \ces_3_6_io_outs_right[31] ;
 wire \ces_3_6_io_outs_right[32] ;
 wire \ces_3_6_io_outs_right[33] ;
 wire \ces_3_6_io_outs_right[34] ;
 wire \ces_3_6_io_outs_right[35] ;
 wire \ces_3_6_io_outs_right[36] ;
 wire \ces_3_6_io_outs_right[37] ;
 wire \ces_3_6_io_outs_right[38] ;
 wire \ces_3_6_io_outs_right[39] ;
 wire \ces_3_6_io_outs_right[3] ;
 wire \ces_3_6_io_outs_right[40] ;
 wire \ces_3_6_io_outs_right[41] ;
 wire \ces_3_6_io_outs_right[42] ;
 wire \ces_3_6_io_outs_right[43] ;
 wire \ces_3_6_io_outs_right[44] ;
 wire \ces_3_6_io_outs_right[45] ;
 wire \ces_3_6_io_outs_right[46] ;
 wire \ces_3_6_io_outs_right[47] ;
 wire \ces_3_6_io_outs_right[48] ;
 wire \ces_3_6_io_outs_right[49] ;
 wire \ces_3_6_io_outs_right[4] ;
 wire \ces_3_6_io_outs_right[50] ;
 wire \ces_3_6_io_outs_right[51] ;
 wire \ces_3_6_io_outs_right[52] ;
 wire \ces_3_6_io_outs_right[53] ;
 wire \ces_3_6_io_outs_right[54] ;
 wire \ces_3_6_io_outs_right[55] ;
 wire \ces_3_6_io_outs_right[56] ;
 wire \ces_3_6_io_outs_right[57] ;
 wire \ces_3_6_io_outs_right[58] ;
 wire \ces_3_6_io_outs_right[59] ;
 wire \ces_3_6_io_outs_right[5] ;
 wire \ces_3_6_io_outs_right[60] ;
 wire \ces_3_6_io_outs_right[61] ;
 wire \ces_3_6_io_outs_right[62] ;
 wire \ces_3_6_io_outs_right[63] ;
 wire \ces_3_6_io_outs_right[6] ;
 wire \ces_3_6_io_outs_right[7] ;
 wire \ces_3_6_io_outs_right[8] ;
 wire \ces_3_6_io_outs_right[9] ;
 wire \ces_3_6_io_outs_up[0] ;
 wire \ces_3_6_io_outs_up[10] ;
 wire \ces_3_6_io_outs_up[11] ;
 wire \ces_3_6_io_outs_up[12] ;
 wire \ces_3_6_io_outs_up[13] ;
 wire \ces_3_6_io_outs_up[14] ;
 wire \ces_3_6_io_outs_up[15] ;
 wire \ces_3_6_io_outs_up[16] ;
 wire \ces_3_6_io_outs_up[17] ;
 wire \ces_3_6_io_outs_up[18] ;
 wire \ces_3_6_io_outs_up[19] ;
 wire \ces_3_6_io_outs_up[1] ;
 wire \ces_3_6_io_outs_up[20] ;
 wire \ces_3_6_io_outs_up[21] ;
 wire \ces_3_6_io_outs_up[22] ;
 wire \ces_3_6_io_outs_up[23] ;
 wire \ces_3_6_io_outs_up[24] ;
 wire \ces_3_6_io_outs_up[25] ;
 wire \ces_3_6_io_outs_up[26] ;
 wire \ces_3_6_io_outs_up[27] ;
 wire \ces_3_6_io_outs_up[28] ;
 wire \ces_3_6_io_outs_up[29] ;
 wire \ces_3_6_io_outs_up[2] ;
 wire \ces_3_6_io_outs_up[30] ;
 wire \ces_3_6_io_outs_up[31] ;
 wire \ces_3_6_io_outs_up[32] ;
 wire \ces_3_6_io_outs_up[33] ;
 wire \ces_3_6_io_outs_up[34] ;
 wire \ces_3_6_io_outs_up[35] ;
 wire \ces_3_6_io_outs_up[36] ;
 wire \ces_3_6_io_outs_up[37] ;
 wire \ces_3_6_io_outs_up[38] ;
 wire \ces_3_6_io_outs_up[39] ;
 wire \ces_3_6_io_outs_up[3] ;
 wire \ces_3_6_io_outs_up[40] ;
 wire \ces_3_6_io_outs_up[41] ;
 wire \ces_3_6_io_outs_up[42] ;
 wire \ces_3_6_io_outs_up[43] ;
 wire \ces_3_6_io_outs_up[44] ;
 wire \ces_3_6_io_outs_up[45] ;
 wire \ces_3_6_io_outs_up[46] ;
 wire \ces_3_6_io_outs_up[47] ;
 wire \ces_3_6_io_outs_up[48] ;
 wire \ces_3_6_io_outs_up[49] ;
 wire \ces_3_6_io_outs_up[4] ;
 wire \ces_3_6_io_outs_up[50] ;
 wire \ces_3_6_io_outs_up[51] ;
 wire \ces_3_6_io_outs_up[52] ;
 wire \ces_3_6_io_outs_up[53] ;
 wire \ces_3_6_io_outs_up[54] ;
 wire \ces_3_6_io_outs_up[55] ;
 wire \ces_3_6_io_outs_up[56] ;
 wire \ces_3_6_io_outs_up[57] ;
 wire \ces_3_6_io_outs_up[58] ;
 wire \ces_3_6_io_outs_up[59] ;
 wire \ces_3_6_io_outs_up[5] ;
 wire \ces_3_6_io_outs_up[60] ;
 wire \ces_3_6_io_outs_up[61] ;
 wire \ces_3_6_io_outs_up[62] ;
 wire \ces_3_6_io_outs_up[63] ;
 wire \ces_3_6_io_outs_up[6] ;
 wire \ces_3_6_io_outs_up[7] ;
 wire \ces_3_6_io_outs_up[8] ;
 wire \ces_3_6_io_outs_up[9] ;
 wire \ces_3_7_io_ins_down[0] ;
 wire \ces_3_7_io_ins_down[10] ;
 wire \ces_3_7_io_ins_down[11] ;
 wire \ces_3_7_io_ins_down[12] ;
 wire \ces_3_7_io_ins_down[13] ;
 wire \ces_3_7_io_ins_down[14] ;
 wire \ces_3_7_io_ins_down[15] ;
 wire \ces_3_7_io_ins_down[16] ;
 wire \ces_3_7_io_ins_down[17] ;
 wire \ces_3_7_io_ins_down[18] ;
 wire \ces_3_7_io_ins_down[19] ;
 wire \ces_3_7_io_ins_down[1] ;
 wire \ces_3_7_io_ins_down[20] ;
 wire \ces_3_7_io_ins_down[21] ;
 wire \ces_3_7_io_ins_down[22] ;
 wire \ces_3_7_io_ins_down[23] ;
 wire \ces_3_7_io_ins_down[24] ;
 wire \ces_3_7_io_ins_down[25] ;
 wire \ces_3_7_io_ins_down[26] ;
 wire \ces_3_7_io_ins_down[27] ;
 wire \ces_3_7_io_ins_down[28] ;
 wire \ces_3_7_io_ins_down[29] ;
 wire \ces_3_7_io_ins_down[2] ;
 wire \ces_3_7_io_ins_down[30] ;
 wire \ces_3_7_io_ins_down[31] ;
 wire \ces_3_7_io_ins_down[32] ;
 wire \ces_3_7_io_ins_down[33] ;
 wire \ces_3_7_io_ins_down[34] ;
 wire \ces_3_7_io_ins_down[35] ;
 wire \ces_3_7_io_ins_down[36] ;
 wire \ces_3_7_io_ins_down[37] ;
 wire \ces_3_7_io_ins_down[38] ;
 wire \ces_3_7_io_ins_down[39] ;
 wire \ces_3_7_io_ins_down[3] ;
 wire \ces_3_7_io_ins_down[40] ;
 wire \ces_3_7_io_ins_down[41] ;
 wire \ces_3_7_io_ins_down[42] ;
 wire \ces_3_7_io_ins_down[43] ;
 wire \ces_3_7_io_ins_down[44] ;
 wire \ces_3_7_io_ins_down[45] ;
 wire \ces_3_7_io_ins_down[46] ;
 wire \ces_3_7_io_ins_down[47] ;
 wire \ces_3_7_io_ins_down[48] ;
 wire \ces_3_7_io_ins_down[49] ;
 wire \ces_3_7_io_ins_down[4] ;
 wire \ces_3_7_io_ins_down[50] ;
 wire \ces_3_7_io_ins_down[51] ;
 wire \ces_3_7_io_ins_down[52] ;
 wire \ces_3_7_io_ins_down[53] ;
 wire \ces_3_7_io_ins_down[54] ;
 wire \ces_3_7_io_ins_down[55] ;
 wire \ces_3_7_io_ins_down[56] ;
 wire \ces_3_7_io_ins_down[57] ;
 wire \ces_3_7_io_ins_down[58] ;
 wire \ces_3_7_io_ins_down[59] ;
 wire \ces_3_7_io_ins_down[5] ;
 wire \ces_3_7_io_ins_down[60] ;
 wire \ces_3_7_io_ins_down[61] ;
 wire \ces_3_7_io_ins_down[62] ;
 wire \ces_3_7_io_ins_down[63] ;
 wire \ces_3_7_io_ins_down[6] ;
 wire \ces_3_7_io_ins_down[7] ;
 wire \ces_3_7_io_ins_down[8] ;
 wire \ces_3_7_io_ins_down[9] ;
 wire ces_3_7_io_lsbOuts_0;
 wire ces_3_7_io_lsbOuts_1;
 wire ces_3_7_io_lsbOuts_2;
 wire ces_3_7_io_lsbOuts_3;
 wire ces_3_7_io_lsbOuts_4;
 wire ces_3_7_io_lsbOuts_5;
 wire ces_3_7_io_lsbOuts_6;
 wire ces_3_7_io_lsbOuts_7;
 wire \ces_3_7_io_outs_up[0] ;
 wire \ces_3_7_io_outs_up[10] ;
 wire \ces_3_7_io_outs_up[11] ;
 wire \ces_3_7_io_outs_up[12] ;
 wire \ces_3_7_io_outs_up[13] ;
 wire \ces_3_7_io_outs_up[14] ;
 wire \ces_3_7_io_outs_up[15] ;
 wire \ces_3_7_io_outs_up[16] ;
 wire \ces_3_7_io_outs_up[17] ;
 wire \ces_3_7_io_outs_up[18] ;
 wire \ces_3_7_io_outs_up[19] ;
 wire \ces_3_7_io_outs_up[1] ;
 wire \ces_3_7_io_outs_up[20] ;
 wire \ces_3_7_io_outs_up[21] ;
 wire \ces_3_7_io_outs_up[22] ;
 wire \ces_3_7_io_outs_up[23] ;
 wire \ces_3_7_io_outs_up[24] ;
 wire \ces_3_7_io_outs_up[25] ;
 wire \ces_3_7_io_outs_up[26] ;
 wire \ces_3_7_io_outs_up[27] ;
 wire \ces_3_7_io_outs_up[28] ;
 wire \ces_3_7_io_outs_up[29] ;
 wire \ces_3_7_io_outs_up[2] ;
 wire \ces_3_7_io_outs_up[30] ;
 wire \ces_3_7_io_outs_up[31] ;
 wire \ces_3_7_io_outs_up[32] ;
 wire \ces_3_7_io_outs_up[33] ;
 wire \ces_3_7_io_outs_up[34] ;
 wire \ces_3_7_io_outs_up[35] ;
 wire \ces_3_7_io_outs_up[36] ;
 wire \ces_3_7_io_outs_up[37] ;
 wire \ces_3_7_io_outs_up[38] ;
 wire \ces_3_7_io_outs_up[39] ;
 wire \ces_3_7_io_outs_up[3] ;
 wire \ces_3_7_io_outs_up[40] ;
 wire \ces_3_7_io_outs_up[41] ;
 wire \ces_3_7_io_outs_up[42] ;
 wire \ces_3_7_io_outs_up[43] ;
 wire \ces_3_7_io_outs_up[44] ;
 wire \ces_3_7_io_outs_up[45] ;
 wire \ces_3_7_io_outs_up[46] ;
 wire \ces_3_7_io_outs_up[47] ;
 wire \ces_3_7_io_outs_up[48] ;
 wire \ces_3_7_io_outs_up[49] ;
 wire \ces_3_7_io_outs_up[4] ;
 wire \ces_3_7_io_outs_up[50] ;
 wire \ces_3_7_io_outs_up[51] ;
 wire \ces_3_7_io_outs_up[52] ;
 wire \ces_3_7_io_outs_up[53] ;
 wire \ces_3_7_io_outs_up[54] ;
 wire \ces_3_7_io_outs_up[55] ;
 wire \ces_3_7_io_outs_up[56] ;
 wire \ces_3_7_io_outs_up[57] ;
 wire \ces_3_7_io_outs_up[58] ;
 wire \ces_3_7_io_outs_up[59] ;
 wire \ces_3_7_io_outs_up[5] ;
 wire \ces_3_7_io_outs_up[60] ;
 wire \ces_3_7_io_outs_up[61] ;
 wire \ces_3_7_io_outs_up[62] ;
 wire \ces_3_7_io_outs_up[63] ;
 wire \ces_3_7_io_outs_up[6] ;
 wire \ces_3_7_io_outs_up[7] ;
 wire \ces_3_7_io_outs_up[8] ;
 wire \ces_3_7_io_outs_up[9] ;
 wire \ces_4_0_io_ins_down[0] ;
 wire \ces_4_0_io_ins_down[10] ;
 wire \ces_4_0_io_ins_down[11] ;
 wire \ces_4_0_io_ins_down[12] ;
 wire \ces_4_0_io_ins_down[13] ;
 wire \ces_4_0_io_ins_down[14] ;
 wire \ces_4_0_io_ins_down[15] ;
 wire \ces_4_0_io_ins_down[16] ;
 wire \ces_4_0_io_ins_down[17] ;
 wire \ces_4_0_io_ins_down[18] ;
 wire \ces_4_0_io_ins_down[19] ;
 wire \ces_4_0_io_ins_down[1] ;
 wire \ces_4_0_io_ins_down[20] ;
 wire \ces_4_0_io_ins_down[21] ;
 wire \ces_4_0_io_ins_down[22] ;
 wire \ces_4_0_io_ins_down[23] ;
 wire \ces_4_0_io_ins_down[24] ;
 wire \ces_4_0_io_ins_down[25] ;
 wire \ces_4_0_io_ins_down[26] ;
 wire \ces_4_0_io_ins_down[27] ;
 wire \ces_4_0_io_ins_down[28] ;
 wire \ces_4_0_io_ins_down[29] ;
 wire \ces_4_0_io_ins_down[2] ;
 wire \ces_4_0_io_ins_down[30] ;
 wire \ces_4_0_io_ins_down[31] ;
 wire \ces_4_0_io_ins_down[32] ;
 wire \ces_4_0_io_ins_down[33] ;
 wire \ces_4_0_io_ins_down[34] ;
 wire \ces_4_0_io_ins_down[35] ;
 wire \ces_4_0_io_ins_down[36] ;
 wire \ces_4_0_io_ins_down[37] ;
 wire \ces_4_0_io_ins_down[38] ;
 wire \ces_4_0_io_ins_down[39] ;
 wire \ces_4_0_io_ins_down[3] ;
 wire \ces_4_0_io_ins_down[40] ;
 wire \ces_4_0_io_ins_down[41] ;
 wire \ces_4_0_io_ins_down[42] ;
 wire \ces_4_0_io_ins_down[43] ;
 wire \ces_4_0_io_ins_down[44] ;
 wire \ces_4_0_io_ins_down[45] ;
 wire \ces_4_0_io_ins_down[46] ;
 wire \ces_4_0_io_ins_down[47] ;
 wire \ces_4_0_io_ins_down[48] ;
 wire \ces_4_0_io_ins_down[49] ;
 wire \ces_4_0_io_ins_down[4] ;
 wire \ces_4_0_io_ins_down[50] ;
 wire \ces_4_0_io_ins_down[51] ;
 wire \ces_4_0_io_ins_down[52] ;
 wire \ces_4_0_io_ins_down[53] ;
 wire \ces_4_0_io_ins_down[54] ;
 wire \ces_4_0_io_ins_down[55] ;
 wire \ces_4_0_io_ins_down[56] ;
 wire \ces_4_0_io_ins_down[57] ;
 wire \ces_4_0_io_ins_down[58] ;
 wire \ces_4_0_io_ins_down[59] ;
 wire \ces_4_0_io_ins_down[5] ;
 wire \ces_4_0_io_ins_down[60] ;
 wire \ces_4_0_io_ins_down[61] ;
 wire \ces_4_0_io_ins_down[62] ;
 wire \ces_4_0_io_ins_down[63] ;
 wire \ces_4_0_io_ins_down[6] ;
 wire \ces_4_0_io_ins_down[7] ;
 wire \ces_4_0_io_ins_down[8] ;
 wire \ces_4_0_io_ins_down[9] ;
 wire \ces_4_0_io_ins_left[0] ;
 wire \ces_4_0_io_ins_left[10] ;
 wire \ces_4_0_io_ins_left[11] ;
 wire \ces_4_0_io_ins_left[12] ;
 wire \ces_4_0_io_ins_left[13] ;
 wire \ces_4_0_io_ins_left[14] ;
 wire \ces_4_0_io_ins_left[15] ;
 wire \ces_4_0_io_ins_left[16] ;
 wire \ces_4_0_io_ins_left[17] ;
 wire \ces_4_0_io_ins_left[18] ;
 wire \ces_4_0_io_ins_left[19] ;
 wire \ces_4_0_io_ins_left[1] ;
 wire \ces_4_0_io_ins_left[20] ;
 wire \ces_4_0_io_ins_left[21] ;
 wire \ces_4_0_io_ins_left[22] ;
 wire \ces_4_0_io_ins_left[23] ;
 wire \ces_4_0_io_ins_left[24] ;
 wire \ces_4_0_io_ins_left[25] ;
 wire \ces_4_0_io_ins_left[26] ;
 wire \ces_4_0_io_ins_left[27] ;
 wire \ces_4_0_io_ins_left[28] ;
 wire \ces_4_0_io_ins_left[29] ;
 wire \ces_4_0_io_ins_left[2] ;
 wire \ces_4_0_io_ins_left[30] ;
 wire \ces_4_0_io_ins_left[31] ;
 wire \ces_4_0_io_ins_left[32] ;
 wire \ces_4_0_io_ins_left[33] ;
 wire \ces_4_0_io_ins_left[34] ;
 wire \ces_4_0_io_ins_left[35] ;
 wire \ces_4_0_io_ins_left[36] ;
 wire \ces_4_0_io_ins_left[37] ;
 wire \ces_4_0_io_ins_left[38] ;
 wire \ces_4_0_io_ins_left[39] ;
 wire \ces_4_0_io_ins_left[3] ;
 wire \ces_4_0_io_ins_left[40] ;
 wire \ces_4_0_io_ins_left[41] ;
 wire \ces_4_0_io_ins_left[42] ;
 wire \ces_4_0_io_ins_left[43] ;
 wire \ces_4_0_io_ins_left[44] ;
 wire \ces_4_0_io_ins_left[45] ;
 wire \ces_4_0_io_ins_left[46] ;
 wire \ces_4_0_io_ins_left[47] ;
 wire \ces_4_0_io_ins_left[48] ;
 wire \ces_4_0_io_ins_left[49] ;
 wire \ces_4_0_io_ins_left[4] ;
 wire \ces_4_0_io_ins_left[50] ;
 wire \ces_4_0_io_ins_left[51] ;
 wire \ces_4_0_io_ins_left[52] ;
 wire \ces_4_0_io_ins_left[53] ;
 wire \ces_4_0_io_ins_left[54] ;
 wire \ces_4_0_io_ins_left[55] ;
 wire \ces_4_0_io_ins_left[56] ;
 wire \ces_4_0_io_ins_left[57] ;
 wire \ces_4_0_io_ins_left[58] ;
 wire \ces_4_0_io_ins_left[59] ;
 wire \ces_4_0_io_ins_left[5] ;
 wire \ces_4_0_io_ins_left[60] ;
 wire \ces_4_0_io_ins_left[61] ;
 wire \ces_4_0_io_ins_left[62] ;
 wire \ces_4_0_io_ins_left[63] ;
 wire \ces_4_0_io_ins_left[6] ;
 wire \ces_4_0_io_ins_left[7] ;
 wire \ces_4_0_io_ins_left[8] ;
 wire \ces_4_0_io_ins_left[9] ;
 wire ces_4_0_io_lsbOuts_0;
 wire ces_4_0_io_lsbOuts_1;
 wire ces_4_0_io_lsbOuts_2;
 wire ces_4_0_io_lsbOuts_3;
 wire ces_4_0_io_lsbOuts_4;
 wire ces_4_0_io_lsbOuts_5;
 wire ces_4_0_io_lsbOuts_6;
 wire ces_4_0_io_lsbOuts_7;
 wire \ces_4_0_io_outs_right[0] ;
 wire \ces_4_0_io_outs_right[10] ;
 wire \ces_4_0_io_outs_right[11] ;
 wire \ces_4_0_io_outs_right[12] ;
 wire \ces_4_0_io_outs_right[13] ;
 wire \ces_4_0_io_outs_right[14] ;
 wire \ces_4_0_io_outs_right[15] ;
 wire \ces_4_0_io_outs_right[16] ;
 wire \ces_4_0_io_outs_right[17] ;
 wire \ces_4_0_io_outs_right[18] ;
 wire \ces_4_0_io_outs_right[19] ;
 wire \ces_4_0_io_outs_right[1] ;
 wire \ces_4_0_io_outs_right[20] ;
 wire \ces_4_0_io_outs_right[21] ;
 wire \ces_4_0_io_outs_right[22] ;
 wire \ces_4_0_io_outs_right[23] ;
 wire \ces_4_0_io_outs_right[24] ;
 wire \ces_4_0_io_outs_right[25] ;
 wire \ces_4_0_io_outs_right[26] ;
 wire \ces_4_0_io_outs_right[27] ;
 wire \ces_4_0_io_outs_right[28] ;
 wire \ces_4_0_io_outs_right[29] ;
 wire \ces_4_0_io_outs_right[2] ;
 wire \ces_4_0_io_outs_right[30] ;
 wire \ces_4_0_io_outs_right[31] ;
 wire \ces_4_0_io_outs_right[32] ;
 wire \ces_4_0_io_outs_right[33] ;
 wire \ces_4_0_io_outs_right[34] ;
 wire \ces_4_0_io_outs_right[35] ;
 wire \ces_4_0_io_outs_right[36] ;
 wire \ces_4_0_io_outs_right[37] ;
 wire \ces_4_0_io_outs_right[38] ;
 wire \ces_4_0_io_outs_right[39] ;
 wire \ces_4_0_io_outs_right[3] ;
 wire \ces_4_0_io_outs_right[40] ;
 wire \ces_4_0_io_outs_right[41] ;
 wire \ces_4_0_io_outs_right[42] ;
 wire \ces_4_0_io_outs_right[43] ;
 wire \ces_4_0_io_outs_right[44] ;
 wire \ces_4_0_io_outs_right[45] ;
 wire \ces_4_0_io_outs_right[46] ;
 wire \ces_4_0_io_outs_right[47] ;
 wire \ces_4_0_io_outs_right[48] ;
 wire \ces_4_0_io_outs_right[49] ;
 wire \ces_4_0_io_outs_right[4] ;
 wire \ces_4_0_io_outs_right[50] ;
 wire \ces_4_0_io_outs_right[51] ;
 wire \ces_4_0_io_outs_right[52] ;
 wire \ces_4_0_io_outs_right[53] ;
 wire \ces_4_0_io_outs_right[54] ;
 wire \ces_4_0_io_outs_right[55] ;
 wire \ces_4_0_io_outs_right[56] ;
 wire \ces_4_0_io_outs_right[57] ;
 wire \ces_4_0_io_outs_right[58] ;
 wire \ces_4_0_io_outs_right[59] ;
 wire \ces_4_0_io_outs_right[5] ;
 wire \ces_4_0_io_outs_right[60] ;
 wire \ces_4_0_io_outs_right[61] ;
 wire \ces_4_0_io_outs_right[62] ;
 wire \ces_4_0_io_outs_right[63] ;
 wire \ces_4_0_io_outs_right[6] ;
 wire \ces_4_0_io_outs_right[7] ;
 wire \ces_4_0_io_outs_right[8] ;
 wire \ces_4_0_io_outs_right[9] ;
 wire \ces_4_0_io_outs_up[0] ;
 wire \ces_4_0_io_outs_up[10] ;
 wire \ces_4_0_io_outs_up[11] ;
 wire \ces_4_0_io_outs_up[12] ;
 wire \ces_4_0_io_outs_up[13] ;
 wire \ces_4_0_io_outs_up[14] ;
 wire \ces_4_0_io_outs_up[15] ;
 wire \ces_4_0_io_outs_up[16] ;
 wire \ces_4_0_io_outs_up[17] ;
 wire \ces_4_0_io_outs_up[18] ;
 wire \ces_4_0_io_outs_up[19] ;
 wire \ces_4_0_io_outs_up[1] ;
 wire \ces_4_0_io_outs_up[20] ;
 wire \ces_4_0_io_outs_up[21] ;
 wire \ces_4_0_io_outs_up[22] ;
 wire \ces_4_0_io_outs_up[23] ;
 wire \ces_4_0_io_outs_up[24] ;
 wire \ces_4_0_io_outs_up[25] ;
 wire \ces_4_0_io_outs_up[26] ;
 wire \ces_4_0_io_outs_up[27] ;
 wire \ces_4_0_io_outs_up[28] ;
 wire \ces_4_0_io_outs_up[29] ;
 wire \ces_4_0_io_outs_up[2] ;
 wire \ces_4_0_io_outs_up[30] ;
 wire \ces_4_0_io_outs_up[31] ;
 wire \ces_4_0_io_outs_up[32] ;
 wire \ces_4_0_io_outs_up[33] ;
 wire \ces_4_0_io_outs_up[34] ;
 wire \ces_4_0_io_outs_up[35] ;
 wire \ces_4_0_io_outs_up[36] ;
 wire \ces_4_0_io_outs_up[37] ;
 wire \ces_4_0_io_outs_up[38] ;
 wire \ces_4_0_io_outs_up[39] ;
 wire \ces_4_0_io_outs_up[3] ;
 wire \ces_4_0_io_outs_up[40] ;
 wire \ces_4_0_io_outs_up[41] ;
 wire \ces_4_0_io_outs_up[42] ;
 wire \ces_4_0_io_outs_up[43] ;
 wire \ces_4_0_io_outs_up[44] ;
 wire \ces_4_0_io_outs_up[45] ;
 wire \ces_4_0_io_outs_up[46] ;
 wire \ces_4_0_io_outs_up[47] ;
 wire \ces_4_0_io_outs_up[48] ;
 wire \ces_4_0_io_outs_up[49] ;
 wire \ces_4_0_io_outs_up[4] ;
 wire \ces_4_0_io_outs_up[50] ;
 wire \ces_4_0_io_outs_up[51] ;
 wire \ces_4_0_io_outs_up[52] ;
 wire \ces_4_0_io_outs_up[53] ;
 wire \ces_4_0_io_outs_up[54] ;
 wire \ces_4_0_io_outs_up[55] ;
 wire \ces_4_0_io_outs_up[56] ;
 wire \ces_4_0_io_outs_up[57] ;
 wire \ces_4_0_io_outs_up[58] ;
 wire \ces_4_0_io_outs_up[59] ;
 wire \ces_4_0_io_outs_up[5] ;
 wire \ces_4_0_io_outs_up[60] ;
 wire \ces_4_0_io_outs_up[61] ;
 wire \ces_4_0_io_outs_up[62] ;
 wire \ces_4_0_io_outs_up[63] ;
 wire \ces_4_0_io_outs_up[6] ;
 wire \ces_4_0_io_outs_up[7] ;
 wire \ces_4_0_io_outs_up[8] ;
 wire \ces_4_0_io_outs_up[9] ;
 wire \ces_4_1_io_ins_down[0] ;
 wire \ces_4_1_io_ins_down[10] ;
 wire \ces_4_1_io_ins_down[11] ;
 wire \ces_4_1_io_ins_down[12] ;
 wire \ces_4_1_io_ins_down[13] ;
 wire \ces_4_1_io_ins_down[14] ;
 wire \ces_4_1_io_ins_down[15] ;
 wire \ces_4_1_io_ins_down[16] ;
 wire \ces_4_1_io_ins_down[17] ;
 wire \ces_4_1_io_ins_down[18] ;
 wire \ces_4_1_io_ins_down[19] ;
 wire \ces_4_1_io_ins_down[1] ;
 wire \ces_4_1_io_ins_down[20] ;
 wire \ces_4_1_io_ins_down[21] ;
 wire \ces_4_1_io_ins_down[22] ;
 wire \ces_4_1_io_ins_down[23] ;
 wire \ces_4_1_io_ins_down[24] ;
 wire \ces_4_1_io_ins_down[25] ;
 wire \ces_4_1_io_ins_down[26] ;
 wire \ces_4_1_io_ins_down[27] ;
 wire \ces_4_1_io_ins_down[28] ;
 wire \ces_4_1_io_ins_down[29] ;
 wire \ces_4_1_io_ins_down[2] ;
 wire \ces_4_1_io_ins_down[30] ;
 wire \ces_4_1_io_ins_down[31] ;
 wire \ces_4_1_io_ins_down[32] ;
 wire \ces_4_1_io_ins_down[33] ;
 wire \ces_4_1_io_ins_down[34] ;
 wire \ces_4_1_io_ins_down[35] ;
 wire \ces_4_1_io_ins_down[36] ;
 wire \ces_4_1_io_ins_down[37] ;
 wire \ces_4_1_io_ins_down[38] ;
 wire \ces_4_1_io_ins_down[39] ;
 wire \ces_4_1_io_ins_down[3] ;
 wire \ces_4_1_io_ins_down[40] ;
 wire \ces_4_1_io_ins_down[41] ;
 wire \ces_4_1_io_ins_down[42] ;
 wire \ces_4_1_io_ins_down[43] ;
 wire \ces_4_1_io_ins_down[44] ;
 wire \ces_4_1_io_ins_down[45] ;
 wire \ces_4_1_io_ins_down[46] ;
 wire \ces_4_1_io_ins_down[47] ;
 wire \ces_4_1_io_ins_down[48] ;
 wire \ces_4_1_io_ins_down[49] ;
 wire \ces_4_1_io_ins_down[4] ;
 wire \ces_4_1_io_ins_down[50] ;
 wire \ces_4_1_io_ins_down[51] ;
 wire \ces_4_1_io_ins_down[52] ;
 wire \ces_4_1_io_ins_down[53] ;
 wire \ces_4_1_io_ins_down[54] ;
 wire \ces_4_1_io_ins_down[55] ;
 wire \ces_4_1_io_ins_down[56] ;
 wire \ces_4_1_io_ins_down[57] ;
 wire \ces_4_1_io_ins_down[58] ;
 wire \ces_4_1_io_ins_down[59] ;
 wire \ces_4_1_io_ins_down[5] ;
 wire \ces_4_1_io_ins_down[60] ;
 wire \ces_4_1_io_ins_down[61] ;
 wire \ces_4_1_io_ins_down[62] ;
 wire \ces_4_1_io_ins_down[63] ;
 wire \ces_4_1_io_ins_down[6] ;
 wire \ces_4_1_io_ins_down[7] ;
 wire \ces_4_1_io_ins_down[8] ;
 wire \ces_4_1_io_ins_down[9] ;
 wire \ces_4_1_io_ins_left[0] ;
 wire \ces_4_1_io_ins_left[10] ;
 wire \ces_4_1_io_ins_left[11] ;
 wire \ces_4_1_io_ins_left[12] ;
 wire \ces_4_1_io_ins_left[13] ;
 wire \ces_4_1_io_ins_left[14] ;
 wire \ces_4_1_io_ins_left[15] ;
 wire \ces_4_1_io_ins_left[16] ;
 wire \ces_4_1_io_ins_left[17] ;
 wire \ces_4_1_io_ins_left[18] ;
 wire \ces_4_1_io_ins_left[19] ;
 wire \ces_4_1_io_ins_left[1] ;
 wire \ces_4_1_io_ins_left[20] ;
 wire \ces_4_1_io_ins_left[21] ;
 wire \ces_4_1_io_ins_left[22] ;
 wire \ces_4_1_io_ins_left[23] ;
 wire \ces_4_1_io_ins_left[24] ;
 wire \ces_4_1_io_ins_left[25] ;
 wire \ces_4_1_io_ins_left[26] ;
 wire \ces_4_1_io_ins_left[27] ;
 wire \ces_4_1_io_ins_left[28] ;
 wire \ces_4_1_io_ins_left[29] ;
 wire \ces_4_1_io_ins_left[2] ;
 wire \ces_4_1_io_ins_left[30] ;
 wire \ces_4_1_io_ins_left[31] ;
 wire \ces_4_1_io_ins_left[32] ;
 wire \ces_4_1_io_ins_left[33] ;
 wire \ces_4_1_io_ins_left[34] ;
 wire \ces_4_1_io_ins_left[35] ;
 wire \ces_4_1_io_ins_left[36] ;
 wire \ces_4_1_io_ins_left[37] ;
 wire \ces_4_1_io_ins_left[38] ;
 wire \ces_4_1_io_ins_left[39] ;
 wire \ces_4_1_io_ins_left[3] ;
 wire \ces_4_1_io_ins_left[40] ;
 wire \ces_4_1_io_ins_left[41] ;
 wire \ces_4_1_io_ins_left[42] ;
 wire \ces_4_1_io_ins_left[43] ;
 wire \ces_4_1_io_ins_left[44] ;
 wire \ces_4_1_io_ins_left[45] ;
 wire \ces_4_1_io_ins_left[46] ;
 wire \ces_4_1_io_ins_left[47] ;
 wire \ces_4_1_io_ins_left[48] ;
 wire \ces_4_1_io_ins_left[49] ;
 wire \ces_4_1_io_ins_left[4] ;
 wire \ces_4_1_io_ins_left[50] ;
 wire \ces_4_1_io_ins_left[51] ;
 wire \ces_4_1_io_ins_left[52] ;
 wire \ces_4_1_io_ins_left[53] ;
 wire \ces_4_1_io_ins_left[54] ;
 wire \ces_4_1_io_ins_left[55] ;
 wire \ces_4_1_io_ins_left[56] ;
 wire \ces_4_1_io_ins_left[57] ;
 wire \ces_4_1_io_ins_left[58] ;
 wire \ces_4_1_io_ins_left[59] ;
 wire \ces_4_1_io_ins_left[5] ;
 wire \ces_4_1_io_ins_left[60] ;
 wire \ces_4_1_io_ins_left[61] ;
 wire \ces_4_1_io_ins_left[62] ;
 wire \ces_4_1_io_ins_left[63] ;
 wire \ces_4_1_io_ins_left[6] ;
 wire \ces_4_1_io_ins_left[7] ;
 wire \ces_4_1_io_ins_left[8] ;
 wire \ces_4_1_io_ins_left[9] ;
 wire ces_4_1_io_lsbOuts_0;
 wire ces_4_1_io_lsbOuts_1;
 wire ces_4_1_io_lsbOuts_2;
 wire ces_4_1_io_lsbOuts_3;
 wire ces_4_1_io_lsbOuts_4;
 wire ces_4_1_io_lsbOuts_5;
 wire ces_4_1_io_lsbOuts_6;
 wire ces_4_1_io_lsbOuts_7;
 wire \ces_4_1_io_outs_right[0] ;
 wire \ces_4_1_io_outs_right[10] ;
 wire \ces_4_1_io_outs_right[11] ;
 wire \ces_4_1_io_outs_right[12] ;
 wire \ces_4_1_io_outs_right[13] ;
 wire \ces_4_1_io_outs_right[14] ;
 wire \ces_4_1_io_outs_right[15] ;
 wire \ces_4_1_io_outs_right[16] ;
 wire \ces_4_1_io_outs_right[17] ;
 wire \ces_4_1_io_outs_right[18] ;
 wire \ces_4_1_io_outs_right[19] ;
 wire \ces_4_1_io_outs_right[1] ;
 wire \ces_4_1_io_outs_right[20] ;
 wire \ces_4_1_io_outs_right[21] ;
 wire \ces_4_1_io_outs_right[22] ;
 wire \ces_4_1_io_outs_right[23] ;
 wire \ces_4_1_io_outs_right[24] ;
 wire \ces_4_1_io_outs_right[25] ;
 wire \ces_4_1_io_outs_right[26] ;
 wire \ces_4_1_io_outs_right[27] ;
 wire \ces_4_1_io_outs_right[28] ;
 wire \ces_4_1_io_outs_right[29] ;
 wire \ces_4_1_io_outs_right[2] ;
 wire \ces_4_1_io_outs_right[30] ;
 wire \ces_4_1_io_outs_right[31] ;
 wire \ces_4_1_io_outs_right[32] ;
 wire \ces_4_1_io_outs_right[33] ;
 wire \ces_4_1_io_outs_right[34] ;
 wire \ces_4_1_io_outs_right[35] ;
 wire \ces_4_1_io_outs_right[36] ;
 wire \ces_4_1_io_outs_right[37] ;
 wire \ces_4_1_io_outs_right[38] ;
 wire \ces_4_1_io_outs_right[39] ;
 wire \ces_4_1_io_outs_right[3] ;
 wire \ces_4_1_io_outs_right[40] ;
 wire \ces_4_1_io_outs_right[41] ;
 wire \ces_4_1_io_outs_right[42] ;
 wire \ces_4_1_io_outs_right[43] ;
 wire \ces_4_1_io_outs_right[44] ;
 wire \ces_4_1_io_outs_right[45] ;
 wire \ces_4_1_io_outs_right[46] ;
 wire \ces_4_1_io_outs_right[47] ;
 wire \ces_4_1_io_outs_right[48] ;
 wire \ces_4_1_io_outs_right[49] ;
 wire \ces_4_1_io_outs_right[4] ;
 wire \ces_4_1_io_outs_right[50] ;
 wire \ces_4_1_io_outs_right[51] ;
 wire \ces_4_1_io_outs_right[52] ;
 wire \ces_4_1_io_outs_right[53] ;
 wire \ces_4_1_io_outs_right[54] ;
 wire \ces_4_1_io_outs_right[55] ;
 wire \ces_4_1_io_outs_right[56] ;
 wire \ces_4_1_io_outs_right[57] ;
 wire \ces_4_1_io_outs_right[58] ;
 wire \ces_4_1_io_outs_right[59] ;
 wire \ces_4_1_io_outs_right[5] ;
 wire \ces_4_1_io_outs_right[60] ;
 wire \ces_4_1_io_outs_right[61] ;
 wire \ces_4_1_io_outs_right[62] ;
 wire \ces_4_1_io_outs_right[63] ;
 wire \ces_4_1_io_outs_right[6] ;
 wire \ces_4_1_io_outs_right[7] ;
 wire \ces_4_1_io_outs_right[8] ;
 wire \ces_4_1_io_outs_right[9] ;
 wire \ces_4_1_io_outs_up[0] ;
 wire \ces_4_1_io_outs_up[10] ;
 wire \ces_4_1_io_outs_up[11] ;
 wire \ces_4_1_io_outs_up[12] ;
 wire \ces_4_1_io_outs_up[13] ;
 wire \ces_4_1_io_outs_up[14] ;
 wire \ces_4_1_io_outs_up[15] ;
 wire \ces_4_1_io_outs_up[16] ;
 wire \ces_4_1_io_outs_up[17] ;
 wire \ces_4_1_io_outs_up[18] ;
 wire \ces_4_1_io_outs_up[19] ;
 wire \ces_4_1_io_outs_up[1] ;
 wire \ces_4_1_io_outs_up[20] ;
 wire \ces_4_1_io_outs_up[21] ;
 wire \ces_4_1_io_outs_up[22] ;
 wire \ces_4_1_io_outs_up[23] ;
 wire \ces_4_1_io_outs_up[24] ;
 wire \ces_4_1_io_outs_up[25] ;
 wire \ces_4_1_io_outs_up[26] ;
 wire \ces_4_1_io_outs_up[27] ;
 wire \ces_4_1_io_outs_up[28] ;
 wire \ces_4_1_io_outs_up[29] ;
 wire \ces_4_1_io_outs_up[2] ;
 wire \ces_4_1_io_outs_up[30] ;
 wire \ces_4_1_io_outs_up[31] ;
 wire \ces_4_1_io_outs_up[32] ;
 wire \ces_4_1_io_outs_up[33] ;
 wire \ces_4_1_io_outs_up[34] ;
 wire \ces_4_1_io_outs_up[35] ;
 wire \ces_4_1_io_outs_up[36] ;
 wire \ces_4_1_io_outs_up[37] ;
 wire \ces_4_1_io_outs_up[38] ;
 wire \ces_4_1_io_outs_up[39] ;
 wire \ces_4_1_io_outs_up[3] ;
 wire \ces_4_1_io_outs_up[40] ;
 wire \ces_4_1_io_outs_up[41] ;
 wire \ces_4_1_io_outs_up[42] ;
 wire \ces_4_1_io_outs_up[43] ;
 wire \ces_4_1_io_outs_up[44] ;
 wire \ces_4_1_io_outs_up[45] ;
 wire \ces_4_1_io_outs_up[46] ;
 wire \ces_4_1_io_outs_up[47] ;
 wire \ces_4_1_io_outs_up[48] ;
 wire \ces_4_1_io_outs_up[49] ;
 wire \ces_4_1_io_outs_up[4] ;
 wire \ces_4_1_io_outs_up[50] ;
 wire \ces_4_1_io_outs_up[51] ;
 wire \ces_4_1_io_outs_up[52] ;
 wire \ces_4_1_io_outs_up[53] ;
 wire \ces_4_1_io_outs_up[54] ;
 wire \ces_4_1_io_outs_up[55] ;
 wire \ces_4_1_io_outs_up[56] ;
 wire \ces_4_1_io_outs_up[57] ;
 wire \ces_4_1_io_outs_up[58] ;
 wire \ces_4_1_io_outs_up[59] ;
 wire \ces_4_1_io_outs_up[5] ;
 wire \ces_4_1_io_outs_up[60] ;
 wire \ces_4_1_io_outs_up[61] ;
 wire \ces_4_1_io_outs_up[62] ;
 wire \ces_4_1_io_outs_up[63] ;
 wire \ces_4_1_io_outs_up[6] ;
 wire \ces_4_1_io_outs_up[7] ;
 wire \ces_4_1_io_outs_up[8] ;
 wire \ces_4_1_io_outs_up[9] ;
 wire \ces_4_2_io_ins_down[0] ;
 wire \ces_4_2_io_ins_down[10] ;
 wire \ces_4_2_io_ins_down[11] ;
 wire \ces_4_2_io_ins_down[12] ;
 wire \ces_4_2_io_ins_down[13] ;
 wire \ces_4_2_io_ins_down[14] ;
 wire \ces_4_2_io_ins_down[15] ;
 wire \ces_4_2_io_ins_down[16] ;
 wire \ces_4_2_io_ins_down[17] ;
 wire \ces_4_2_io_ins_down[18] ;
 wire \ces_4_2_io_ins_down[19] ;
 wire \ces_4_2_io_ins_down[1] ;
 wire \ces_4_2_io_ins_down[20] ;
 wire \ces_4_2_io_ins_down[21] ;
 wire \ces_4_2_io_ins_down[22] ;
 wire \ces_4_2_io_ins_down[23] ;
 wire \ces_4_2_io_ins_down[24] ;
 wire \ces_4_2_io_ins_down[25] ;
 wire \ces_4_2_io_ins_down[26] ;
 wire \ces_4_2_io_ins_down[27] ;
 wire \ces_4_2_io_ins_down[28] ;
 wire \ces_4_2_io_ins_down[29] ;
 wire \ces_4_2_io_ins_down[2] ;
 wire \ces_4_2_io_ins_down[30] ;
 wire \ces_4_2_io_ins_down[31] ;
 wire \ces_4_2_io_ins_down[32] ;
 wire \ces_4_2_io_ins_down[33] ;
 wire \ces_4_2_io_ins_down[34] ;
 wire \ces_4_2_io_ins_down[35] ;
 wire \ces_4_2_io_ins_down[36] ;
 wire \ces_4_2_io_ins_down[37] ;
 wire \ces_4_2_io_ins_down[38] ;
 wire \ces_4_2_io_ins_down[39] ;
 wire \ces_4_2_io_ins_down[3] ;
 wire \ces_4_2_io_ins_down[40] ;
 wire \ces_4_2_io_ins_down[41] ;
 wire \ces_4_2_io_ins_down[42] ;
 wire \ces_4_2_io_ins_down[43] ;
 wire \ces_4_2_io_ins_down[44] ;
 wire \ces_4_2_io_ins_down[45] ;
 wire \ces_4_2_io_ins_down[46] ;
 wire \ces_4_2_io_ins_down[47] ;
 wire \ces_4_2_io_ins_down[48] ;
 wire \ces_4_2_io_ins_down[49] ;
 wire \ces_4_2_io_ins_down[4] ;
 wire \ces_4_2_io_ins_down[50] ;
 wire \ces_4_2_io_ins_down[51] ;
 wire \ces_4_2_io_ins_down[52] ;
 wire \ces_4_2_io_ins_down[53] ;
 wire \ces_4_2_io_ins_down[54] ;
 wire \ces_4_2_io_ins_down[55] ;
 wire \ces_4_2_io_ins_down[56] ;
 wire \ces_4_2_io_ins_down[57] ;
 wire \ces_4_2_io_ins_down[58] ;
 wire \ces_4_2_io_ins_down[59] ;
 wire \ces_4_2_io_ins_down[5] ;
 wire \ces_4_2_io_ins_down[60] ;
 wire \ces_4_2_io_ins_down[61] ;
 wire \ces_4_2_io_ins_down[62] ;
 wire \ces_4_2_io_ins_down[63] ;
 wire \ces_4_2_io_ins_down[6] ;
 wire \ces_4_2_io_ins_down[7] ;
 wire \ces_4_2_io_ins_down[8] ;
 wire \ces_4_2_io_ins_down[9] ;
 wire \ces_4_2_io_ins_left[0] ;
 wire \ces_4_2_io_ins_left[10] ;
 wire \ces_4_2_io_ins_left[11] ;
 wire \ces_4_2_io_ins_left[12] ;
 wire \ces_4_2_io_ins_left[13] ;
 wire \ces_4_2_io_ins_left[14] ;
 wire \ces_4_2_io_ins_left[15] ;
 wire \ces_4_2_io_ins_left[16] ;
 wire \ces_4_2_io_ins_left[17] ;
 wire \ces_4_2_io_ins_left[18] ;
 wire \ces_4_2_io_ins_left[19] ;
 wire \ces_4_2_io_ins_left[1] ;
 wire \ces_4_2_io_ins_left[20] ;
 wire \ces_4_2_io_ins_left[21] ;
 wire \ces_4_2_io_ins_left[22] ;
 wire \ces_4_2_io_ins_left[23] ;
 wire \ces_4_2_io_ins_left[24] ;
 wire \ces_4_2_io_ins_left[25] ;
 wire \ces_4_2_io_ins_left[26] ;
 wire \ces_4_2_io_ins_left[27] ;
 wire \ces_4_2_io_ins_left[28] ;
 wire \ces_4_2_io_ins_left[29] ;
 wire \ces_4_2_io_ins_left[2] ;
 wire \ces_4_2_io_ins_left[30] ;
 wire \ces_4_2_io_ins_left[31] ;
 wire \ces_4_2_io_ins_left[32] ;
 wire \ces_4_2_io_ins_left[33] ;
 wire \ces_4_2_io_ins_left[34] ;
 wire \ces_4_2_io_ins_left[35] ;
 wire \ces_4_2_io_ins_left[36] ;
 wire \ces_4_2_io_ins_left[37] ;
 wire \ces_4_2_io_ins_left[38] ;
 wire \ces_4_2_io_ins_left[39] ;
 wire \ces_4_2_io_ins_left[3] ;
 wire \ces_4_2_io_ins_left[40] ;
 wire \ces_4_2_io_ins_left[41] ;
 wire \ces_4_2_io_ins_left[42] ;
 wire \ces_4_2_io_ins_left[43] ;
 wire \ces_4_2_io_ins_left[44] ;
 wire \ces_4_2_io_ins_left[45] ;
 wire \ces_4_2_io_ins_left[46] ;
 wire \ces_4_2_io_ins_left[47] ;
 wire \ces_4_2_io_ins_left[48] ;
 wire \ces_4_2_io_ins_left[49] ;
 wire \ces_4_2_io_ins_left[4] ;
 wire \ces_4_2_io_ins_left[50] ;
 wire \ces_4_2_io_ins_left[51] ;
 wire \ces_4_2_io_ins_left[52] ;
 wire \ces_4_2_io_ins_left[53] ;
 wire \ces_4_2_io_ins_left[54] ;
 wire \ces_4_2_io_ins_left[55] ;
 wire \ces_4_2_io_ins_left[56] ;
 wire \ces_4_2_io_ins_left[57] ;
 wire \ces_4_2_io_ins_left[58] ;
 wire \ces_4_2_io_ins_left[59] ;
 wire \ces_4_2_io_ins_left[5] ;
 wire \ces_4_2_io_ins_left[60] ;
 wire \ces_4_2_io_ins_left[61] ;
 wire \ces_4_2_io_ins_left[62] ;
 wire \ces_4_2_io_ins_left[63] ;
 wire \ces_4_2_io_ins_left[6] ;
 wire \ces_4_2_io_ins_left[7] ;
 wire \ces_4_2_io_ins_left[8] ;
 wire \ces_4_2_io_ins_left[9] ;
 wire ces_4_2_io_lsbOuts_0;
 wire ces_4_2_io_lsbOuts_1;
 wire ces_4_2_io_lsbOuts_2;
 wire ces_4_2_io_lsbOuts_3;
 wire ces_4_2_io_lsbOuts_4;
 wire ces_4_2_io_lsbOuts_5;
 wire ces_4_2_io_lsbOuts_6;
 wire ces_4_2_io_lsbOuts_7;
 wire \ces_4_2_io_outs_right[0] ;
 wire \ces_4_2_io_outs_right[10] ;
 wire \ces_4_2_io_outs_right[11] ;
 wire \ces_4_2_io_outs_right[12] ;
 wire \ces_4_2_io_outs_right[13] ;
 wire \ces_4_2_io_outs_right[14] ;
 wire \ces_4_2_io_outs_right[15] ;
 wire \ces_4_2_io_outs_right[16] ;
 wire \ces_4_2_io_outs_right[17] ;
 wire \ces_4_2_io_outs_right[18] ;
 wire \ces_4_2_io_outs_right[19] ;
 wire \ces_4_2_io_outs_right[1] ;
 wire \ces_4_2_io_outs_right[20] ;
 wire \ces_4_2_io_outs_right[21] ;
 wire \ces_4_2_io_outs_right[22] ;
 wire \ces_4_2_io_outs_right[23] ;
 wire \ces_4_2_io_outs_right[24] ;
 wire \ces_4_2_io_outs_right[25] ;
 wire \ces_4_2_io_outs_right[26] ;
 wire \ces_4_2_io_outs_right[27] ;
 wire \ces_4_2_io_outs_right[28] ;
 wire \ces_4_2_io_outs_right[29] ;
 wire \ces_4_2_io_outs_right[2] ;
 wire \ces_4_2_io_outs_right[30] ;
 wire \ces_4_2_io_outs_right[31] ;
 wire \ces_4_2_io_outs_right[32] ;
 wire \ces_4_2_io_outs_right[33] ;
 wire \ces_4_2_io_outs_right[34] ;
 wire \ces_4_2_io_outs_right[35] ;
 wire \ces_4_2_io_outs_right[36] ;
 wire \ces_4_2_io_outs_right[37] ;
 wire \ces_4_2_io_outs_right[38] ;
 wire \ces_4_2_io_outs_right[39] ;
 wire \ces_4_2_io_outs_right[3] ;
 wire \ces_4_2_io_outs_right[40] ;
 wire \ces_4_2_io_outs_right[41] ;
 wire \ces_4_2_io_outs_right[42] ;
 wire \ces_4_2_io_outs_right[43] ;
 wire \ces_4_2_io_outs_right[44] ;
 wire \ces_4_2_io_outs_right[45] ;
 wire \ces_4_2_io_outs_right[46] ;
 wire \ces_4_2_io_outs_right[47] ;
 wire \ces_4_2_io_outs_right[48] ;
 wire \ces_4_2_io_outs_right[49] ;
 wire \ces_4_2_io_outs_right[4] ;
 wire \ces_4_2_io_outs_right[50] ;
 wire \ces_4_2_io_outs_right[51] ;
 wire \ces_4_2_io_outs_right[52] ;
 wire \ces_4_2_io_outs_right[53] ;
 wire \ces_4_2_io_outs_right[54] ;
 wire \ces_4_2_io_outs_right[55] ;
 wire \ces_4_2_io_outs_right[56] ;
 wire \ces_4_2_io_outs_right[57] ;
 wire \ces_4_2_io_outs_right[58] ;
 wire \ces_4_2_io_outs_right[59] ;
 wire \ces_4_2_io_outs_right[5] ;
 wire \ces_4_2_io_outs_right[60] ;
 wire \ces_4_2_io_outs_right[61] ;
 wire \ces_4_2_io_outs_right[62] ;
 wire \ces_4_2_io_outs_right[63] ;
 wire \ces_4_2_io_outs_right[6] ;
 wire \ces_4_2_io_outs_right[7] ;
 wire \ces_4_2_io_outs_right[8] ;
 wire \ces_4_2_io_outs_right[9] ;
 wire \ces_4_2_io_outs_up[0] ;
 wire \ces_4_2_io_outs_up[10] ;
 wire \ces_4_2_io_outs_up[11] ;
 wire \ces_4_2_io_outs_up[12] ;
 wire \ces_4_2_io_outs_up[13] ;
 wire \ces_4_2_io_outs_up[14] ;
 wire \ces_4_2_io_outs_up[15] ;
 wire \ces_4_2_io_outs_up[16] ;
 wire \ces_4_2_io_outs_up[17] ;
 wire \ces_4_2_io_outs_up[18] ;
 wire \ces_4_2_io_outs_up[19] ;
 wire \ces_4_2_io_outs_up[1] ;
 wire \ces_4_2_io_outs_up[20] ;
 wire \ces_4_2_io_outs_up[21] ;
 wire \ces_4_2_io_outs_up[22] ;
 wire \ces_4_2_io_outs_up[23] ;
 wire \ces_4_2_io_outs_up[24] ;
 wire \ces_4_2_io_outs_up[25] ;
 wire \ces_4_2_io_outs_up[26] ;
 wire \ces_4_2_io_outs_up[27] ;
 wire \ces_4_2_io_outs_up[28] ;
 wire \ces_4_2_io_outs_up[29] ;
 wire \ces_4_2_io_outs_up[2] ;
 wire \ces_4_2_io_outs_up[30] ;
 wire \ces_4_2_io_outs_up[31] ;
 wire \ces_4_2_io_outs_up[32] ;
 wire \ces_4_2_io_outs_up[33] ;
 wire \ces_4_2_io_outs_up[34] ;
 wire \ces_4_2_io_outs_up[35] ;
 wire \ces_4_2_io_outs_up[36] ;
 wire \ces_4_2_io_outs_up[37] ;
 wire \ces_4_2_io_outs_up[38] ;
 wire \ces_4_2_io_outs_up[39] ;
 wire \ces_4_2_io_outs_up[3] ;
 wire \ces_4_2_io_outs_up[40] ;
 wire \ces_4_2_io_outs_up[41] ;
 wire \ces_4_2_io_outs_up[42] ;
 wire \ces_4_2_io_outs_up[43] ;
 wire \ces_4_2_io_outs_up[44] ;
 wire \ces_4_2_io_outs_up[45] ;
 wire \ces_4_2_io_outs_up[46] ;
 wire \ces_4_2_io_outs_up[47] ;
 wire \ces_4_2_io_outs_up[48] ;
 wire \ces_4_2_io_outs_up[49] ;
 wire \ces_4_2_io_outs_up[4] ;
 wire \ces_4_2_io_outs_up[50] ;
 wire \ces_4_2_io_outs_up[51] ;
 wire \ces_4_2_io_outs_up[52] ;
 wire \ces_4_2_io_outs_up[53] ;
 wire \ces_4_2_io_outs_up[54] ;
 wire \ces_4_2_io_outs_up[55] ;
 wire \ces_4_2_io_outs_up[56] ;
 wire \ces_4_2_io_outs_up[57] ;
 wire \ces_4_2_io_outs_up[58] ;
 wire \ces_4_2_io_outs_up[59] ;
 wire \ces_4_2_io_outs_up[5] ;
 wire \ces_4_2_io_outs_up[60] ;
 wire \ces_4_2_io_outs_up[61] ;
 wire \ces_4_2_io_outs_up[62] ;
 wire \ces_4_2_io_outs_up[63] ;
 wire \ces_4_2_io_outs_up[6] ;
 wire \ces_4_2_io_outs_up[7] ;
 wire \ces_4_2_io_outs_up[8] ;
 wire \ces_4_2_io_outs_up[9] ;
 wire \ces_4_3_io_ins_down[0] ;
 wire \ces_4_3_io_ins_down[10] ;
 wire \ces_4_3_io_ins_down[11] ;
 wire \ces_4_3_io_ins_down[12] ;
 wire \ces_4_3_io_ins_down[13] ;
 wire \ces_4_3_io_ins_down[14] ;
 wire \ces_4_3_io_ins_down[15] ;
 wire \ces_4_3_io_ins_down[16] ;
 wire \ces_4_3_io_ins_down[17] ;
 wire \ces_4_3_io_ins_down[18] ;
 wire \ces_4_3_io_ins_down[19] ;
 wire \ces_4_3_io_ins_down[1] ;
 wire \ces_4_3_io_ins_down[20] ;
 wire \ces_4_3_io_ins_down[21] ;
 wire \ces_4_3_io_ins_down[22] ;
 wire \ces_4_3_io_ins_down[23] ;
 wire \ces_4_3_io_ins_down[24] ;
 wire \ces_4_3_io_ins_down[25] ;
 wire \ces_4_3_io_ins_down[26] ;
 wire \ces_4_3_io_ins_down[27] ;
 wire \ces_4_3_io_ins_down[28] ;
 wire \ces_4_3_io_ins_down[29] ;
 wire \ces_4_3_io_ins_down[2] ;
 wire \ces_4_3_io_ins_down[30] ;
 wire \ces_4_3_io_ins_down[31] ;
 wire \ces_4_3_io_ins_down[32] ;
 wire \ces_4_3_io_ins_down[33] ;
 wire \ces_4_3_io_ins_down[34] ;
 wire \ces_4_3_io_ins_down[35] ;
 wire \ces_4_3_io_ins_down[36] ;
 wire \ces_4_3_io_ins_down[37] ;
 wire \ces_4_3_io_ins_down[38] ;
 wire \ces_4_3_io_ins_down[39] ;
 wire \ces_4_3_io_ins_down[3] ;
 wire \ces_4_3_io_ins_down[40] ;
 wire \ces_4_3_io_ins_down[41] ;
 wire \ces_4_3_io_ins_down[42] ;
 wire \ces_4_3_io_ins_down[43] ;
 wire \ces_4_3_io_ins_down[44] ;
 wire \ces_4_3_io_ins_down[45] ;
 wire \ces_4_3_io_ins_down[46] ;
 wire \ces_4_3_io_ins_down[47] ;
 wire \ces_4_3_io_ins_down[48] ;
 wire \ces_4_3_io_ins_down[49] ;
 wire \ces_4_3_io_ins_down[4] ;
 wire \ces_4_3_io_ins_down[50] ;
 wire \ces_4_3_io_ins_down[51] ;
 wire \ces_4_3_io_ins_down[52] ;
 wire \ces_4_3_io_ins_down[53] ;
 wire \ces_4_3_io_ins_down[54] ;
 wire \ces_4_3_io_ins_down[55] ;
 wire \ces_4_3_io_ins_down[56] ;
 wire \ces_4_3_io_ins_down[57] ;
 wire \ces_4_3_io_ins_down[58] ;
 wire \ces_4_3_io_ins_down[59] ;
 wire \ces_4_3_io_ins_down[5] ;
 wire \ces_4_3_io_ins_down[60] ;
 wire \ces_4_3_io_ins_down[61] ;
 wire \ces_4_3_io_ins_down[62] ;
 wire \ces_4_3_io_ins_down[63] ;
 wire \ces_4_3_io_ins_down[6] ;
 wire \ces_4_3_io_ins_down[7] ;
 wire \ces_4_3_io_ins_down[8] ;
 wire \ces_4_3_io_ins_down[9] ;
 wire \ces_4_3_io_ins_left[0] ;
 wire \ces_4_3_io_ins_left[10] ;
 wire \ces_4_3_io_ins_left[11] ;
 wire \ces_4_3_io_ins_left[12] ;
 wire \ces_4_3_io_ins_left[13] ;
 wire \ces_4_3_io_ins_left[14] ;
 wire \ces_4_3_io_ins_left[15] ;
 wire \ces_4_3_io_ins_left[16] ;
 wire \ces_4_3_io_ins_left[17] ;
 wire \ces_4_3_io_ins_left[18] ;
 wire \ces_4_3_io_ins_left[19] ;
 wire \ces_4_3_io_ins_left[1] ;
 wire \ces_4_3_io_ins_left[20] ;
 wire \ces_4_3_io_ins_left[21] ;
 wire \ces_4_3_io_ins_left[22] ;
 wire \ces_4_3_io_ins_left[23] ;
 wire \ces_4_3_io_ins_left[24] ;
 wire \ces_4_3_io_ins_left[25] ;
 wire \ces_4_3_io_ins_left[26] ;
 wire \ces_4_3_io_ins_left[27] ;
 wire \ces_4_3_io_ins_left[28] ;
 wire \ces_4_3_io_ins_left[29] ;
 wire \ces_4_3_io_ins_left[2] ;
 wire \ces_4_3_io_ins_left[30] ;
 wire \ces_4_3_io_ins_left[31] ;
 wire \ces_4_3_io_ins_left[32] ;
 wire \ces_4_3_io_ins_left[33] ;
 wire \ces_4_3_io_ins_left[34] ;
 wire \ces_4_3_io_ins_left[35] ;
 wire \ces_4_3_io_ins_left[36] ;
 wire \ces_4_3_io_ins_left[37] ;
 wire \ces_4_3_io_ins_left[38] ;
 wire \ces_4_3_io_ins_left[39] ;
 wire \ces_4_3_io_ins_left[3] ;
 wire \ces_4_3_io_ins_left[40] ;
 wire \ces_4_3_io_ins_left[41] ;
 wire \ces_4_3_io_ins_left[42] ;
 wire \ces_4_3_io_ins_left[43] ;
 wire \ces_4_3_io_ins_left[44] ;
 wire \ces_4_3_io_ins_left[45] ;
 wire \ces_4_3_io_ins_left[46] ;
 wire \ces_4_3_io_ins_left[47] ;
 wire \ces_4_3_io_ins_left[48] ;
 wire \ces_4_3_io_ins_left[49] ;
 wire \ces_4_3_io_ins_left[4] ;
 wire \ces_4_3_io_ins_left[50] ;
 wire \ces_4_3_io_ins_left[51] ;
 wire \ces_4_3_io_ins_left[52] ;
 wire \ces_4_3_io_ins_left[53] ;
 wire \ces_4_3_io_ins_left[54] ;
 wire \ces_4_3_io_ins_left[55] ;
 wire \ces_4_3_io_ins_left[56] ;
 wire \ces_4_3_io_ins_left[57] ;
 wire \ces_4_3_io_ins_left[58] ;
 wire \ces_4_3_io_ins_left[59] ;
 wire \ces_4_3_io_ins_left[5] ;
 wire \ces_4_3_io_ins_left[60] ;
 wire \ces_4_3_io_ins_left[61] ;
 wire \ces_4_3_io_ins_left[62] ;
 wire \ces_4_3_io_ins_left[63] ;
 wire \ces_4_3_io_ins_left[6] ;
 wire \ces_4_3_io_ins_left[7] ;
 wire \ces_4_3_io_ins_left[8] ;
 wire \ces_4_3_io_ins_left[9] ;
 wire ces_4_3_io_lsbOuts_0;
 wire ces_4_3_io_lsbOuts_1;
 wire ces_4_3_io_lsbOuts_2;
 wire ces_4_3_io_lsbOuts_3;
 wire ces_4_3_io_lsbOuts_4;
 wire ces_4_3_io_lsbOuts_5;
 wire ces_4_3_io_lsbOuts_6;
 wire ces_4_3_io_lsbOuts_7;
 wire \ces_4_3_io_outs_right[0] ;
 wire \ces_4_3_io_outs_right[10] ;
 wire \ces_4_3_io_outs_right[11] ;
 wire \ces_4_3_io_outs_right[12] ;
 wire \ces_4_3_io_outs_right[13] ;
 wire \ces_4_3_io_outs_right[14] ;
 wire \ces_4_3_io_outs_right[15] ;
 wire \ces_4_3_io_outs_right[16] ;
 wire \ces_4_3_io_outs_right[17] ;
 wire \ces_4_3_io_outs_right[18] ;
 wire \ces_4_3_io_outs_right[19] ;
 wire \ces_4_3_io_outs_right[1] ;
 wire \ces_4_3_io_outs_right[20] ;
 wire \ces_4_3_io_outs_right[21] ;
 wire \ces_4_3_io_outs_right[22] ;
 wire \ces_4_3_io_outs_right[23] ;
 wire \ces_4_3_io_outs_right[24] ;
 wire \ces_4_3_io_outs_right[25] ;
 wire \ces_4_3_io_outs_right[26] ;
 wire \ces_4_3_io_outs_right[27] ;
 wire \ces_4_3_io_outs_right[28] ;
 wire \ces_4_3_io_outs_right[29] ;
 wire \ces_4_3_io_outs_right[2] ;
 wire \ces_4_3_io_outs_right[30] ;
 wire \ces_4_3_io_outs_right[31] ;
 wire \ces_4_3_io_outs_right[32] ;
 wire \ces_4_3_io_outs_right[33] ;
 wire \ces_4_3_io_outs_right[34] ;
 wire \ces_4_3_io_outs_right[35] ;
 wire \ces_4_3_io_outs_right[36] ;
 wire \ces_4_3_io_outs_right[37] ;
 wire \ces_4_3_io_outs_right[38] ;
 wire \ces_4_3_io_outs_right[39] ;
 wire \ces_4_3_io_outs_right[3] ;
 wire \ces_4_3_io_outs_right[40] ;
 wire \ces_4_3_io_outs_right[41] ;
 wire \ces_4_3_io_outs_right[42] ;
 wire \ces_4_3_io_outs_right[43] ;
 wire \ces_4_3_io_outs_right[44] ;
 wire \ces_4_3_io_outs_right[45] ;
 wire \ces_4_3_io_outs_right[46] ;
 wire \ces_4_3_io_outs_right[47] ;
 wire \ces_4_3_io_outs_right[48] ;
 wire \ces_4_3_io_outs_right[49] ;
 wire \ces_4_3_io_outs_right[4] ;
 wire \ces_4_3_io_outs_right[50] ;
 wire \ces_4_3_io_outs_right[51] ;
 wire \ces_4_3_io_outs_right[52] ;
 wire \ces_4_3_io_outs_right[53] ;
 wire \ces_4_3_io_outs_right[54] ;
 wire \ces_4_3_io_outs_right[55] ;
 wire \ces_4_3_io_outs_right[56] ;
 wire \ces_4_3_io_outs_right[57] ;
 wire \ces_4_3_io_outs_right[58] ;
 wire \ces_4_3_io_outs_right[59] ;
 wire \ces_4_3_io_outs_right[5] ;
 wire \ces_4_3_io_outs_right[60] ;
 wire \ces_4_3_io_outs_right[61] ;
 wire \ces_4_3_io_outs_right[62] ;
 wire \ces_4_3_io_outs_right[63] ;
 wire \ces_4_3_io_outs_right[6] ;
 wire \ces_4_3_io_outs_right[7] ;
 wire \ces_4_3_io_outs_right[8] ;
 wire \ces_4_3_io_outs_right[9] ;
 wire \ces_4_3_io_outs_up[0] ;
 wire \ces_4_3_io_outs_up[10] ;
 wire \ces_4_3_io_outs_up[11] ;
 wire \ces_4_3_io_outs_up[12] ;
 wire \ces_4_3_io_outs_up[13] ;
 wire \ces_4_3_io_outs_up[14] ;
 wire \ces_4_3_io_outs_up[15] ;
 wire \ces_4_3_io_outs_up[16] ;
 wire \ces_4_3_io_outs_up[17] ;
 wire \ces_4_3_io_outs_up[18] ;
 wire \ces_4_3_io_outs_up[19] ;
 wire \ces_4_3_io_outs_up[1] ;
 wire \ces_4_3_io_outs_up[20] ;
 wire \ces_4_3_io_outs_up[21] ;
 wire \ces_4_3_io_outs_up[22] ;
 wire \ces_4_3_io_outs_up[23] ;
 wire \ces_4_3_io_outs_up[24] ;
 wire \ces_4_3_io_outs_up[25] ;
 wire \ces_4_3_io_outs_up[26] ;
 wire \ces_4_3_io_outs_up[27] ;
 wire \ces_4_3_io_outs_up[28] ;
 wire \ces_4_3_io_outs_up[29] ;
 wire \ces_4_3_io_outs_up[2] ;
 wire \ces_4_3_io_outs_up[30] ;
 wire \ces_4_3_io_outs_up[31] ;
 wire \ces_4_3_io_outs_up[32] ;
 wire \ces_4_3_io_outs_up[33] ;
 wire \ces_4_3_io_outs_up[34] ;
 wire \ces_4_3_io_outs_up[35] ;
 wire \ces_4_3_io_outs_up[36] ;
 wire \ces_4_3_io_outs_up[37] ;
 wire \ces_4_3_io_outs_up[38] ;
 wire \ces_4_3_io_outs_up[39] ;
 wire \ces_4_3_io_outs_up[3] ;
 wire \ces_4_3_io_outs_up[40] ;
 wire \ces_4_3_io_outs_up[41] ;
 wire \ces_4_3_io_outs_up[42] ;
 wire \ces_4_3_io_outs_up[43] ;
 wire \ces_4_3_io_outs_up[44] ;
 wire \ces_4_3_io_outs_up[45] ;
 wire \ces_4_3_io_outs_up[46] ;
 wire \ces_4_3_io_outs_up[47] ;
 wire \ces_4_3_io_outs_up[48] ;
 wire \ces_4_3_io_outs_up[49] ;
 wire \ces_4_3_io_outs_up[4] ;
 wire \ces_4_3_io_outs_up[50] ;
 wire \ces_4_3_io_outs_up[51] ;
 wire \ces_4_3_io_outs_up[52] ;
 wire \ces_4_3_io_outs_up[53] ;
 wire \ces_4_3_io_outs_up[54] ;
 wire \ces_4_3_io_outs_up[55] ;
 wire \ces_4_3_io_outs_up[56] ;
 wire \ces_4_3_io_outs_up[57] ;
 wire \ces_4_3_io_outs_up[58] ;
 wire \ces_4_3_io_outs_up[59] ;
 wire \ces_4_3_io_outs_up[5] ;
 wire \ces_4_3_io_outs_up[60] ;
 wire \ces_4_3_io_outs_up[61] ;
 wire \ces_4_3_io_outs_up[62] ;
 wire \ces_4_3_io_outs_up[63] ;
 wire \ces_4_3_io_outs_up[6] ;
 wire \ces_4_3_io_outs_up[7] ;
 wire \ces_4_3_io_outs_up[8] ;
 wire \ces_4_3_io_outs_up[9] ;
 wire \ces_4_4_io_ins_down[0] ;
 wire \ces_4_4_io_ins_down[10] ;
 wire \ces_4_4_io_ins_down[11] ;
 wire \ces_4_4_io_ins_down[12] ;
 wire \ces_4_4_io_ins_down[13] ;
 wire \ces_4_4_io_ins_down[14] ;
 wire \ces_4_4_io_ins_down[15] ;
 wire \ces_4_4_io_ins_down[16] ;
 wire \ces_4_4_io_ins_down[17] ;
 wire \ces_4_4_io_ins_down[18] ;
 wire \ces_4_4_io_ins_down[19] ;
 wire \ces_4_4_io_ins_down[1] ;
 wire \ces_4_4_io_ins_down[20] ;
 wire \ces_4_4_io_ins_down[21] ;
 wire \ces_4_4_io_ins_down[22] ;
 wire \ces_4_4_io_ins_down[23] ;
 wire \ces_4_4_io_ins_down[24] ;
 wire \ces_4_4_io_ins_down[25] ;
 wire \ces_4_4_io_ins_down[26] ;
 wire \ces_4_4_io_ins_down[27] ;
 wire \ces_4_4_io_ins_down[28] ;
 wire \ces_4_4_io_ins_down[29] ;
 wire \ces_4_4_io_ins_down[2] ;
 wire \ces_4_4_io_ins_down[30] ;
 wire \ces_4_4_io_ins_down[31] ;
 wire \ces_4_4_io_ins_down[32] ;
 wire \ces_4_4_io_ins_down[33] ;
 wire \ces_4_4_io_ins_down[34] ;
 wire \ces_4_4_io_ins_down[35] ;
 wire \ces_4_4_io_ins_down[36] ;
 wire \ces_4_4_io_ins_down[37] ;
 wire \ces_4_4_io_ins_down[38] ;
 wire \ces_4_4_io_ins_down[39] ;
 wire \ces_4_4_io_ins_down[3] ;
 wire \ces_4_4_io_ins_down[40] ;
 wire \ces_4_4_io_ins_down[41] ;
 wire \ces_4_4_io_ins_down[42] ;
 wire \ces_4_4_io_ins_down[43] ;
 wire \ces_4_4_io_ins_down[44] ;
 wire \ces_4_4_io_ins_down[45] ;
 wire \ces_4_4_io_ins_down[46] ;
 wire \ces_4_4_io_ins_down[47] ;
 wire \ces_4_4_io_ins_down[48] ;
 wire \ces_4_4_io_ins_down[49] ;
 wire \ces_4_4_io_ins_down[4] ;
 wire \ces_4_4_io_ins_down[50] ;
 wire \ces_4_4_io_ins_down[51] ;
 wire \ces_4_4_io_ins_down[52] ;
 wire \ces_4_4_io_ins_down[53] ;
 wire \ces_4_4_io_ins_down[54] ;
 wire \ces_4_4_io_ins_down[55] ;
 wire \ces_4_4_io_ins_down[56] ;
 wire \ces_4_4_io_ins_down[57] ;
 wire \ces_4_4_io_ins_down[58] ;
 wire \ces_4_4_io_ins_down[59] ;
 wire \ces_4_4_io_ins_down[5] ;
 wire \ces_4_4_io_ins_down[60] ;
 wire \ces_4_4_io_ins_down[61] ;
 wire \ces_4_4_io_ins_down[62] ;
 wire \ces_4_4_io_ins_down[63] ;
 wire \ces_4_4_io_ins_down[6] ;
 wire \ces_4_4_io_ins_down[7] ;
 wire \ces_4_4_io_ins_down[8] ;
 wire \ces_4_4_io_ins_down[9] ;
 wire \ces_4_4_io_ins_left[0] ;
 wire \ces_4_4_io_ins_left[10] ;
 wire \ces_4_4_io_ins_left[11] ;
 wire \ces_4_4_io_ins_left[12] ;
 wire \ces_4_4_io_ins_left[13] ;
 wire \ces_4_4_io_ins_left[14] ;
 wire \ces_4_4_io_ins_left[15] ;
 wire \ces_4_4_io_ins_left[16] ;
 wire \ces_4_4_io_ins_left[17] ;
 wire \ces_4_4_io_ins_left[18] ;
 wire \ces_4_4_io_ins_left[19] ;
 wire \ces_4_4_io_ins_left[1] ;
 wire \ces_4_4_io_ins_left[20] ;
 wire \ces_4_4_io_ins_left[21] ;
 wire \ces_4_4_io_ins_left[22] ;
 wire \ces_4_4_io_ins_left[23] ;
 wire \ces_4_4_io_ins_left[24] ;
 wire \ces_4_4_io_ins_left[25] ;
 wire \ces_4_4_io_ins_left[26] ;
 wire \ces_4_4_io_ins_left[27] ;
 wire \ces_4_4_io_ins_left[28] ;
 wire \ces_4_4_io_ins_left[29] ;
 wire \ces_4_4_io_ins_left[2] ;
 wire \ces_4_4_io_ins_left[30] ;
 wire \ces_4_4_io_ins_left[31] ;
 wire \ces_4_4_io_ins_left[32] ;
 wire \ces_4_4_io_ins_left[33] ;
 wire \ces_4_4_io_ins_left[34] ;
 wire \ces_4_4_io_ins_left[35] ;
 wire \ces_4_4_io_ins_left[36] ;
 wire \ces_4_4_io_ins_left[37] ;
 wire \ces_4_4_io_ins_left[38] ;
 wire \ces_4_4_io_ins_left[39] ;
 wire \ces_4_4_io_ins_left[3] ;
 wire \ces_4_4_io_ins_left[40] ;
 wire \ces_4_4_io_ins_left[41] ;
 wire \ces_4_4_io_ins_left[42] ;
 wire \ces_4_4_io_ins_left[43] ;
 wire \ces_4_4_io_ins_left[44] ;
 wire \ces_4_4_io_ins_left[45] ;
 wire \ces_4_4_io_ins_left[46] ;
 wire \ces_4_4_io_ins_left[47] ;
 wire \ces_4_4_io_ins_left[48] ;
 wire \ces_4_4_io_ins_left[49] ;
 wire \ces_4_4_io_ins_left[4] ;
 wire \ces_4_4_io_ins_left[50] ;
 wire \ces_4_4_io_ins_left[51] ;
 wire \ces_4_4_io_ins_left[52] ;
 wire \ces_4_4_io_ins_left[53] ;
 wire \ces_4_4_io_ins_left[54] ;
 wire \ces_4_4_io_ins_left[55] ;
 wire \ces_4_4_io_ins_left[56] ;
 wire \ces_4_4_io_ins_left[57] ;
 wire \ces_4_4_io_ins_left[58] ;
 wire \ces_4_4_io_ins_left[59] ;
 wire \ces_4_4_io_ins_left[5] ;
 wire \ces_4_4_io_ins_left[60] ;
 wire \ces_4_4_io_ins_left[61] ;
 wire \ces_4_4_io_ins_left[62] ;
 wire \ces_4_4_io_ins_left[63] ;
 wire \ces_4_4_io_ins_left[6] ;
 wire \ces_4_4_io_ins_left[7] ;
 wire \ces_4_4_io_ins_left[8] ;
 wire \ces_4_4_io_ins_left[9] ;
 wire ces_4_4_io_lsbOuts_0;
 wire ces_4_4_io_lsbOuts_1;
 wire ces_4_4_io_lsbOuts_2;
 wire ces_4_4_io_lsbOuts_3;
 wire ces_4_4_io_lsbOuts_4;
 wire ces_4_4_io_lsbOuts_5;
 wire ces_4_4_io_lsbOuts_6;
 wire ces_4_4_io_lsbOuts_7;
 wire \ces_4_4_io_outs_right[0] ;
 wire \ces_4_4_io_outs_right[10] ;
 wire \ces_4_4_io_outs_right[11] ;
 wire \ces_4_4_io_outs_right[12] ;
 wire \ces_4_4_io_outs_right[13] ;
 wire \ces_4_4_io_outs_right[14] ;
 wire \ces_4_4_io_outs_right[15] ;
 wire \ces_4_4_io_outs_right[16] ;
 wire \ces_4_4_io_outs_right[17] ;
 wire \ces_4_4_io_outs_right[18] ;
 wire \ces_4_4_io_outs_right[19] ;
 wire \ces_4_4_io_outs_right[1] ;
 wire \ces_4_4_io_outs_right[20] ;
 wire \ces_4_4_io_outs_right[21] ;
 wire \ces_4_4_io_outs_right[22] ;
 wire \ces_4_4_io_outs_right[23] ;
 wire \ces_4_4_io_outs_right[24] ;
 wire \ces_4_4_io_outs_right[25] ;
 wire \ces_4_4_io_outs_right[26] ;
 wire \ces_4_4_io_outs_right[27] ;
 wire \ces_4_4_io_outs_right[28] ;
 wire \ces_4_4_io_outs_right[29] ;
 wire \ces_4_4_io_outs_right[2] ;
 wire \ces_4_4_io_outs_right[30] ;
 wire \ces_4_4_io_outs_right[31] ;
 wire \ces_4_4_io_outs_right[32] ;
 wire \ces_4_4_io_outs_right[33] ;
 wire \ces_4_4_io_outs_right[34] ;
 wire \ces_4_4_io_outs_right[35] ;
 wire \ces_4_4_io_outs_right[36] ;
 wire \ces_4_4_io_outs_right[37] ;
 wire \ces_4_4_io_outs_right[38] ;
 wire \ces_4_4_io_outs_right[39] ;
 wire \ces_4_4_io_outs_right[3] ;
 wire \ces_4_4_io_outs_right[40] ;
 wire \ces_4_4_io_outs_right[41] ;
 wire \ces_4_4_io_outs_right[42] ;
 wire \ces_4_4_io_outs_right[43] ;
 wire \ces_4_4_io_outs_right[44] ;
 wire \ces_4_4_io_outs_right[45] ;
 wire \ces_4_4_io_outs_right[46] ;
 wire \ces_4_4_io_outs_right[47] ;
 wire \ces_4_4_io_outs_right[48] ;
 wire \ces_4_4_io_outs_right[49] ;
 wire \ces_4_4_io_outs_right[4] ;
 wire \ces_4_4_io_outs_right[50] ;
 wire \ces_4_4_io_outs_right[51] ;
 wire \ces_4_4_io_outs_right[52] ;
 wire \ces_4_4_io_outs_right[53] ;
 wire \ces_4_4_io_outs_right[54] ;
 wire \ces_4_4_io_outs_right[55] ;
 wire \ces_4_4_io_outs_right[56] ;
 wire \ces_4_4_io_outs_right[57] ;
 wire \ces_4_4_io_outs_right[58] ;
 wire \ces_4_4_io_outs_right[59] ;
 wire \ces_4_4_io_outs_right[5] ;
 wire \ces_4_4_io_outs_right[60] ;
 wire \ces_4_4_io_outs_right[61] ;
 wire \ces_4_4_io_outs_right[62] ;
 wire \ces_4_4_io_outs_right[63] ;
 wire \ces_4_4_io_outs_right[6] ;
 wire \ces_4_4_io_outs_right[7] ;
 wire \ces_4_4_io_outs_right[8] ;
 wire \ces_4_4_io_outs_right[9] ;
 wire \ces_4_4_io_outs_up[0] ;
 wire \ces_4_4_io_outs_up[10] ;
 wire \ces_4_4_io_outs_up[11] ;
 wire \ces_4_4_io_outs_up[12] ;
 wire \ces_4_4_io_outs_up[13] ;
 wire \ces_4_4_io_outs_up[14] ;
 wire \ces_4_4_io_outs_up[15] ;
 wire \ces_4_4_io_outs_up[16] ;
 wire \ces_4_4_io_outs_up[17] ;
 wire \ces_4_4_io_outs_up[18] ;
 wire \ces_4_4_io_outs_up[19] ;
 wire \ces_4_4_io_outs_up[1] ;
 wire \ces_4_4_io_outs_up[20] ;
 wire \ces_4_4_io_outs_up[21] ;
 wire \ces_4_4_io_outs_up[22] ;
 wire \ces_4_4_io_outs_up[23] ;
 wire \ces_4_4_io_outs_up[24] ;
 wire \ces_4_4_io_outs_up[25] ;
 wire \ces_4_4_io_outs_up[26] ;
 wire \ces_4_4_io_outs_up[27] ;
 wire \ces_4_4_io_outs_up[28] ;
 wire \ces_4_4_io_outs_up[29] ;
 wire \ces_4_4_io_outs_up[2] ;
 wire \ces_4_4_io_outs_up[30] ;
 wire \ces_4_4_io_outs_up[31] ;
 wire \ces_4_4_io_outs_up[32] ;
 wire \ces_4_4_io_outs_up[33] ;
 wire \ces_4_4_io_outs_up[34] ;
 wire \ces_4_4_io_outs_up[35] ;
 wire \ces_4_4_io_outs_up[36] ;
 wire \ces_4_4_io_outs_up[37] ;
 wire \ces_4_4_io_outs_up[38] ;
 wire \ces_4_4_io_outs_up[39] ;
 wire \ces_4_4_io_outs_up[3] ;
 wire \ces_4_4_io_outs_up[40] ;
 wire \ces_4_4_io_outs_up[41] ;
 wire \ces_4_4_io_outs_up[42] ;
 wire \ces_4_4_io_outs_up[43] ;
 wire \ces_4_4_io_outs_up[44] ;
 wire \ces_4_4_io_outs_up[45] ;
 wire \ces_4_4_io_outs_up[46] ;
 wire \ces_4_4_io_outs_up[47] ;
 wire \ces_4_4_io_outs_up[48] ;
 wire \ces_4_4_io_outs_up[49] ;
 wire \ces_4_4_io_outs_up[4] ;
 wire \ces_4_4_io_outs_up[50] ;
 wire \ces_4_4_io_outs_up[51] ;
 wire \ces_4_4_io_outs_up[52] ;
 wire \ces_4_4_io_outs_up[53] ;
 wire \ces_4_4_io_outs_up[54] ;
 wire \ces_4_4_io_outs_up[55] ;
 wire \ces_4_4_io_outs_up[56] ;
 wire \ces_4_4_io_outs_up[57] ;
 wire \ces_4_4_io_outs_up[58] ;
 wire \ces_4_4_io_outs_up[59] ;
 wire \ces_4_4_io_outs_up[5] ;
 wire \ces_4_4_io_outs_up[60] ;
 wire \ces_4_4_io_outs_up[61] ;
 wire \ces_4_4_io_outs_up[62] ;
 wire \ces_4_4_io_outs_up[63] ;
 wire \ces_4_4_io_outs_up[6] ;
 wire \ces_4_4_io_outs_up[7] ;
 wire \ces_4_4_io_outs_up[8] ;
 wire \ces_4_4_io_outs_up[9] ;
 wire \ces_4_5_io_ins_down[0] ;
 wire \ces_4_5_io_ins_down[10] ;
 wire \ces_4_5_io_ins_down[11] ;
 wire \ces_4_5_io_ins_down[12] ;
 wire \ces_4_5_io_ins_down[13] ;
 wire \ces_4_5_io_ins_down[14] ;
 wire \ces_4_5_io_ins_down[15] ;
 wire \ces_4_5_io_ins_down[16] ;
 wire \ces_4_5_io_ins_down[17] ;
 wire \ces_4_5_io_ins_down[18] ;
 wire \ces_4_5_io_ins_down[19] ;
 wire \ces_4_5_io_ins_down[1] ;
 wire \ces_4_5_io_ins_down[20] ;
 wire \ces_4_5_io_ins_down[21] ;
 wire \ces_4_5_io_ins_down[22] ;
 wire \ces_4_5_io_ins_down[23] ;
 wire \ces_4_5_io_ins_down[24] ;
 wire \ces_4_5_io_ins_down[25] ;
 wire \ces_4_5_io_ins_down[26] ;
 wire \ces_4_5_io_ins_down[27] ;
 wire \ces_4_5_io_ins_down[28] ;
 wire \ces_4_5_io_ins_down[29] ;
 wire \ces_4_5_io_ins_down[2] ;
 wire \ces_4_5_io_ins_down[30] ;
 wire \ces_4_5_io_ins_down[31] ;
 wire \ces_4_5_io_ins_down[32] ;
 wire \ces_4_5_io_ins_down[33] ;
 wire \ces_4_5_io_ins_down[34] ;
 wire \ces_4_5_io_ins_down[35] ;
 wire \ces_4_5_io_ins_down[36] ;
 wire \ces_4_5_io_ins_down[37] ;
 wire \ces_4_5_io_ins_down[38] ;
 wire \ces_4_5_io_ins_down[39] ;
 wire \ces_4_5_io_ins_down[3] ;
 wire \ces_4_5_io_ins_down[40] ;
 wire \ces_4_5_io_ins_down[41] ;
 wire \ces_4_5_io_ins_down[42] ;
 wire \ces_4_5_io_ins_down[43] ;
 wire \ces_4_5_io_ins_down[44] ;
 wire \ces_4_5_io_ins_down[45] ;
 wire \ces_4_5_io_ins_down[46] ;
 wire \ces_4_5_io_ins_down[47] ;
 wire \ces_4_5_io_ins_down[48] ;
 wire \ces_4_5_io_ins_down[49] ;
 wire \ces_4_5_io_ins_down[4] ;
 wire \ces_4_5_io_ins_down[50] ;
 wire \ces_4_5_io_ins_down[51] ;
 wire \ces_4_5_io_ins_down[52] ;
 wire \ces_4_5_io_ins_down[53] ;
 wire \ces_4_5_io_ins_down[54] ;
 wire \ces_4_5_io_ins_down[55] ;
 wire \ces_4_5_io_ins_down[56] ;
 wire \ces_4_5_io_ins_down[57] ;
 wire \ces_4_5_io_ins_down[58] ;
 wire \ces_4_5_io_ins_down[59] ;
 wire \ces_4_5_io_ins_down[5] ;
 wire \ces_4_5_io_ins_down[60] ;
 wire \ces_4_5_io_ins_down[61] ;
 wire \ces_4_5_io_ins_down[62] ;
 wire \ces_4_5_io_ins_down[63] ;
 wire \ces_4_5_io_ins_down[6] ;
 wire \ces_4_5_io_ins_down[7] ;
 wire \ces_4_5_io_ins_down[8] ;
 wire \ces_4_5_io_ins_down[9] ;
 wire \ces_4_5_io_ins_left[0] ;
 wire \ces_4_5_io_ins_left[10] ;
 wire \ces_4_5_io_ins_left[11] ;
 wire \ces_4_5_io_ins_left[12] ;
 wire \ces_4_5_io_ins_left[13] ;
 wire \ces_4_5_io_ins_left[14] ;
 wire \ces_4_5_io_ins_left[15] ;
 wire \ces_4_5_io_ins_left[16] ;
 wire \ces_4_5_io_ins_left[17] ;
 wire \ces_4_5_io_ins_left[18] ;
 wire \ces_4_5_io_ins_left[19] ;
 wire \ces_4_5_io_ins_left[1] ;
 wire \ces_4_5_io_ins_left[20] ;
 wire \ces_4_5_io_ins_left[21] ;
 wire \ces_4_5_io_ins_left[22] ;
 wire \ces_4_5_io_ins_left[23] ;
 wire \ces_4_5_io_ins_left[24] ;
 wire \ces_4_5_io_ins_left[25] ;
 wire \ces_4_5_io_ins_left[26] ;
 wire \ces_4_5_io_ins_left[27] ;
 wire \ces_4_5_io_ins_left[28] ;
 wire \ces_4_5_io_ins_left[29] ;
 wire \ces_4_5_io_ins_left[2] ;
 wire \ces_4_5_io_ins_left[30] ;
 wire \ces_4_5_io_ins_left[31] ;
 wire \ces_4_5_io_ins_left[32] ;
 wire \ces_4_5_io_ins_left[33] ;
 wire \ces_4_5_io_ins_left[34] ;
 wire \ces_4_5_io_ins_left[35] ;
 wire \ces_4_5_io_ins_left[36] ;
 wire \ces_4_5_io_ins_left[37] ;
 wire \ces_4_5_io_ins_left[38] ;
 wire \ces_4_5_io_ins_left[39] ;
 wire \ces_4_5_io_ins_left[3] ;
 wire \ces_4_5_io_ins_left[40] ;
 wire \ces_4_5_io_ins_left[41] ;
 wire \ces_4_5_io_ins_left[42] ;
 wire \ces_4_5_io_ins_left[43] ;
 wire \ces_4_5_io_ins_left[44] ;
 wire \ces_4_5_io_ins_left[45] ;
 wire \ces_4_5_io_ins_left[46] ;
 wire \ces_4_5_io_ins_left[47] ;
 wire \ces_4_5_io_ins_left[48] ;
 wire \ces_4_5_io_ins_left[49] ;
 wire \ces_4_5_io_ins_left[4] ;
 wire \ces_4_5_io_ins_left[50] ;
 wire \ces_4_5_io_ins_left[51] ;
 wire \ces_4_5_io_ins_left[52] ;
 wire \ces_4_5_io_ins_left[53] ;
 wire \ces_4_5_io_ins_left[54] ;
 wire \ces_4_5_io_ins_left[55] ;
 wire \ces_4_5_io_ins_left[56] ;
 wire \ces_4_5_io_ins_left[57] ;
 wire \ces_4_5_io_ins_left[58] ;
 wire \ces_4_5_io_ins_left[59] ;
 wire \ces_4_5_io_ins_left[5] ;
 wire \ces_4_5_io_ins_left[60] ;
 wire \ces_4_5_io_ins_left[61] ;
 wire \ces_4_5_io_ins_left[62] ;
 wire \ces_4_5_io_ins_left[63] ;
 wire \ces_4_5_io_ins_left[6] ;
 wire \ces_4_5_io_ins_left[7] ;
 wire \ces_4_5_io_ins_left[8] ;
 wire \ces_4_5_io_ins_left[9] ;
 wire ces_4_5_io_lsbOuts_0;
 wire ces_4_5_io_lsbOuts_1;
 wire ces_4_5_io_lsbOuts_2;
 wire ces_4_5_io_lsbOuts_3;
 wire ces_4_5_io_lsbOuts_4;
 wire ces_4_5_io_lsbOuts_5;
 wire ces_4_5_io_lsbOuts_6;
 wire ces_4_5_io_lsbOuts_7;
 wire \ces_4_5_io_outs_right[0] ;
 wire \ces_4_5_io_outs_right[10] ;
 wire \ces_4_5_io_outs_right[11] ;
 wire \ces_4_5_io_outs_right[12] ;
 wire \ces_4_5_io_outs_right[13] ;
 wire \ces_4_5_io_outs_right[14] ;
 wire \ces_4_5_io_outs_right[15] ;
 wire \ces_4_5_io_outs_right[16] ;
 wire \ces_4_5_io_outs_right[17] ;
 wire \ces_4_5_io_outs_right[18] ;
 wire \ces_4_5_io_outs_right[19] ;
 wire \ces_4_5_io_outs_right[1] ;
 wire \ces_4_5_io_outs_right[20] ;
 wire \ces_4_5_io_outs_right[21] ;
 wire \ces_4_5_io_outs_right[22] ;
 wire \ces_4_5_io_outs_right[23] ;
 wire \ces_4_5_io_outs_right[24] ;
 wire \ces_4_5_io_outs_right[25] ;
 wire \ces_4_5_io_outs_right[26] ;
 wire \ces_4_5_io_outs_right[27] ;
 wire \ces_4_5_io_outs_right[28] ;
 wire \ces_4_5_io_outs_right[29] ;
 wire \ces_4_5_io_outs_right[2] ;
 wire \ces_4_5_io_outs_right[30] ;
 wire \ces_4_5_io_outs_right[31] ;
 wire \ces_4_5_io_outs_right[32] ;
 wire \ces_4_5_io_outs_right[33] ;
 wire \ces_4_5_io_outs_right[34] ;
 wire \ces_4_5_io_outs_right[35] ;
 wire \ces_4_5_io_outs_right[36] ;
 wire \ces_4_5_io_outs_right[37] ;
 wire \ces_4_5_io_outs_right[38] ;
 wire \ces_4_5_io_outs_right[39] ;
 wire \ces_4_5_io_outs_right[3] ;
 wire \ces_4_5_io_outs_right[40] ;
 wire \ces_4_5_io_outs_right[41] ;
 wire \ces_4_5_io_outs_right[42] ;
 wire \ces_4_5_io_outs_right[43] ;
 wire \ces_4_5_io_outs_right[44] ;
 wire \ces_4_5_io_outs_right[45] ;
 wire \ces_4_5_io_outs_right[46] ;
 wire \ces_4_5_io_outs_right[47] ;
 wire \ces_4_5_io_outs_right[48] ;
 wire \ces_4_5_io_outs_right[49] ;
 wire \ces_4_5_io_outs_right[4] ;
 wire \ces_4_5_io_outs_right[50] ;
 wire \ces_4_5_io_outs_right[51] ;
 wire \ces_4_5_io_outs_right[52] ;
 wire \ces_4_5_io_outs_right[53] ;
 wire \ces_4_5_io_outs_right[54] ;
 wire \ces_4_5_io_outs_right[55] ;
 wire \ces_4_5_io_outs_right[56] ;
 wire \ces_4_5_io_outs_right[57] ;
 wire \ces_4_5_io_outs_right[58] ;
 wire \ces_4_5_io_outs_right[59] ;
 wire \ces_4_5_io_outs_right[5] ;
 wire \ces_4_5_io_outs_right[60] ;
 wire \ces_4_5_io_outs_right[61] ;
 wire \ces_4_5_io_outs_right[62] ;
 wire \ces_4_5_io_outs_right[63] ;
 wire \ces_4_5_io_outs_right[6] ;
 wire \ces_4_5_io_outs_right[7] ;
 wire \ces_4_5_io_outs_right[8] ;
 wire \ces_4_5_io_outs_right[9] ;
 wire \ces_4_5_io_outs_up[0] ;
 wire \ces_4_5_io_outs_up[10] ;
 wire \ces_4_5_io_outs_up[11] ;
 wire \ces_4_5_io_outs_up[12] ;
 wire \ces_4_5_io_outs_up[13] ;
 wire \ces_4_5_io_outs_up[14] ;
 wire \ces_4_5_io_outs_up[15] ;
 wire \ces_4_5_io_outs_up[16] ;
 wire \ces_4_5_io_outs_up[17] ;
 wire \ces_4_5_io_outs_up[18] ;
 wire \ces_4_5_io_outs_up[19] ;
 wire \ces_4_5_io_outs_up[1] ;
 wire \ces_4_5_io_outs_up[20] ;
 wire \ces_4_5_io_outs_up[21] ;
 wire \ces_4_5_io_outs_up[22] ;
 wire \ces_4_5_io_outs_up[23] ;
 wire \ces_4_5_io_outs_up[24] ;
 wire \ces_4_5_io_outs_up[25] ;
 wire \ces_4_5_io_outs_up[26] ;
 wire \ces_4_5_io_outs_up[27] ;
 wire \ces_4_5_io_outs_up[28] ;
 wire \ces_4_5_io_outs_up[29] ;
 wire \ces_4_5_io_outs_up[2] ;
 wire \ces_4_5_io_outs_up[30] ;
 wire \ces_4_5_io_outs_up[31] ;
 wire \ces_4_5_io_outs_up[32] ;
 wire \ces_4_5_io_outs_up[33] ;
 wire \ces_4_5_io_outs_up[34] ;
 wire \ces_4_5_io_outs_up[35] ;
 wire \ces_4_5_io_outs_up[36] ;
 wire \ces_4_5_io_outs_up[37] ;
 wire \ces_4_5_io_outs_up[38] ;
 wire \ces_4_5_io_outs_up[39] ;
 wire \ces_4_5_io_outs_up[3] ;
 wire \ces_4_5_io_outs_up[40] ;
 wire \ces_4_5_io_outs_up[41] ;
 wire \ces_4_5_io_outs_up[42] ;
 wire \ces_4_5_io_outs_up[43] ;
 wire \ces_4_5_io_outs_up[44] ;
 wire \ces_4_5_io_outs_up[45] ;
 wire \ces_4_5_io_outs_up[46] ;
 wire \ces_4_5_io_outs_up[47] ;
 wire \ces_4_5_io_outs_up[48] ;
 wire \ces_4_5_io_outs_up[49] ;
 wire \ces_4_5_io_outs_up[4] ;
 wire \ces_4_5_io_outs_up[50] ;
 wire \ces_4_5_io_outs_up[51] ;
 wire \ces_4_5_io_outs_up[52] ;
 wire \ces_4_5_io_outs_up[53] ;
 wire \ces_4_5_io_outs_up[54] ;
 wire \ces_4_5_io_outs_up[55] ;
 wire \ces_4_5_io_outs_up[56] ;
 wire \ces_4_5_io_outs_up[57] ;
 wire \ces_4_5_io_outs_up[58] ;
 wire \ces_4_5_io_outs_up[59] ;
 wire \ces_4_5_io_outs_up[5] ;
 wire \ces_4_5_io_outs_up[60] ;
 wire \ces_4_5_io_outs_up[61] ;
 wire \ces_4_5_io_outs_up[62] ;
 wire \ces_4_5_io_outs_up[63] ;
 wire \ces_4_5_io_outs_up[6] ;
 wire \ces_4_5_io_outs_up[7] ;
 wire \ces_4_5_io_outs_up[8] ;
 wire \ces_4_5_io_outs_up[9] ;
 wire \ces_4_6_io_ins_down[0] ;
 wire \ces_4_6_io_ins_down[10] ;
 wire \ces_4_6_io_ins_down[11] ;
 wire \ces_4_6_io_ins_down[12] ;
 wire \ces_4_6_io_ins_down[13] ;
 wire \ces_4_6_io_ins_down[14] ;
 wire \ces_4_6_io_ins_down[15] ;
 wire \ces_4_6_io_ins_down[16] ;
 wire \ces_4_6_io_ins_down[17] ;
 wire \ces_4_6_io_ins_down[18] ;
 wire \ces_4_6_io_ins_down[19] ;
 wire \ces_4_6_io_ins_down[1] ;
 wire \ces_4_6_io_ins_down[20] ;
 wire \ces_4_6_io_ins_down[21] ;
 wire \ces_4_6_io_ins_down[22] ;
 wire \ces_4_6_io_ins_down[23] ;
 wire \ces_4_6_io_ins_down[24] ;
 wire \ces_4_6_io_ins_down[25] ;
 wire \ces_4_6_io_ins_down[26] ;
 wire \ces_4_6_io_ins_down[27] ;
 wire \ces_4_6_io_ins_down[28] ;
 wire \ces_4_6_io_ins_down[29] ;
 wire \ces_4_6_io_ins_down[2] ;
 wire \ces_4_6_io_ins_down[30] ;
 wire \ces_4_6_io_ins_down[31] ;
 wire \ces_4_6_io_ins_down[32] ;
 wire \ces_4_6_io_ins_down[33] ;
 wire \ces_4_6_io_ins_down[34] ;
 wire \ces_4_6_io_ins_down[35] ;
 wire \ces_4_6_io_ins_down[36] ;
 wire \ces_4_6_io_ins_down[37] ;
 wire \ces_4_6_io_ins_down[38] ;
 wire \ces_4_6_io_ins_down[39] ;
 wire \ces_4_6_io_ins_down[3] ;
 wire \ces_4_6_io_ins_down[40] ;
 wire \ces_4_6_io_ins_down[41] ;
 wire \ces_4_6_io_ins_down[42] ;
 wire \ces_4_6_io_ins_down[43] ;
 wire \ces_4_6_io_ins_down[44] ;
 wire \ces_4_6_io_ins_down[45] ;
 wire \ces_4_6_io_ins_down[46] ;
 wire \ces_4_6_io_ins_down[47] ;
 wire \ces_4_6_io_ins_down[48] ;
 wire \ces_4_6_io_ins_down[49] ;
 wire \ces_4_6_io_ins_down[4] ;
 wire \ces_4_6_io_ins_down[50] ;
 wire \ces_4_6_io_ins_down[51] ;
 wire \ces_4_6_io_ins_down[52] ;
 wire \ces_4_6_io_ins_down[53] ;
 wire \ces_4_6_io_ins_down[54] ;
 wire \ces_4_6_io_ins_down[55] ;
 wire \ces_4_6_io_ins_down[56] ;
 wire \ces_4_6_io_ins_down[57] ;
 wire \ces_4_6_io_ins_down[58] ;
 wire \ces_4_6_io_ins_down[59] ;
 wire \ces_4_6_io_ins_down[5] ;
 wire \ces_4_6_io_ins_down[60] ;
 wire \ces_4_6_io_ins_down[61] ;
 wire \ces_4_6_io_ins_down[62] ;
 wire \ces_4_6_io_ins_down[63] ;
 wire \ces_4_6_io_ins_down[6] ;
 wire \ces_4_6_io_ins_down[7] ;
 wire \ces_4_6_io_ins_down[8] ;
 wire \ces_4_6_io_ins_down[9] ;
 wire \ces_4_6_io_ins_left[0] ;
 wire \ces_4_6_io_ins_left[10] ;
 wire \ces_4_6_io_ins_left[11] ;
 wire \ces_4_6_io_ins_left[12] ;
 wire \ces_4_6_io_ins_left[13] ;
 wire \ces_4_6_io_ins_left[14] ;
 wire \ces_4_6_io_ins_left[15] ;
 wire \ces_4_6_io_ins_left[16] ;
 wire \ces_4_6_io_ins_left[17] ;
 wire \ces_4_6_io_ins_left[18] ;
 wire \ces_4_6_io_ins_left[19] ;
 wire \ces_4_6_io_ins_left[1] ;
 wire \ces_4_6_io_ins_left[20] ;
 wire \ces_4_6_io_ins_left[21] ;
 wire \ces_4_6_io_ins_left[22] ;
 wire \ces_4_6_io_ins_left[23] ;
 wire \ces_4_6_io_ins_left[24] ;
 wire \ces_4_6_io_ins_left[25] ;
 wire \ces_4_6_io_ins_left[26] ;
 wire \ces_4_6_io_ins_left[27] ;
 wire \ces_4_6_io_ins_left[28] ;
 wire \ces_4_6_io_ins_left[29] ;
 wire \ces_4_6_io_ins_left[2] ;
 wire \ces_4_6_io_ins_left[30] ;
 wire \ces_4_6_io_ins_left[31] ;
 wire \ces_4_6_io_ins_left[32] ;
 wire \ces_4_6_io_ins_left[33] ;
 wire \ces_4_6_io_ins_left[34] ;
 wire \ces_4_6_io_ins_left[35] ;
 wire \ces_4_6_io_ins_left[36] ;
 wire \ces_4_6_io_ins_left[37] ;
 wire \ces_4_6_io_ins_left[38] ;
 wire \ces_4_6_io_ins_left[39] ;
 wire \ces_4_6_io_ins_left[3] ;
 wire \ces_4_6_io_ins_left[40] ;
 wire \ces_4_6_io_ins_left[41] ;
 wire \ces_4_6_io_ins_left[42] ;
 wire \ces_4_6_io_ins_left[43] ;
 wire \ces_4_6_io_ins_left[44] ;
 wire \ces_4_6_io_ins_left[45] ;
 wire \ces_4_6_io_ins_left[46] ;
 wire \ces_4_6_io_ins_left[47] ;
 wire \ces_4_6_io_ins_left[48] ;
 wire \ces_4_6_io_ins_left[49] ;
 wire \ces_4_6_io_ins_left[4] ;
 wire \ces_4_6_io_ins_left[50] ;
 wire \ces_4_6_io_ins_left[51] ;
 wire \ces_4_6_io_ins_left[52] ;
 wire \ces_4_6_io_ins_left[53] ;
 wire \ces_4_6_io_ins_left[54] ;
 wire \ces_4_6_io_ins_left[55] ;
 wire \ces_4_6_io_ins_left[56] ;
 wire \ces_4_6_io_ins_left[57] ;
 wire \ces_4_6_io_ins_left[58] ;
 wire \ces_4_6_io_ins_left[59] ;
 wire \ces_4_6_io_ins_left[5] ;
 wire \ces_4_6_io_ins_left[60] ;
 wire \ces_4_6_io_ins_left[61] ;
 wire \ces_4_6_io_ins_left[62] ;
 wire \ces_4_6_io_ins_left[63] ;
 wire \ces_4_6_io_ins_left[6] ;
 wire \ces_4_6_io_ins_left[7] ;
 wire \ces_4_6_io_ins_left[8] ;
 wire \ces_4_6_io_ins_left[9] ;
 wire ces_4_6_io_lsbOuts_0;
 wire ces_4_6_io_lsbOuts_1;
 wire ces_4_6_io_lsbOuts_2;
 wire ces_4_6_io_lsbOuts_3;
 wire ces_4_6_io_lsbOuts_4;
 wire ces_4_6_io_lsbOuts_5;
 wire ces_4_6_io_lsbOuts_6;
 wire ces_4_6_io_lsbOuts_7;
 wire \ces_4_6_io_outs_right[0] ;
 wire \ces_4_6_io_outs_right[10] ;
 wire \ces_4_6_io_outs_right[11] ;
 wire \ces_4_6_io_outs_right[12] ;
 wire \ces_4_6_io_outs_right[13] ;
 wire \ces_4_6_io_outs_right[14] ;
 wire \ces_4_6_io_outs_right[15] ;
 wire \ces_4_6_io_outs_right[16] ;
 wire \ces_4_6_io_outs_right[17] ;
 wire \ces_4_6_io_outs_right[18] ;
 wire \ces_4_6_io_outs_right[19] ;
 wire \ces_4_6_io_outs_right[1] ;
 wire \ces_4_6_io_outs_right[20] ;
 wire \ces_4_6_io_outs_right[21] ;
 wire \ces_4_6_io_outs_right[22] ;
 wire \ces_4_6_io_outs_right[23] ;
 wire \ces_4_6_io_outs_right[24] ;
 wire \ces_4_6_io_outs_right[25] ;
 wire \ces_4_6_io_outs_right[26] ;
 wire \ces_4_6_io_outs_right[27] ;
 wire \ces_4_6_io_outs_right[28] ;
 wire \ces_4_6_io_outs_right[29] ;
 wire \ces_4_6_io_outs_right[2] ;
 wire \ces_4_6_io_outs_right[30] ;
 wire \ces_4_6_io_outs_right[31] ;
 wire \ces_4_6_io_outs_right[32] ;
 wire \ces_4_6_io_outs_right[33] ;
 wire \ces_4_6_io_outs_right[34] ;
 wire \ces_4_6_io_outs_right[35] ;
 wire \ces_4_6_io_outs_right[36] ;
 wire \ces_4_6_io_outs_right[37] ;
 wire \ces_4_6_io_outs_right[38] ;
 wire \ces_4_6_io_outs_right[39] ;
 wire \ces_4_6_io_outs_right[3] ;
 wire \ces_4_6_io_outs_right[40] ;
 wire \ces_4_6_io_outs_right[41] ;
 wire \ces_4_6_io_outs_right[42] ;
 wire \ces_4_6_io_outs_right[43] ;
 wire \ces_4_6_io_outs_right[44] ;
 wire \ces_4_6_io_outs_right[45] ;
 wire \ces_4_6_io_outs_right[46] ;
 wire \ces_4_6_io_outs_right[47] ;
 wire \ces_4_6_io_outs_right[48] ;
 wire \ces_4_6_io_outs_right[49] ;
 wire \ces_4_6_io_outs_right[4] ;
 wire \ces_4_6_io_outs_right[50] ;
 wire \ces_4_6_io_outs_right[51] ;
 wire \ces_4_6_io_outs_right[52] ;
 wire \ces_4_6_io_outs_right[53] ;
 wire \ces_4_6_io_outs_right[54] ;
 wire \ces_4_6_io_outs_right[55] ;
 wire \ces_4_6_io_outs_right[56] ;
 wire \ces_4_6_io_outs_right[57] ;
 wire \ces_4_6_io_outs_right[58] ;
 wire \ces_4_6_io_outs_right[59] ;
 wire \ces_4_6_io_outs_right[5] ;
 wire \ces_4_6_io_outs_right[60] ;
 wire \ces_4_6_io_outs_right[61] ;
 wire \ces_4_6_io_outs_right[62] ;
 wire \ces_4_6_io_outs_right[63] ;
 wire \ces_4_6_io_outs_right[6] ;
 wire \ces_4_6_io_outs_right[7] ;
 wire \ces_4_6_io_outs_right[8] ;
 wire \ces_4_6_io_outs_right[9] ;
 wire \ces_4_6_io_outs_up[0] ;
 wire \ces_4_6_io_outs_up[10] ;
 wire \ces_4_6_io_outs_up[11] ;
 wire \ces_4_6_io_outs_up[12] ;
 wire \ces_4_6_io_outs_up[13] ;
 wire \ces_4_6_io_outs_up[14] ;
 wire \ces_4_6_io_outs_up[15] ;
 wire \ces_4_6_io_outs_up[16] ;
 wire \ces_4_6_io_outs_up[17] ;
 wire \ces_4_6_io_outs_up[18] ;
 wire \ces_4_6_io_outs_up[19] ;
 wire \ces_4_6_io_outs_up[1] ;
 wire \ces_4_6_io_outs_up[20] ;
 wire \ces_4_6_io_outs_up[21] ;
 wire \ces_4_6_io_outs_up[22] ;
 wire \ces_4_6_io_outs_up[23] ;
 wire \ces_4_6_io_outs_up[24] ;
 wire \ces_4_6_io_outs_up[25] ;
 wire \ces_4_6_io_outs_up[26] ;
 wire \ces_4_6_io_outs_up[27] ;
 wire \ces_4_6_io_outs_up[28] ;
 wire \ces_4_6_io_outs_up[29] ;
 wire \ces_4_6_io_outs_up[2] ;
 wire \ces_4_6_io_outs_up[30] ;
 wire \ces_4_6_io_outs_up[31] ;
 wire \ces_4_6_io_outs_up[32] ;
 wire \ces_4_6_io_outs_up[33] ;
 wire \ces_4_6_io_outs_up[34] ;
 wire \ces_4_6_io_outs_up[35] ;
 wire \ces_4_6_io_outs_up[36] ;
 wire \ces_4_6_io_outs_up[37] ;
 wire \ces_4_6_io_outs_up[38] ;
 wire \ces_4_6_io_outs_up[39] ;
 wire \ces_4_6_io_outs_up[3] ;
 wire \ces_4_6_io_outs_up[40] ;
 wire \ces_4_6_io_outs_up[41] ;
 wire \ces_4_6_io_outs_up[42] ;
 wire \ces_4_6_io_outs_up[43] ;
 wire \ces_4_6_io_outs_up[44] ;
 wire \ces_4_6_io_outs_up[45] ;
 wire \ces_4_6_io_outs_up[46] ;
 wire \ces_4_6_io_outs_up[47] ;
 wire \ces_4_6_io_outs_up[48] ;
 wire \ces_4_6_io_outs_up[49] ;
 wire \ces_4_6_io_outs_up[4] ;
 wire \ces_4_6_io_outs_up[50] ;
 wire \ces_4_6_io_outs_up[51] ;
 wire \ces_4_6_io_outs_up[52] ;
 wire \ces_4_6_io_outs_up[53] ;
 wire \ces_4_6_io_outs_up[54] ;
 wire \ces_4_6_io_outs_up[55] ;
 wire \ces_4_6_io_outs_up[56] ;
 wire \ces_4_6_io_outs_up[57] ;
 wire \ces_4_6_io_outs_up[58] ;
 wire \ces_4_6_io_outs_up[59] ;
 wire \ces_4_6_io_outs_up[5] ;
 wire \ces_4_6_io_outs_up[60] ;
 wire \ces_4_6_io_outs_up[61] ;
 wire \ces_4_6_io_outs_up[62] ;
 wire \ces_4_6_io_outs_up[63] ;
 wire \ces_4_6_io_outs_up[6] ;
 wire \ces_4_6_io_outs_up[7] ;
 wire \ces_4_6_io_outs_up[8] ;
 wire \ces_4_6_io_outs_up[9] ;
 wire \ces_4_7_io_ins_down[0] ;
 wire \ces_4_7_io_ins_down[10] ;
 wire \ces_4_7_io_ins_down[11] ;
 wire \ces_4_7_io_ins_down[12] ;
 wire \ces_4_7_io_ins_down[13] ;
 wire \ces_4_7_io_ins_down[14] ;
 wire \ces_4_7_io_ins_down[15] ;
 wire \ces_4_7_io_ins_down[16] ;
 wire \ces_4_7_io_ins_down[17] ;
 wire \ces_4_7_io_ins_down[18] ;
 wire \ces_4_7_io_ins_down[19] ;
 wire \ces_4_7_io_ins_down[1] ;
 wire \ces_4_7_io_ins_down[20] ;
 wire \ces_4_7_io_ins_down[21] ;
 wire \ces_4_7_io_ins_down[22] ;
 wire \ces_4_7_io_ins_down[23] ;
 wire \ces_4_7_io_ins_down[24] ;
 wire \ces_4_7_io_ins_down[25] ;
 wire \ces_4_7_io_ins_down[26] ;
 wire \ces_4_7_io_ins_down[27] ;
 wire \ces_4_7_io_ins_down[28] ;
 wire \ces_4_7_io_ins_down[29] ;
 wire \ces_4_7_io_ins_down[2] ;
 wire \ces_4_7_io_ins_down[30] ;
 wire \ces_4_7_io_ins_down[31] ;
 wire \ces_4_7_io_ins_down[32] ;
 wire \ces_4_7_io_ins_down[33] ;
 wire \ces_4_7_io_ins_down[34] ;
 wire \ces_4_7_io_ins_down[35] ;
 wire \ces_4_7_io_ins_down[36] ;
 wire \ces_4_7_io_ins_down[37] ;
 wire \ces_4_7_io_ins_down[38] ;
 wire \ces_4_7_io_ins_down[39] ;
 wire \ces_4_7_io_ins_down[3] ;
 wire \ces_4_7_io_ins_down[40] ;
 wire \ces_4_7_io_ins_down[41] ;
 wire \ces_4_7_io_ins_down[42] ;
 wire \ces_4_7_io_ins_down[43] ;
 wire \ces_4_7_io_ins_down[44] ;
 wire \ces_4_7_io_ins_down[45] ;
 wire \ces_4_7_io_ins_down[46] ;
 wire \ces_4_7_io_ins_down[47] ;
 wire \ces_4_7_io_ins_down[48] ;
 wire \ces_4_7_io_ins_down[49] ;
 wire \ces_4_7_io_ins_down[4] ;
 wire \ces_4_7_io_ins_down[50] ;
 wire \ces_4_7_io_ins_down[51] ;
 wire \ces_4_7_io_ins_down[52] ;
 wire \ces_4_7_io_ins_down[53] ;
 wire \ces_4_7_io_ins_down[54] ;
 wire \ces_4_7_io_ins_down[55] ;
 wire \ces_4_7_io_ins_down[56] ;
 wire \ces_4_7_io_ins_down[57] ;
 wire \ces_4_7_io_ins_down[58] ;
 wire \ces_4_7_io_ins_down[59] ;
 wire \ces_4_7_io_ins_down[5] ;
 wire \ces_4_7_io_ins_down[60] ;
 wire \ces_4_7_io_ins_down[61] ;
 wire \ces_4_7_io_ins_down[62] ;
 wire \ces_4_7_io_ins_down[63] ;
 wire \ces_4_7_io_ins_down[6] ;
 wire \ces_4_7_io_ins_down[7] ;
 wire \ces_4_7_io_ins_down[8] ;
 wire \ces_4_7_io_ins_down[9] ;
 wire ces_4_7_io_lsbOuts_0;
 wire ces_4_7_io_lsbOuts_1;
 wire ces_4_7_io_lsbOuts_2;
 wire ces_4_7_io_lsbOuts_3;
 wire ces_4_7_io_lsbOuts_4;
 wire ces_4_7_io_lsbOuts_5;
 wire ces_4_7_io_lsbOuts_6;
 wire ces_4_7_io_lsbOuts_7;
 wire \ces_4_7_io_outs_up[0] ;
 wire \ces_4_7_io_outs_up[10] ;
 wire \ces_4_7_io_outs_up[11] ;
 wire \ces_4_7_io_outs_up[12] ;
 wire \ces_4_7_io_outs_up[13] ;
 wire \ces_4_7_io_outs_up[14] ;
 wire \ces_4_7_io_outs_up[15] ;
 wire \ces_4_7_io_outs_up[16] ;
 wire \ces_4_7_io_outs_up[17] ;
 wire \ces_4_7_io_outs_up[18] ;
 wire \ces_4_7_io_outs_up[19] ;
 wire \ces_4_7_io_outs_up[1] ;
 wire \ces_4_7_io_outs_up[20] ;
 wire \ces_4_7_io_outs_up[21] ;
 wire \ces_4_7_io_outs_up[22] ;
 wire \ces_4_7_io_outs_up[23] ;
 wire \ces_4_7_io_outs_up[24] ;
 wire \ces_4_7_io_outs_up[25] ;
 wire \ces_4_7_io_outs_up[26] ;
 wire \ces_4_7_io_outs_up[27] ;
 wire \ces_4_7_io_outs_up[28] ;
 wire \ces_4_7_io_outs_up[29] ;
 wire \ces_4_7_io_outs_up[2] ;
 wire \ces_4_7_io_outs_up[30] ;
 wire \ces_4_7_io_outs_up[31] ;
 wire \ces_4_7_io_outs_up[32] ;
 wire \ces_4_7_io_outs_up[33] ;
 wire \ces_4_7_io_outs_up[34] ;
 wire \ces_4_7_io_outs_up[35] ;
 wire \ces_4_7_io_outs_up[36] ;
 wire \ces_4_7_io_outs_up[37] ;
 wire \ces_4_7_io_outs_up[38] ;
 wire \ces_4_7_io_outs_up[39] ;
 wire \ces_4_7_io_outs_up[3] ;
 wire \ces_4_7_io_outs_up[40] ;
 wire \ces_4_7_io_outs_up[41] ;
 wire \ces_4_7_io_outs_up[42] ;
 wire \ces_4_7_io_outs_up[43] ;
 wire \ces_4_7_io_outs_up[44] ;
 wire \ces_4_7_io_outs_up[45] ;
 wire \ces_4_7_io_outs_up[46] ;
 wire \ces_4_7_io_outs_up[47] ;
 wire \ces_4_7_io_outs_up[48] ;
 wire \ces_4_7_io_outs_up[49] ;
 wire \ces_4_7_io_outs_up[4] ;
 wire \ces_4_7_io_outs_up[50] ;
 wire \ces_4_7_io_outs_up[51] ;
 wire \ces_4_7_io_outs_up[52] ;
 wire \ces_4_7_io_outs_up[53] ;
 wire \ces_4_7_io_outs_up[54] ;
 wire \ces_4_7_io_outs_up[55] ;
 wire \ces_4_7_io_outs_up[56] ;
 wire \ces_4_7_io_outs_up[57] ;
 wire \ces_4_7_io_outs_up[58] ;
 wire \ces_4_7_io_outs_up[59] ;
 wire \ces_4_7_io_outs_up[5] ;
 wire \ces_4_7_io_outs_up[60] ;
 wire \ces_4_7_io_outs_up[61] ;
 wire \ces_4_7_io_outs_up[62] ;
 wire \ces_4_7_io_outs_up[63] ;
 wire \ces_4_7_io_outs_up[6] ;
 wire \ces_4_7_io_outs_up[7] ;
 wire \ces_4_7_io_outs_up[8] ;
 wire \ces_4_7_io_outs_up[9] ;
 wire \ces_5_0_io_ins_down[0] ;
 wire \ces_5_0_io_ins_down[10] ;
 wire \ces_5_0_io_ins_down[11] ;
 wire \ces_5_0_io_ins_down[12] ;
 wire \ces_5_0_io_ins_down[13] ;
 wire \ces_5_0_io_ins_down[14] ;
 wire \ces_5_0_io_ins_down[15] ;
 wire \ces_5_0_io_ins_down[16] ;
 wire \ces_5_0_io_ins_down[17] ;
 wire \ces_5_0_io_ins_down[18] ;
 wire \ces_5_0_io_ins_down[19] ;
 wire \ces_5_0_io_ins_down[1] ;
 wire \ces_5_0_io_ins_down[20] ;
 wire \ces_5_0_io_ins_down[21] ;
 wire \ces_5_0_io_ins_down[22] ;
 wire \ces_5_0_io_ins_down[23] ;
 wire \ces_5_0_io_ins_down[24] ;
 wire \ces_5_0_io_ins_down[25] ;
 wire \ces_5_0_io_ins_down[26] ;
 wire \ces_5_0_io_ins_down[27] ;
 wire \ces_5_0_io_ins_down[28] ;
 wire \ces_5_0_io_ins_down[29] ;
 wire \ces_5_0_io_ins_down[2] ;
 wire \ces_5_0_io_ins_down[30] ;
 wire \ces_5_0_io_ins_down[31] ;
 wire \ces_5_0_io_ins_down[32] ;
 wire \ces_5_0_io_ins_down[33] ;
 wire \ces_5_0_io_ins_down[34] ;
 wire \ces_5_0_io_ins_down[35] ;
 wire \ces_5_0_io_ins_down[36] ;
 wire \ces_5_0_io_ins_down[37] ;
 wire \ces_5_0_io_ins_down[38] ;
 wire \ces_5_0_io_ins_down[39] ;
 wire \ces_5_0_io_ins_down[3] ;
 wire \ces_5_0_io_ins_down[40] ;
 wire \ces_5_0_io_ins_down[41] ;
 wire \ces_5_0_io_ins_down[42] ;
 wire \ces_5_0_io_ins_down[43] ;
 wire \ces_5_0_io_ins_down[44] ;
 wire \ces_5_0_io_ins_down[45] ;
 wire \ces_5_0_io_ins_down[46] ;
 wire \ces_5_0_io_ins_down[47] ;
 wire \ces_5_0_io_ins_down[48] ;
 wire \ces_5_0_io_ins_down[49] ;
 wire \ces_5_0_io_ins_down[4] ;
 wire \ces_5_0_io_ins_down[50] ;
 wire \ces_5_0_io_ins_down[51] ;
 wire \ces_5_0_io_ins_down[52] ;
 wire \ces_5_0_io_ins_down[53] ;
 wire \ces_5_0_io_ins_down[54] ;
 wire \ces_5_0_io_ins_down[55] ;
 wire \ces_5_0_io_ins_down[56] ;
 wire \ces_5_0_io_ins_down[57] ;
 wire \ces_5_0_io_ins_down[58] ;
 wire \ces_5_0_io_ins_down[59] ;
 wire \ces_5_0_io_ins_down[5] ;
 wire \ces_5_0_io_ins_down[60] ;
 wire \ces_5_0_io_ins_down[61] ;
 wire \ces_5_0_io_ins_down[62] ;
 wire \ces_5_0_io_ins_down[63] ;
 wire \ces_5_0_io_ins_down[6] ;
 wire \ces_5_0_io_ins_down[7] ;
 wire \ces_5_0_io_ins_down[8] ;
 wire \ces_5_0_io_ins_down[9] ;
 wire \ces_5_0_io_ins_left[0] ;
 wire \ces_5_0_io_ins_left[10] ;
 wire \ces_5_0_io_ins_left[11] ;
 wire \ces_5_0_io_ins_left[12] ;
 wire \ces_5_0_io_ins_left[13] ;
 wire \ces_5_0_io_ins_left[14] ;
 wire \ces_5_0_io_ins_left[15] ;
 wire \ces_5_0_io_ins_left[16] ;
 wire \ces_5_0_io_ins_left[17] ;
 wire \ces_5_0_io_ins_left[18] ;
 wire \ces_5_0_io_ins_left[19] ;
 wire \ces_5_0_io_ins_left[1] ;
 wire \ces_5_0_io_ins_left[20] ;
 wire \ces_5_0_io_ins_left[21] ;
 wire \ces_5_0_io_ins_left[22] ;
 wire \ces_5_0_io_ins_left[23] ;
 wire \ces_5_0_io_ins_left[24] ;
 wire \ces_5_0_io_ins_left[25] ;
 wire \ces_5_0_io_ins_left[26] ;
 wire \ces_5_0_io_ins_left[27] ;
 wire \ces_5_0_io_ins_left[28] ;
 wire \ces_5_0_io_ins_left[29] ;
 wire \ces_5_0_io_ins_left[2] ;
 wire \ces_5_0_io_ins_left[30] ;
 wire \ces_5_0_io_ins_left[31] ;
 wire \ces_5_0_io_ins_left[32] ;
 wire \ces_5_0_io_ins_left[33] ;
 wire \ces_5_0_io_ins_left[34] ;
 wire \ces_5_0_io_ins_left[35] ;
 wire \ces_5_0_io_ins_left[36] ;
 wire \ces_5_0_io_ins_left[37] ;
 wire \ces_5_0_io_ins_left[38] ;
 wire \ces_5_0_io_ins_left[39] ;
 wire \ces_5_0_io_ins_left[3] ;
 wire \ces_5_0_io_ins_left[40] ;
 wire \ces_5_0_io_ins_left[41] ;
 wire \ces_5_0_io_ins_left[42] ;
 wire \ces_5_0_io_ins_left[43] ;
 wire \ces_5_0_io_ins_left[44] ;
 wire \ces_5_0_io_ins_left[45] ;
 wire \ces_5_0_io_ins_left[46] ;
 wire \ces_5_0_io_ins_left[47] ;
 wire \ces_5_0_io_ins_left[48] ;
 wire \ces_5_0_io_ins_left[49] ;
 wire \ces_5_0_io_ins_left[4] ;
 wire \ces_5_0_io_ins_left[50] ;
 wire \ces_5_0_io_ins_left[51] ;
 wire \ces_5_0_io_ins_left[52] ;
 wire \ces_5_0_io_ins_left[53] ;
 wire \ces_5_0_io_ins_left[54] ;
 wire \ces_5_0_io_ins_left[55] ;
 wire \ces_5_0_io_ins_left[56] ;
 wire \ces_5_0_io_ins_left[57] ;
 wire \ces_5_0_io_ins_left[58] ;
 wire \ces_5_0_io_ins_left[59] ;
 wire \ces_5_0_io_ins_left[5] ;
 wire \ces_5_0_io_ins_left[60] ;
 wire \ces_5_0_io_ins_left[61] ;
 wire \ces_5_0_io_ins_left[62] ;
 wire \ces_5_0_io_ins_left[63] ;
 wire \ces_5_0_io_ins_left[6] ;
 wire \ces_5_0_io_ins_left[7] ;
 wire \ces_5_0_io_ins_left[8] ;
 wire \ces_5_0_io_ins_left[9] ;
 wire ces_5_0_io_lsbOuts_0;
 wire ces_5_0_io_lsbOuts_1;
 wire ces_5_0_io_lsbOuts_2;
 wire ces_5_0_io_lsbOuts_3;
 wire ces_5_0_io_lsbOuts_4;
 wire ces_5_0_io_lsbOuts_5;
 wire ces_5_0_io_lsbOuts_6;
 wire ces_5_0_io_lsbOuts_7;
 wire \ces_5_0_io_outs_right[0] ;
 wire \ces_5_0_io_outs_right[10] ;
 wire \ces_5_0_io_outs_right[11] ;
 wire \ces_5_0_io_outs_right[12] ;
 wire \ces_5_0_io_outs_right[13] ;
 wire \ces_5_0_io_outs_right[14] ;
 wire \ces_5_0_io_outs_right[15] ;
 wire \ces_5_0_io_outs_right[16] ;
 wire \ces_5_0_io_outs_right[17] ;
 wire \ces_5_0_io_outs_right[18] ;
 wire \ces_5_0_io_outs_right[19] ;
 wire \ces_5_0_io_outs_right[1] ;
 wire \ces_5_0_io_outs_right[20] ;
 wire \ces_5_0_io_outs_right[21] ;
 wire \ces_5_0_io_outs_right[22] ;
 wire \ces_5_0_io_outs_right[23] ;
 wire \ces_5_0_io_outs_right[24] ;
 wire \ces_5_0_io_outs_right[25] ;
 wire \ces_5_0_io_outs_right[26] ;
 wire \ces_5_0_io_outs_right[27] ;
 wire \ces_5_0_io_outs_right[28] ;
 wire \ces_5_0_io_outs_right[29] ;
 wire \ces_5_0_io_outs_right[2] ;
 wire \ces_5_0_io_outs_right[30] ;
 wire \ces_5_0_io_outs_right[31] ;
 wire \ces_5_0_io_outs_right[32] ;
 wire \ces_5_0_io_outs_right[33] ;
 wire \ces_5_0_io_outs_right[34] ;
 wire \ces_5_0_io_outs_right[35] ;
 wire \ces_5_0_io_outs_right[36] ;
 wire \ces_5_0_io_outs_right[37] ;
 wire \ces_5_0_io_outs_right[38] ;
 wire \ces_5_0_io_outs_right[39] ;
 wire \ces_5_0_io_outs_right[3] ;
 wire \ces_5_0_io_outs_right[40] ;
 wire \ces_5_0_io_outs_right[41] ;
 wire \ces_5_0_io_outs_right[42] ;
 wire \ces_5_0_io_outs_right[43] ;
 wire \ces_5_0_io_outs_right[44] ;
 wire \ces_5_0_io_outs_right[45] ;
 wire \ces_5_0_io_outs_right[46] ;
 wire \ces_5_0_io_outs_right[47] ;
 wire \ces_5_0_io_outs_right[48] ;
 wire \ces_5_0_io_outs_right[49] ;
 wire \ces_5_0_io_outs_right[4] ;
 wire \ces_5_0_io_outs_right[50] ;
 wire \ces_5_0_io_outs_right[51] ;
 wire \ces_5_0_io_outs_right[52] ;
 wire \ces_5_0_io_outs_right[53] ;
 wire \ces_5_0_io_outs_right[54] ;
 wire \ces_5_0_io_outs_right[55] ;
 wire \ces_5_0_io_outs_right[56] ;
 wire \ces_5_0_io_outs_right[57] ;
 wire \ces_5_0_io_outs_right[58] ;
 wire \ces_5_0_io_outs_right[59] ;
 wire \ces_5_0_io_outs_right[5] ;
 wire \ces_5_0_io_outs_right[60] ;
 wire \ces_5_0_io_outs_right[61] ;
 wire \ces_5_0_io_outs_right[62] ;
 wire \ces_5_0_io_outs_right[63] ;
 wire \ces_5_0_io_outs_right[6] ;
 wire \ces_5_0_io_outs_right[7] ;
 wire \ces_5_0_io_outs_right[8] ;
 wire \ces_5_0_io_outs_right[9] ;
 wire \ces_5_0_io_outs_up[0] ;
 wire \ces_5_0_io_outs_up[10] ;
 wire \ces_5_0_io_outs_up[11] ;
 wire \ces_5_0_io_outs_up[12] ;
 wire \ces_5_0_io_outs_up[13] ;
 wire \ces_5_0_io_outs_up[14] ;
 wire \ces_5_0_io_outs_up[15] ;
 wire \ces_5_0_io_outs_up[16] ;
 wire \ces_5_0_io_outs_up[17] ;
 wire \ces_5_0_io_outs_up[18] ;
 wire \ces_5_0_io_outs_up[19] ;
 wire \ces_5_0_io_outs_up[1] ;
 wire \ces_5_0_io_outs_up[20] ;
 wire \ces_5_0_io_outs_up[21] ;
 wire \ces_5_0_io_outs_up[22] ;
 wire \ces_5_0_io_outs_up[23] ;
 wire \ces_5_0_io_outs_up[24] ;
 wire \ces_5_0_io_outs_up[25] ;
 wire \ces_5_0_io_outs_up[26] ;
 wire \ces_5_0_io_outs_up[27] ;
 wire \ces_5_0_io_outs_up[28] ;
 wire \ces_5_0_io_outs_up[29] ;
 wire \ces_5_0_io_outs_up[2] ;
 wire \ces_5_0_io_outs_up[30] ;
 wire \ces_5_0_io_outs_up[31] ;
 wire \ces_5_0_io_outs_up[32] ;
 wire \ces_5_0_io_outs_up[33] ;
 wire \ces_5_0_io_outs_up[34] ;
 wire \ces_5_0_io_outs_up[35] ;
 wire \ces_5_0_io_outs_up[36] ;
 wire \ces_5_0_io_outs_up[37] ;
 wire \ces_5_0_io_outs_up[38] ;
 wire \ces_5_0_io_outs_up[39] ;
 wire \ces_5_0_io_outs_up[3] ;
 wire \ces_5_0_io_outs_up[40] ;
 wire \ces_5_0_io_outs_up[41] ;
 wire \ces_5_0_io_outs_up[42] ;
 wire \ces_5_0_io_outs_up[43] ;
 wire \ces_5_0_io_outs_up[44] ;
 wire \ces_5_0_io_outs_up[45] ;
 wire \ces_5_0_io_outs_up[46] ;
 wire \ces_5_0_io_outs_up[47] ;
 wire \ces_5_0_io_outs_up[48] ;
 wire \ces_5_0_io_outs_up[49] ;
 wire \ces_5_0_io_outs_up[4] ;
 wire \ces_5_0_io_outs_up[50] ;
 wire \ces_5_0_io_outs_up[51] ;
 wire \ces_5_0_io_outs_up[52] ;
 wire \ces_5_0_io_outs_up[53] ;
 wire \ces_5_0_io_outs_up[54] ;
 wire \ces_5_0_io_outs_up[55] ;
 wire \ces_5_0_io_outs_up[56] ;
 wire \ces_5_0_io_outs_up[57] ;
 wire \ces_5_0_io_outs_up[58] ;
 wire \ces_5_0_io_outs_up[59] ;
 wire \ces_5_0_io_outs_up[5] ;
 wire \ces_5_0_io_outs_up[60] ;
 wire \ces_5_0_io_outs_up[61] ;
 wire \ces_5_0_io_outs_up[62] ;
 wire \ces_5_0_io_outs_up[63] ;
 wire \ces_5_0_io_outs_up[6] ;
 wire \ces_5_0_io_outs_up[7] ;
 wire \ces_5_0_io_outs_up[8] ;
 wire \ces_5_0_io_outs_up[9] ;
 wire \ces_5_1_io_ins_down[0] ;
 wire \ces_5_1_io_ins_down[10] ;
 wire \ces_5_1_io_ins_down[11] ;
 wire \ces_5_1_io_ins_down[12] ;
 wire \ces_5_1_io_ins_down[13] ;
 wire \ces_5_1_io_ins_down[14] ;
 wire \ces_5_1_io_ins_down[15] ;
 wire \ces_5_1_io_ins_down[16] ;
 wire \ces_5_1_io_ins_down[17] ;
 wire \ces_5_1_io_ins_down[18] ;
 wire \ces_5_1_io_ins_down[19] ;
 wire \ces_5_1_io_ins_down[1] ;
 wire \ces_5_1_io_ins_down[20] ;
 wire \ces_5_1_io_ins_down[21] ;
 wire \ces_5_1_io_ins_down[22] ;
 wire \ces_5_1_io_ins_down[23] ;
 wire \ces_5_1_io_ins_down[24] ;
 wire \ces_5_1_io_ins_down[25] ;
 wire \ces_5_1_io_ins_down[26] ;
 wire \ces_5_1_io_ins_down[27] ;
 wire \ces_5_1_io_ins_down[28] ;
 wire \ces_5_1_io_ins_down[29] ;
 wire \ces_5_1_io_ins_down[2] ;
 wire \ces_5_1_io_ins_down[30] ;
 wire \ces_5_1_io_ins_down[31] ;
 wire \ces_5_1_io_ins_down[32] ;
 wire \ces_5_1_io_ins_down[33] ;
 wire \ces_5_1_io_ins_down[34] ;
 wire \ces_5_1_io_ins_down[35] ;
 wire \ces_5_1_io_ins_down[36] ;
 wire \ces_5_1_io_ins_down[37] ;
 wire \ces_5_1_io_ins_down[38] ;
 wire \ces_5_1_io_ins_down[39] ;
 wire \ces_5_1_io_ins_down[3] ;
 wire \ces_5_1_io_ins_down[40] ;
 wire \ces_5_1_io_ins_down[41] ;
 wire \ces_5_1_io_ins_down[42] ;
 wire \ces_5_1_io_ins_down[43] ;
 wire \ces_5_1_io_ins_down[44] ;
 wire \ces_5_1_io_ins_down[45] ;
 wire \ces_5_1_io_ins_down[46] ;
 wire \ces_5_1_io_ins_down[47] ;
 wire \ces_5_1_io_ins_down[48] ;
 wire \ces_5_1_io_ins_down[49] ;
 wire \ces_5_1_io_ins_down[4] ;
 wire \ces_5_1_io_ins_down[50] ;
 wire \ces_5_1_io_ins_down[51] ;
 wire \ces_5_1_io_ins_down[52] ;
 wire \ces_5_1_io_ins_down[53] ;
 wire \ces_5_1_io_ins_down[54] ;
 wire \ces_5_1_io_ins_down[55] ;
 wire \ces_5_1_io_ins_down[56] ;
 wire \ces_5_1_io_ins_down[57] ;
 wire \ces_5_1_io_ins_down[58] ;
 wire \ces_5_1_io_ins_down[59] ;
 wire \ces_5_1_io_ins_down[5] ;
 wire \ces_5_1_io_ins_down[60] ;
 wire \ces_5_1_io_ins_down[61] ;
 wire \ces_5_1_io_ins_down[62] ;
 wire \ces_5_1_io_ins_down[63] ;
 wire \ces_5_1_io_ins_down[6] ;
 wire \ces_5_1_io_ins_down[7] ;
 wire \ces_5_1_io_ins_down[8] ;
 wire \ces_5_1_io_ins_down[9] ;
 wire \ces_5_1_io_ins_left[0] ;
 wire \ces_5_1_io_ins_left[10] ;
 wire \ces_5_1_io_ins_left[11] ;
 wire \ces_5_1_io_ins_left[12] ;
 wire \ces_5_1_io_ins_left[13] ;
 wire \ces_5_1_io_ins_left[14] ;
 wire \ces_5_1_io_ins_left[15] ;
 wire \ces_5_1_io_ins_left[16] ;
 wire \ces_5_1_io_ins_left[17] ;
 wire \ces_5_1_io_ins_left[18] ;
 wire \ces_5_1_io_ins_left[19] ;
 wire \ces_5_1_io_ins_left[1] ;
 wire \ces_5_1_io_ins_left[20] ;
 wire \ces_5_1_io_ins_left[21] ;
 wire \ces_5_1_io_ins_left[22] ;
 wire \ces_5_1_io_ins_left[23] ;
 wire \ces_5_1_io_ins_left[24] ;
 wire \ces_5_1_io_ins_left[25] ;
 wire \ces_5_1_io_ins_left[26] ;
 wire \ces_5_1_io_ins_left[27] ;
 wire \ces_5_1_io_ins_left[28] ;
 wire \ces_5_1_io_ins_left[29] ;
 wire \ces_5_1_io_ins_left[2] ;
 wire \ces_5_1_io_ins_left[30] ;
 wire \ces_5_1_io_ins_left[31] ;
 wire \ces_5_1_io_ins_left[32] ;
 wire \ces_5_1_io_ins_left[33] ;
 wire \ces_5_1_io_ins_left[34] ;
 wire \ces_5_1_io_ins_left[35] ;
 wire \ces_5_1_io_ins_left[36] ;
 wire \ces_5_1_io_ins_left[37] ;
 wire \ces_5_1_io_ins_left[38] ;
 wire \ces_5_1_io_ins_left[39] ;
 wire \ces_5_1_io_ins_left[3] ;
 wire \ces_5_1_io_ins_left[40] ;
 wire \ces_5_1_io_ins_left[41] ;
 wire \ces_5_1_io_ins_left[42] ;
 wire \ces_5_1_io_ins_left[43] ;
 wire \ces_5_1_io_ins_left[44] ;
 wire \ces_5_1_io_ins_left[45] ;
 wire \ces_5_1_io_ins_left[46] ;
 wire \ces_5_1_io_ins_left[47] ;
 wire \ces_5_1_io_ins_left[48] ;
 wire \ces_5_1_io_ins_left[49] ;
 wire \ces_5_1_io_ins_left[4] ;
 wire \ces_5_1_io_ins_left[50] ;
 wire \ces_5_1_io_ins_left[51] ;
 wire \ces_5_1_io_ins_left[52] ;
 wire \ces_5_1_io_ins_left[53] ;
 wire \ces_5_1_io_ins_left[54] ;
 wire \ces_5_1_io_ins_left[55] ;
 wire \ces_5_1_io_ins_left[56] ;
 wire \ces_5_1_io_ins_left[57] ;
 wire \ces_5_1_io_ins_left[58] ;
 wire \ces_5_1_io_ins_left[59] ;
 wire \ces_5_1_io_ins_left[5] ;
 wire \ces_5_1_io_ins_left[60] ;
 wire \ces_5_1_io_ins_left[61] ;
 wire \ces_5_1_io_ins_left[62] ;
 wire \ces_5_1_io_ins_left[63] ;
 wire \ces_5_1_io_ins_left[6] ;
 wire \ces_5_1_io_ins_left[7] ;
 wire \ces_5_1_io_ins_left[8] ;
 wire \ces_5_1_io_ins_left[9] ;
 wire ces_5_1_io_lsbOuts_0;
 wire ces_5_1_io_lsbOuts_1;
 wire ces_5_1_io_lsbOuts_2;
 wire ces_5_1_io_lsbOuts_3;
 wire ces_5_1_io_lsbOuts_4;
 wire ces_5_1_io_lsbOuts_5;
 wire ces_5_1_io_lsbOuts_6;
 wire ces_5_1_io_lsbOuts_7;
 wire \ces_5_1_io_outs_right[0] ;
 wire \ces_5_1_io_outs_right[10] ;
 wire \ces_5_1_io_outs_right[11] ;
 wire \ces_5_1_io_outs_right[12] ;
 wire \ces_5_1_io_outs_right[13] ;
 wire \ces_5_1_io_outs_right[14] ;
 wire \ces_5_1_io_outs_right[15] ;
 wire \ces_5_1_io_outs_right[16] ;
 wire \ces_5_1_io_outs_right[17] ;
 wire \ces_5_1_io_outs_right[18] ;
 wire \ces_5_1_io_outs_right[19] ;
 wire \ces_5_1_io_outs_right[1] ;
 wire \ces_5_1_io_outs_right[20] ;
 wire \ces_5_1_io_outs_right[21] ;
 wire \ces_5_1_io_outs_right[22] ;
 wire \ces_5_1_io_outs_right[23] ;
 wire \ces_5_1_io_outs_right[24] ;
 wire \ces_5_1_io_outs_right[25] ;
 wire \ces_5_1_io_outs_right[26] ;
 wire \ces_5_1_io_outs_right[27] ;
 wire \ces_5_1_io_outs_right[28] ;
 wire \ces_5_1_io_outs_right[29] ;
 wire \ces_5_1_io_outs_right[2] ;
 wire \ces_5_1_io_outs_right[30] ;
 wire \ces_5_1_io_outs_right[31] ;
 wire \ces_5_1_io_outs_right[32] ;
 wire \ces_5_1_io_outs_right[33] ;
 wire \ces_5_1_io_outs_right[34] ;
 wire \ces_5_1_io_outs_right[35] ;
 wire \ces_5_1_io_outs_right[36] ;
 wire \ces_5_1_io_outs_right[37] ;
 wire \ces_5_1_io_outs_right[38] ;
 wire \ces_5_1_io_outs_right[39] ;
 wire \ces_5_1_io_outs_right[3] ;
 wire \ces_5_1_io_outs_right[40] ;
 wire \ces_5_1_io_outs_right[41] ;
 wire \ces_5_1_io_outs_right[42] ;
 wire \ces_5_1_io_outs_right[43] ;
 wire \ces_5_1_io_outs_right[44] ;
 wire \ces_5_1_io_outs_right[45] ;
 wire \ces_5_1_io_outs_right[46] ;
 wire \ces_5_1_io_outs_right[47] ;
 wire \ces_5_1_io_outs_right[48] ;
 wire \ces_5_1_io_outs_right[49] ;
 wire \ces_5_1_io_outs_right[4] ;
 wire \ces_5_1_io_outs_right[50] ;
 wire \ces_5_1_io_outs_right[51] ;
 wire \ces_5_1_io_outs_right[52] ;
 wire \ces_5_1_io_outs_right[53] ;
 wire \ces_5_1_io_outs_right[54] ;
 wire \ces_5_1_io_outs_right[55] ;
 wire \ces_5_1_io_outs_right[56] ;
 wire \ces_5_1_io_outs_right[57] ;
 wire \ces_5_1_io_outs_right[58] ;
 wire \ces_5_1_io_outs_right[59] ;
 wire \ces_5_1_io_outs_right[5] ;
 wire \ces_5_1_io_outs_right[60] ;
 wire \ces_5_1_io_outs_right[61] ;
 wire \ces_5_1_io_outs_right[62] ;
 wire \ces_5_1_io_outs_right[63] ;
 wire \ces_5_1_io_outs_right[6] ;
 wire \ces_5_1_io_outs_right[7] ;
 wire \ces_5_1_io_outs_right[8] ;
 wire \ces_5_1_io_outs_right[9] ;
 wire \ces_5_1_io_outs_up[0] ;
 wire \ces_5_1_io_outs_up[10] ;
 wire \ces_5_1_io_outs_up[11] ;
 wire \ces_5_1_io_outs_up[12] ;
 wire \ces_5_1_io_outs_up[13] ;
 wire \ces_5_1_io_outs_up[14] ;
 wire \ces_5_1_io_outs_up[15] ;
 wire \ces_5_1_io_outs_up[16] ;
 wire \ces_5_1_io_outs_up[17] ;
 wire \ces_5_1_io_outs_up[18] ;
 wire \ces_5_1_io_outs_up[19] ;
 wire \ces_5_1_io_outs_up[1] ;
 wire \ces_5_1_io_outs_up[20] ;
 wire \ces_5_1_io_outs_up[21] ;
 wire \ces_5_1_io_outs_up[22] ;
 wire \ces_5_1_io_outs_up[23] ;
 wire \ces_5_1_io_outs_up[24] ;
 wire \ces_5_1_io_outs_up[25] ;
 wire \ces_5_1_io_outs_up[26] ;
 wire \ces_5_1_io_outs_up[27] ;
 wire \ces_5_1_io_outs_up[28] ;
 wire \ces_5_1_io_outs_up[29] ;
 wire \ces_5_1_io_outs_up[2] ;
 wire \ces_5_1_io_outs_up[30] ;
 wire \ces_5_1_io_outs_up[31] ;
 wire \ces_5_1_io_outs_up[32] ;
 wire \ces_5_1_io_outs_up[33] ;
 wire \ces_5_1_io_outs_up[34] ;
 wire \ces_5_1_io_outs_up[35] ;
 wire \ces_5_1_io_outs_up[36] ;
 wire \ces_5_1_io_outs_up[37] ;
 wire \ces_5_1_io_outs_up[38] ;
 wire \ces_5_1_io_outs_up[39] ;
 wire \ces_5_1_io_outs_up[3] ;
 wire \ces_5_1_io_outs_up[40] ;
 wire \ces_5_1_io_outs_up[41] ;
 wire \ces_5_1_io_outs_up[42] ;
 wire \ces_5_1_io_outs_up[43] ;
 wire \ces_5_1_io_outs_up[44] ;
 wire \ces_5_1_io_outs_up[45] ;
 wire \ces_5_1_io_outs_up[46] ;
 wire \ces_5_1_io_outs_up[47] ;
 wire \ces_5_1_io_outs_up[48] ;
 wire \ces_5_1_io_outs_up[49] ;
 wire \ces_5_1_io_outs_up[4] ;
 wire \ces_5_1_io_outs_up[50] ;
 wire \ces_5_1_io_outs_up[51] ;
 wire \ces_5_1_io_outs_up[52] ;
 wire \ces_5_1_io_outs_up[53] ;
 wire \ces_5_1_io_outs_up[54] ;
 wire \ces_5_1_io_outs_up[55] ;
 wire \ces_5_1_io_outs_up[56] ;
 wire \ces_5_1_io_outs_up[57] ;
 wire \ces_5_1_io_outs_up[58] ;
 wire \ces_5_1_io_outs_up[59] ;
 wire \ces_5_1_io_outs_up[5] ;
 wire \ces_5_1_io_outs_up[60] ;
 wire \ces_5_1_io_outs_up[61] ;
 wire \ces_5_1_io_outs_up[62] ;
 wire \ces_5_1_io_outs_up[63] ;
 wire \ces_5_1_io_outs_up[6] ;
 wire \ces_5_1_io_outs_up[7] ;
 wire \ces_5_1_io_outs_up[8] ;
 wire \ces_5_1_io_outs_up[9] ;
 wire \ces_5_2_io_ins_down[0] ;
 wire \ces_5_2_io_ins_down[10] ;
 wire \ces_5_2_io_ins_down[11] ;
 wire \ces_5_2_io_ins_down[12] ;
 wire \ces_5_2_io_ins_down[13] ;
 wire \ces_5_2_io_ins_down[14] ;
 wire \ces_5_2_io_ins_down[15] ;
 wire \ces_5_2_io_ins_down[16] ;
 wire \ces_5_2_io_ins_down[17] ;
 wire \ces_5_2_io_ins_down[18] ;
 wire \ces_5_2_io_ins_down[19] ;
 wire \ces_5_2_io_ins_down[1] ;
 wire \ces_5_2_io_ins_down[20] ;
 wire \ces_5_2_io_ins_down[21] ;
 wire \ces_5_2_io_ins_down[22] ;
 wire \ces_5_2_io_ins_down[23] ;
 wire \ces_5_2_io_ins_down[24] ;
 wire \ces_5_2_io_ins_down[25] ;
 wire \ces_5_2_io_ins_down[26] ;
 wire \ces_5_2_io_ins_down[27] ;
 wire \ces_5_2_io_ins_down[28] ;
 wire \ces_5_2_io_ins_down[29] ;
 wire \ces_5_2_io_ins_down[2] ;
 wire \ces_5_2_io_ins_down[30] ;
 wire \ces_5_2_io_ins_down[31] ;
 wire \ces_5_2_io_ins_down[32] ;
 wire \ces_5_2_io_ins_down[33] ;
 wire \ces_5_2_io_ins_down[34] ;
 wire \ces_5_2_io_ins_down[35] ;
 wire \ces_5_2_io_ins_down[36] ;
 wire \ces_5_2_io_ins_down[37] ;
 wire \ces_5_2_io_ins_down[38] ;
 wire \ces_5_2_io_ins_down[39] ;
 wire \ces_5_2_io_ins_down[3] ;
 wire \ces_5_2_io_ins_down[40] ;
 wire \ces_5_2_io_ins_down[41] ;
 wire \ces_5_2_io_ins_down[42] ;
 wire \ces_5_2_io_ins_down[43] ;
 wire \ces_5_2_io_ins_down[44] ;
 wire \ces_5_2_io_ins_down[45] ;
 wire \ces_5_2_io_ins_down[46] ;
 wire \ces_5_2_io_ins_down[47] ;
 wire \ces_5_2_io_ins_down[48] ;
 wire \ces_5_2_io_ins_down[49] ;
 wire \ces_5_2_io_ins_down[4] ;
 wire \ces_5_2_io_ins_down[50] ;
 wire \ces_5_2_io_ins_down[51] ;
 wire \ces_5_2_io_ins_down[52] ;
 wire \ces_5_2_io_ins_down[53] ;
 wire \ces_5_2_io_ins_down[54] ;
 wire \ces_5_2_io_ins_down[55] ;
 wire \ces_5_2_io_ins_down[56] ;
 wire \ces_5_2_io_ins_down[57] ;
 wire \ces_5_2_io_ins_down[58] ;
 wire \ces_5_2_io_ins_down[59] ;
 wire \ces_5_2_io_ins_down[5] ;
 wire \ces_5_2_io_ins_down[60] ;
 wire \ces_5_2_io_ins_down[61] ;
 wire \ces_5_2_io_ins_down[62] ;
 wire \ces_5_2_io_ins_down[63] ;
 wire \ces_5_2_io_ins_down[6] ;
 wire \ces_5_2_io_ins_down[7] ;
 wire \ces_5_2_io_ins_down[8] ;
 wire \ces_5_2_io_ins_down[9] ;
 wire \ces_5_2_io_ins_left[0] ;
 wire \ces_5_2_io_ins_left[10] ;
 wire \ces_5_2_io_ins_left[11] ;
 wire \ces_5_2_io_ins_left[12] ;
 wire \ces_5_2_io_ins_left[13] ;
 wire \ces_5_2_io_ins_left[14] ;
 wire \ces_5_2_io_ins_left[15] ;
 wire \ces_5_2_io_ins_left[16] ;
 wire \ces_5_2_io_ins_left[17] ;
 wire \ces_5_2_io_ins_left[18] ;
 wire \ces_5_2_io_ins_left[19] ;
 wire \ces_5_2_io_ins_left[1] ;
 wire \ces_5_2_io_ins_left[20] ;
 wire \ces_5_2_io_ins_left[21] ;
 wire \ces_5_2_io_ins_left[22] ;
 wire \ces_5_2_io_ins_left[23] ;
 wire \ces_5_2_io_ins_left[24] ;
 wire \ces_5_2_io_ins_left[25] ;
 wire \ces_5_2_io_ins_left[26] ;
 wire \ces_5_2_io_ins_left[27] ;
 wire \ces_5_2_io_ins_left[28] ;
 wire \ces_5_2_io_ins_left[29] ;
 wire \ces_5_2_io_ins_left[2] ;
 wire \ces_5_2_io_ins_left[30] ;
 wire \ces_5_2_io_ins_left[31] ;
 wire \ces_5_2_io_ins_left[32] ;
 wire \ces_5_2_io_ins_left[33] ;
 wire \ces_5_2_io_ins_left[34] ;
 wire \ces_5_2_io_ins_left[35] ;
 wire \ces_5_2_io_ins_left[36] ;
 wire \ces_5_2_io_ins_left[37] ;
 wire \ces_5_2_io_ins_left[38] ;
 wire \ces_5_2_io_ins_left[39] ;
 wire \ces_5_2_io_ins_left[3] ;
 wire \ces_5_2_io_ins_left[40] ;
 wire \ces_5_2_io_ins_left[41] ;
 wire \ces_5_2_io_ins_left[42] ;
 wire \ces_5_2_io_ins_left[43] ;
 wire \ces_5_2_io_ins_left[44] ;
 wire \ces_5_2_io_ins_left[45] ;
 wire \ces_5_2_io_ins_left[46] ;
 wire \ces_5_2_io_ins_left[47] ;
 wire \ces_5_2_io_ins_left[48] ;
 wire \ces_5_2_io_ins_left[49] ;
 wire \ces_5_2_io_ins_left[4] ;
 wire \ces_5_2_io_ins_left[50] ;
 wire \ces_5_2_io_ins_left[51] ;
 wire \ces_5_2_io_ins_left[52] ;
 wire \ces_5_2_io_ins_left[53] ;
 wire \ces_5_2_io_ins_left[54] ;
 wire \ces_5_2_io_ins_left[55] ;
 wire \ces_5_2_io_ins_left[56] ;
 wire \ces_5_2_io_ins_left[57] ;
 wire \ces_5_2_io_ins_left[58] ;
 wire \ces_5_2_io_ins_left[59] ;
 wire \ces_5_2_io_ins_left[5] ;
 wire \ces_5_2_io_ins_left[60] ;
 wire \ces_5_2_io_ins_left[61] ;
 wire \ces_5_2_io_ins_left[62] ;
 wire \ces_5_2_io_ins_left[63] ;
 wire \ces_5_2_io_ins_left[6] ;
 wire \ces_5_2_io_ins_left[7] ;
 wire \ces_5_2_io_ins_left[8] ;
 wire \ces_5_2_io_ins_left[9] ;
 wire ces_5_2_io_lsbOuts_0;
 wire ces_5_2_io_lsbOuts_1;
 wire ces_5_2_io_lsbOuts_2;
 wire ces_5_2_io_lsbOuts_3;
 wire ces_5_2_io_lsbOuts_4;
 wire ces_5_2_io_lsbOuts_5;
 wire ces_5_2_io_lsbOuts_6;
 wire ces_5_2_io_lsbOuts_7;
 wire \ces_5_2_io_outs_right[0] ;
 wire \ces_5_2_io_outs_right[10] ;
 wire \ces_5_2_io_outs_right[11] ;
 wire \ces_5_2_io_outs_right[12] ;
 wire \ces_5_2_io_outs_right[13] ;
 wire \ces_5_2_io_outs_right[14] ;
 wire \ces_5_2_io_outs_right[15] ;
 wire \ces_5_2_io_outs_right[16] ;
 wire \ces_5_2_io_outs_right[17] ;
 wire \ces_5_2_io_outs_right[18] ;
 wire \ces_5_2_io_outs_right[19] ;
 wire \ces_5_2_io_outs_right[1] ;
 wire \ces_5_2_io_outs_right[20] ;
 wire \ces_5_2_io_outs_right[21] ;
 wire \ces_5_2_io_outs_right[22] ;
 wire \ces_5_2_io_outs_right[23] ;
 wire \ces_5_2_io_outs_right[24] ;
 wire \ces_5_2_io_outs_right[25] ;
 wire \ces_5_2_io_outs_right[26] ;
 wire \ces_5_2_io_outs_right[27] ;
 wire \ces_5_2_io_outs_right[28] ;
 wire \ces_5_2_io_outs_right[29] ;
 wire \ces_5_2_io_outs_right[2] ;
 wire \ces_5_2_io_outs_right[30] ;
 wire \ces_5_2_io_outs_right[31] ;
 wire \ces_5_2_io_outs_right[32] ;
 wire \ces_5_2_io_outs_right[33] ;
 wire \ces_5_2_io_outs_right[34] ;
 wire \ces_5_2_io_outs_right[35] ;
 wire \ces_5_2_io_outs_right[36] ;
 wire \ces_5_2_io_outs_right[37] ;
 wire \ces_5_2_io_outs_right[38] ;
 wire \ces_5_2_io_outs_right[39] ;
 wire \ces_5_2_io_outs_right[3] ;
 wire \ces_5_2_io_outs_right[40] ;
 wire \ces_5_2_io_outs_right[41] ;
 wire \ces_5_2_io_outs_right[42] ;
 wire \ces_5_2_io_outs_right[43] ;
 wire \ces_5_2_io_outs_right[44] ;
 wire \ces_5_2_io_outs_right[45] ;
 wire \ces_5_2_io_outs_right[46] ;
 wire \ces_5_2_io_outs_right[47] ;
 wire \ces_5_2_io_outs_right[48] ;
 wire \ces_5_2_io_outs_right[49] ;
 wire \ces_5_2_io_outs_right[4] ;
 wire \ces_5_2_io_outs_right[50] ;
 wire \ces_5_2_io_outs_right[51] ;
 wire \ces_5_2_io_outs_right[52] ;
 wire \ces_5_2_io_outs_right[53] ;
 wire \ces_5_2_io_outs_right[54] ;
 wire \ces_5_2_io_outs_right[55] ;
 wire \ces_5_2_io_outs_right[56] ;
 wire \ces_5_2_io_outs_right[57] ;
 wire \ces_5_2_io_outs_right[58] ;
 wire \ces_5_2_io_outs_right[59] ;
 wire \ces_5_2_io_outs_right[5] ;
 wire \ces_5_2_io_outs_right[60] ;
 wire \ces_5_2_io_outs_right[61] ;
 wire \ces_5_2_io_outs_right[62] ;
 wire \ces_5_2_io_outs_right[63] ;
 wire \ces_5_2_io_outs_right[6] ;
 wire \ces_5_2_io_outs_right[7] ;
 wire \ces_5_2_io_outs_right[8] ;
 wire \ces_5_2_io_outs_right[9] ;
 wire \ces_5_2_io_outs_up[0] ;
 wire \ces_5_2_io_outs_up[10] ;
 wire \ces_5_2_io_outs_up[11] ;
 wire \ces_5_2_io_outs_up[12] ;
 wire \ces_5_2_io_outs_up[13] ;
 wire \ces_5_2_io_outs_up[14] ;
 wire \ces_5_2_io_outs_up[15] ;
 wire \ces_5_2_io_outs_up[16] ;
 wire \ces_5_2_io_outs_up[17] ;
 wire \ces_5_2_io_outs_up[18] ;
 wire \ces_5_2_io_outs_up[19] ;
 wire \ces_5_2_io_outs_up[1] ;
 wire \ces_5_2_io_outs_up[20] ;
 wire \ces_5_2_io_outs_up[21] ;
 wire \ces_5_2_io_outs_up[22] ;
 wire \ces_5_2_io_outs_up[23] ;
 wire \ces_5_2_io_outs_up[24] ;
 wire \ces_5_2_io_outs_up[25] ;
 wire \ces_5_2_io_outs_up[26] ;
 wire \ces_5_2_io_outs_up[27] ;
 wire \ces_5_2_io_outs_up[28] ;
 wire \ces_5_2_io_outs_up[29] ;
 wire \ces_5_2_io_outs_up[2] ;
 wire \ces_5_2_io_outs_up[30] ;
 wire \ces_5_2_io_outs_up[31] ;
 wire \ces_5_2_io_outs_up[32] ;
 wire \ces_5_2_io_outs_up[33] ;
 wire \ces_5_2_io_outs_up[34] ;
 wire \ces_5_2_io_outs_up[35] ;
 wire \ces_5_2_io_outs_up[36] ;
 wire \ces_5_2_io_outs_up[37] ;
 wire \ces_5_2_io_outs_up[38] ;
 wire \ces_5_2_io_outs_up[39] ;
 wire \ces_5_2_io_outs_up[3] ;
 wire \ces_5_2_io_outs_up[40] ;
 wire \ces_5_2_io_outs_up[41] ;
 wire \ces_5_2_io_outs_up[42] ;
 wire \ces_5_2_io_outs_up[43] ;
 wire \ces_5_2_io_outs_up[44] ;
 wire \ces_5_2_io_outs_up[45] ;
 wire \ces_5_2_io_outs_up[46] ;
 wire \ces_5_2_io_outs_up[47] ;
 wire \ces_5_2_io_outs_up[48] ;
 wire \ces_5_2_io_outs_up[49] ;
 wire \ces_5_2_io_outs_up[4] ;
 wire \ces_5_2_io_outs_up[50] ;
 wire \ces_5_2_io_outs_up[51] ;
 wire \ces_5_2_io_outs_up[52] ;
 wire \ces_5_2_io_outs_up[53] ;
 wire \ces_5_2_io_outs_up[54] ;
 wire \ces_5_2_io_outs_up[55] ;
 wire \ces_5_2_io_outs_up[56] ;
 wire \ces_5_2_io_outs_up[57] ;
 wire \ces_5_2_io_outs_up[58] ;
 wire \ces_5_2_io_outs_up[59] ;
 wire \ces_5_2_io_outs_up[5] ;
 wire \ces_5_2_io_outs_up[60] ;
 wire \ces_5_2_io_outs_up[61] ;
 wire \ces_5_2_io_outs_up[62] ;
 wire \ces_5_2_io_outs_up[63] ;
 wire \ces_5_2_io_outs_up[6] ;
 wire \ces_5_2_io_outs_up[7] ;
 wire \ces_5_2_io_outs_up[8] ;
 wire \ces_5_2_io_outs_up[9] ;
 wire \ces_5_3_io_ins_down[0] ;
 wire \ces_5_3_io_ins_down[10] ;
 wire \ces_5_3_io_ins_down[11] ;
 wire \ces_5_3_io_ins_down[12] ;
 wire \ces_5_3_io_ins_down[13] ;
 wire \ces_5_3_io_ins_down[14] ;
 wire \ces_5_3_io_ins_down[15] ;
 wire \ces_5_3_io_ins_down[16] ;
 wire \ces_5_3_io_ins_down[17] ;
 wire \ces_5_3_io_ins_down[18] ;
 wire \ces_5_3_io_ins_down[19] ;
 wire \ces_5_3_io_ins_down[1] ;
 wire \ces_5_3_io_ins_down[20] ;
 wire \ces_5_3_io_ins_down[21] ;
 wire \ces_5_3_io_ins_down[22] ;
 wire \ces_5_3_io_ins_down[23] ;
 wire \ces_5_3_io_ins_down[24] ;
 wire \ces_5_3_io_ins_down[25] ;
 wire \ces_5_3_io_ins_down[26] ;
 wire \ces_5_3_io_ins_down[27] ;
 wire \ces_5_3_io_ins_down[28] ;
 wire \ces_5_3_io_ins_down[29] ;
 wire \ces_5_3_io_ins_down[2] ;
 wire \ces_5_3_io_ins_down[30] ;
 wire \ces_5_3_io_ins_down[31] ;
 wire \ces_5_3_io_ins_down[32] ;
 wire \ces_5_3_io_ins_down[33] ;
 wire \ces_5_3_io_ins_down[34] ;
 wire \ces_5_3_io_ins_down[35] ;
 wire \ces_5_3_io_ins_down[36] ;
 wire \ces_5_3_io_ins_down[37] ;
 wire \ces_5_3_io_ins_down[38] ;
 wire \ces_5_3_io_ins_down[39] ;
 wire \ces_5_3_io_ins_down[3] ;
 wire \ces_5_3_io_ins_down[40] ;
 wire \ces_5_3_io_ins_down[41] ;
 wire \ces_5_3_io_ins_down[42] ;
 wire \ces_5_3_io_ins_down[43] ;
 wire \ces_5_3_io_ins_down[44] ;
 wire \ces_5_3_io_ins_down[45] ;
 wire \ces_5_3_io_ins_down[46] ;
 wire \ces_5_3_io_ins_down[47] ;
 wire \ces_5_3_io_ins_down[48] ;
 wire \ces_5_3_io_ins_down[49] ;
 wire \ces_5_3_io_ins_down[4] ;
 wire \ces_5_3_io_ins_down[50] ;
 wire \ces_5_3_io_ins_down[51] ;
 wire \ces_5_3_io_ins_down[52] ;
 wire \ces_5_3_io_ins_down[53] ;
 wire \ces_5_3_io_ins_down[54] ;
 wire \ces_5_3_io_ins_down[55] ;
 wire \ces_5_3_io_ins_down[56] ;
 wire \ces_5_3_io_ins_down[57] ;
 wire \ces_5_3_io_ins_down[58] ;
 wire \ces_5_3_io_ins_down[59] ;
 wire \ces_5_3_io_ins_down[5] ;
 wire \ces_5_3_io_ins_down[60] ;
 wire \ces_5_3_io_ins_down[61] ;
 wire \ces_5_3_io_ins_down[62] ;
 wire \ces_5_3_io_ins_down[63] ;
 wire \ces_5_3_io_ins_down[6] ;
 wire \ces_5_3_io_ins_down[7] ;
 wire \ces_5_3_io_ins_down[8] ;
 wire \ces_5_3_io_ins_down[9] ;
 wire \ces_5_3_io_ins_left[0] ;
 wire \ces_5_3_io_ins_left[10] ;
 wire \ces_5_3_io_ins_left[11] ;
 wire \ces_5_3_io_ins_left[12] ;
 wire \ces_5_3_io_ins_left[13] ;
 wire \ces_5_3_io_ins_left[14] ;
 wire \ces_5_3_io_ins_left[15] ;
 wire \ces_5_3_io_ins_left[16] ;
 wire \ces_5_3_io_ins_left[17] ;
 wire \ces_5_3_io_ins_left[18] ;
 wire \ces_5_3_io_ins_left[19] ;
 wire \ces_5_3_io_ins_left[1] ;
 wire \ces_5_3_io_ins_left[20] ;
 wire \ces_5_3_io_ins_left[21] ;
 wire \ces_5_3_io_ins_left[22] ;
 wire \ces_5_3_io_ins_left[23] ;
 wire \ces_5_3_io_ins_left[24] ;
 wire \ces_5_3_io_ins_left[25] ;
 wire \ces_5_3_io_ins_left[26] ;
 wire \ces_5_3_io_ins_left[27] ;
 wire \ces_5_3_io_ins_left[28] ;
 wire \ces_5_3_io_ins_left[29] ;
 wire \ces_5_3_io_ins_left[2] ;
 wire \ces_5_3_io_ins_left[30] ;
 wire \ces_5_3_io_ins_left[31] ;
 wire \ces_5_3_io_ins_left[32] ;
 wire \ces_5_3_io_ins_left[33] ;
 wire \ces_5_3_io_ins_left[34] ;
 wire \ces_5_3_io_ins_left[35] ;
 wire \ces_5_3_io_ins_left[36] ;
 wire \ces_5_3_io_ins_left[37] ;
 wire \ces_5_3_io_ins_left[38] ;
 wire \ces_5_3_io_ins_left[39] ;
 wire \ces_5_3_io_ins_left[3] ;
 wire \ces_5_3_io_ins_left[40] ;
 wire \ces_5_3_io_ins_left[41] ;
 wire \ces_5_3_io_ins_left[42] ;
 wire \ces_5_3_io_ins_left[43] ;
 wire \ces_5_3_io_ins_left[44] ;
 wire \ces_5_3_io_ins_left[45] ;
 wire \ces_5_3_io_ins_left[46] ;
 wire \ces_5_3_io_ins_left[47] ;
 wire \ces_5_3_io_ins_left[48] ;
 wire \ces_5_3_io_ins_left[49] ;
 wire \ces_5_3_io_ins_left[4] ;
 wire \ces_5_3_io_ins_left[50] ;
 wire \ces_5_3_io_ins_left[51] ;
 wire \ces_5_3_io_ins_left[52] ;
 wire \ces_5_3_io_ins_left[53] ;
 wire \ces_5_3_io_ins_left[54] ;
 wire \ces_5_3_io_ins_left[55] ;
 wire \ces_5_3_io_ins_left[56] ;
 wire \ces_5_3_io_ins_left[57] ;
 wire \ces_5_3_io_ins_left[58] ;
 wire \ces_5_3_io_ins_left[59] ;
 wire \ces_5_3_io_ins_left[5] ;
 wire \ces_5_3_io_ins_left[60] ;
 wire \ces_5_3_io_ins_left[61] ;
 wire \ces_5_3_io_ins_left[62] ;
 wire \ces_5_3_io_ins_left[63] ;
 wire \ces_5_3_io_ins_left[6] ;
 wire \ces_5_3_io_ins_left[7] ;
 wire \ces_5_3_io_ins_left[8] ;
 wire \ces_5_3_io_ins_left[9] ;
 wire ces_5_3_io_lsbOuts_0;
 wire ces_5_3_io_lsbOuts_1;
 wire ces_5_3_io_lsbOuts_2;
 wire ces_5_3_io_lsbOuts_3;
 wire ces_5_3_io_lsbOuts_4;
 wire ces_5_3_io_lsbOuts_5;
 wire ces_5_3_io_lsbOuts_6;
 wire ces_5_3_io_lsbOuts_7;
 wire \ces_5_3_io_outs_right[0] ;
 wire \ces_5_3_io_outs_right[10] ;
 wire \ces_5_3_io_outs_right[11] ;
 wire \ces_5_3_io_outs_right[12] ;
 wire \ces_5_3_io_outs_right[13] ;
 wire \ces_5_3_io_outs_right[14] ;
 wire \ces_5_3_io_outs_right[15] ;
 wire \ces_5_3_io_outs_right[16] ;
 wire \ces_5_3_io_outs_right[17] ;
 wire \ces_5_3_io_outs_right[18] ;
 wire \ces_5_3_io_outs_right[19] ;
 wire \ces_5_3_io_outs_right[1] ;
 wire \ces_5_3_io_outs_right[20] ;
 wire \ces_5_3_io_outs_right[21] ;
 wire \ces_5_3_io_outs_right[22] ;
 wire \ces_5_3_io_outs_right[23] ;
 wire \ces_5_3_io_outs_right[24] ;
 wire \ces_5_3_io_outs_right[25] ;
 wire \ces_5_3_io_outs_right[26] ;
 wire \ces_5_3_io_outs_right[27] ;
 wire \ces_5_3_io_outs_right[28] ;
 wire \ces_5_3_io_outs_right[29] ;
 wire \ces_5_3_io_outs_right[2] ;
 wire \ces_5_3_io_outs_right[30] ;
 wire \ces_5_3_io_outs_right[31] ;
 wire \ces_5_3_io_outs_right[32] ;
 wire \ces_5_3_io_outs_right[33] ;
 wire \ces_5_3_io_outs_right[34] ;
 wire \ces_5_3_io_outs_right[35] ;
 wire \ces_5_3_io_outs_right[36] ;
 wire \ces_5_3_io_outs_right[37] ;
 wire \ces_5_3_io_outs_right[38] ;
 wire \ces_5_3_io_outs_right[39] ;
 wire \ces_5_3_io_outs_right[3] ;
 wire \ces_5_3_io_outs_right[40] ;
 wire \ces_5_3_io_outs_right[41] ;
 wire \ces_5_3_io_outs_right[42] ;
 wire \ces_5_3_io_outs_right[43] ;
 wire \ces_5_3_io_outs_right[44] ;
 wire \ces_5_3_io_outs_right[45] ;
 wire \ces_5_3_io_outs_right[46] ;
 wire \ces_5_3_io_outs_right[47] ;
 wire \ces_5_3_io_outs_right[48] ;
 wire \ces_5_3_io_outs_right[49] ;
 wire \ces_5_3_io_outs_right[4] ;
 wire \ces_5_3_io_outs_right[50] ;
 wire \ces_5_3_io_outs_right[51] ;
 wire \ces_5_3_io_outs_right[52] ;
 wire \ces_5_3_io_outs_right[53] ;
 wire \ces_5_3_io_outs_right[54] ;
 wire \ces_5_3_io_outs_right[55] ;
 wire \ces_5_3_io_outs_right[56] ;
 wire \ces_5_3_io_outs_right[57] ;
 wire \ces_5_3_io_outs_right[58] ;
 wire \ces_5_3_io_outs_right[59] ;
 wire \ces_5_3_io_outs_right[5] ;
 wire \ces_5_3_io_outs_right[60] ;
 wire \ces_5_3_io_outs_right[61] ;
 wire \ces_5_3_io_outs_right[62] ;
 wire \ces_5_3_io_outs_right[63] ;
 wire \ces_5_3_io_outs_right[6] ;
 wire \ces_5_3_io_outs_right[7] ;
 wire \ces_5_3_io_outs_right[8] ;
 wire \ces_5_3_io_outs_right[9] ;
 wire \ces_5_3_io_outs_up[0] ;
 wire \ces_5_3_io_outs_up[10] ;
 wire \ces_5_3_io_outs_up[11] ;
 wire \ces_5_3_io_outs_up[12] ;
 wire \ces_5_3_io_outs_up[13] ;
 wire \ces_5_3_io_outs_up[14] ;
 wire \ces_5_3_io_outs_up[15] ;
 wire \ces_5_3_io_outs_up[16] ;
 wire \ces_5_3_io_outs_up[17] ;
 wire \ces_5_3_io_outs_up[18] ;
 wire \ces_5_3_io_outs_up[19] ;
 wire \ces_5_3_io_outs_up[1] ;
 wire \ces_5_3_io_outs_up[20] ;
 wire \ces_5_3_io_outs_up[21] ;
 wire \ces_5_3_io_outs_up[22] ;
 wire \ces_5_3_io_outs_up[23] ;
 wire \ces_5_3_io_outs_up[24] ;
 wire \ces_5_3_io_outs_up[25] ;
 wire \ces_5_3_io_outs_up[26] ;
 wire \ces_5_3_io_outs_up[27] ;
 wire \ces_5_3_io_outs_up[28] ;
 wire \ces_5_3_io_outs_up[29] ;
 wire \ces_5_3_io_outs_up[2] ;
 wire \ces_5_3_io_outs_up[30] ;
 wire \ces_5_3_io_outs_up[31] ;
 wire \ces_5_3_io_outs_up[32] ;
 wire \ces_5_3_io_outs_up[33] ;
 wire \ces_5_3_io_outs_up[34] ;
 wire \ces_5_3_io_outs_up[35] ;
 wire \ces_5_3_io_outs_up[36] ;
 wire \ces_5_3_io_outs_up[37] ;
 wire \ces_5_3_io_outs_up[38] ;
 wire \ces_5_3_io_outs_up[39] ;
 wire \ces_5_3_io_outs_up[3] ;
 wire \ces_5_3_io_outs_up[40] ;
 wire \ces_5_3_io_outs_up[41] ;
 wire \ces_5_3_io_outs_up[42] ;
 wire \ces_5_3_io_outs_up[43] ;
 wire \ces_5_3_io_outs_up[44] ;
 wire \ces_5_3_io_outs_up[45] ;
 wire \ces_5_3_io_outs_up[46] ;
 wire \ces_5_3_io_outs_up[47] ;
 wire \ces_5_3_io_outs_up[48] ;
 wire \ces_5_3_io_outs_up[49] ;
 wire \ces_5_3_io_outs_up[4] ;
 wire \ces_5_3_io_outs_up[50] ;
 wire \ces_5_3_io_outs_up[51] ;
 wire \ces_5_3_io_outs_up[52] ;
 wire \ces_5_3_io_outs_up[53] ;
 wire \ces_5_3_io_outs_up[54] ;
 wire \ces_5_3_io_outs_up[55] ;
 wire \ces_5_3_io_outs_up[56] ;
 wire \ces_5_3_io_outs_up[57] ;
 wire \ces_5_3_io_outs_up[58] ;
 wire \ces_5_3_io_outs_up[59] ;
 wire \ces_5_3_io_outs_up[5] ;
 wire \ces_5_3_io_outs_up[60] ;
 wire \ces_5_3_io_outs_up[61] ;
 wire \ces_5_3_io_outs_up[62] ;
 wire \ces_5_3_io_outs_up[63] ;
 wire \ces_5_3_io_outs_up[6] ;
 wire \ces_5_3_io_outs_up[7] ;
 wire \ces_5_3_io_outs_up[8] ;
 wire \ces_5_3_io_outs_up[9] ;
 wire \ces_5_4_io_ins_down[0] ;
 wire \ces_5_4_io_ins_down[10] ;
 wire \ces_5_4_io_ins_down[11] ;
 wire \ces_5_4_io_ins_down[12] ;
 wire \ces_5_4_io_ins_down[13] ;
 wire \ces_5_4_io_ins_down[14] ;
 wire \ces_5_4_io_ins_down[15] ;
 wire \ces_5_4_io_ins_down[16] ;
 wire \ces_5_4_io_ins_down[17] ;
 wire \ces_5_4_io_ins_down[18] ;
 wire \ces_5_4_io_ins_down[19] ;
 wire \ces_5_4_io_ins_down[1] ;
 wire \ces_5_4_io_ins_down[20] ;
 wire \ces_5_4_io_ins_down[21] ;
 wire \ces_5_4_io_ins_down[22] ;
 wire \ces_5_4_io_ins_down[23] ;
 wire \ces_5_4_io_ins_down[24] ;
 wire \ces_5_4_io_ins_down[25] ;
 wire \ces_5_4_io_ins_down[26] ;
 wire \ces_5_4_io_ins_down[27] ;
 wire \ces_5_4_io_ins_down[28] ;
 wire \ces_5_4_io_ins_down[29] ;
 wire \ces_5_4_io_ins_down[2] ;
 wire \ces_5_4_io_ins_down[30] ;
 wire \ces_5_4_io_ins_down[31] ;
 wire \ces_5_4_io_ins_down[32] ;
 wire \ces_5_4_io_ins_down[33] ;
 wire \ces_5_4_io_ins_down[34] ;
 wire \ces_5_4_io_ins_down[35] ;
 wire \ces_5_4_io_ins_down[36] ;
 wire \ces_5_4_io_ins_down[37] ;
 wire \ces_5_4_io_ins_down[38] ;
 wire \ces_5_4_io_ins_down[39] ;
 wire \ces_5_4_io_ins_down[3] ;
 wire \ces_5_4_io_ins_down[40] ;
 wire \ces_5_4_io_ins_down[41] ;
 wire \ces_5_4_io_ins_down[42] ;
 wire \ces_5_4_io_ins_down[43] ;
 wire \ces_5_4_io_ins_down[44] ;
 wire \ces_5_4_io_ins_down[45] ;
 wire \ces_5_4_io_ins_down[46] ;
 wire \ces_5_4_io_ins_down[47] ;
 wire \ces_5_4_io_ins_down[48] ;
 wire \ces_5_4_io_ins_down[49] ;
 wire \ces_5_4_io_ins_down[4] ;
 wire \ces_5_4_io_ins_down[50] ;
 wire \ces_5_4_io_ins_down[51] ;
 wire \ces_5_4_io_ins_down[52] ;
 wire \ces_5_4_io_ins_down[53] ;
 wire \ces_5_4_io_ins_down[54] ;
 wire \ces_5_4_io_ins_down[55] ;
 wire \ces_5_4_io_ins_down[56] ;
 wire \ces_5_4_io_ins_down[57] ;
 wire \ces_5_4_io_ins_down[58] ;
 wire \ces_5_4_io_ins_down[59] ;
 wire \ces_5_4_io_ins_down[5] ;
 wire \ces_5_4_io_ins_down[60] ;
 wire \ces_5_4_io_ins_down[61] ;
 wire \ces_5_4_io_ins_down[62] ;
 wire \ces_5_4_io_ins_down[63] ;
 wire \ces_5_4_io_ins_down[6] ;
 wire \ces_5_4_io_ins_down[7] ;
 wire \ces_5_4_io_ins_down[8] ;
 wire \ces_5_4_io_ins_down[9] ;
 wire \ces_5_4_io_ins_left[0] ;
 wire \ces_5_4_io_ins_left[10] ;
 wire \ces_5_4_io_ins_left[11] ;
 wire \ces_5_4_io_ins_left[12] ;
 wire \ces_5_4_io_ins_left[13] ;
 wire \ces_5_4_io_ins_left[14] ;
 wire \ces_5_4_io_ins_left[15] ;
 wire \ces_5_4_io_ins_left[16] ;
 wire \ces_5_4_io_ins_left[17] ;
 wire \ces_5_4_io_ins_left[18] ;
 wire \ces_5_4_io_ins_left[19] ;
 wire \ces_5_4_io_ins_left[1] ;
 wire \ces_5_4_io_ins_left[20] ;
 wire \ces_5_4_io_ins_left[21] ;
 wire \ces_5_4_io_ins_left[22] ;
 wire \ces_5_4_io_ins_left[23] ;
 wire \ces_5_4_io_ins_left[24] ;
 wire \ces_5_4_io_ins_left[25] ;
 wire \ces_5_4_io_ins_left[26] ;
 wire \ces_5_4_io_ins_left[27] ;
 wire \ces_5_4_io_ins_left[28] ;
 wire \ces_5_4_io_ins_left[29] ;
 wire \ces_5_4_io_ins_left[2] ;
 wire \ces_5_4_io_ins_left[30] ;
 wire \ces_5_4_io_ins_left[31] ;
 wire \ces_5_4_io_ins_left[32] ;
 wire \ces_5_4_io_ins_left[33] ;
 wire \ces_5_4_io_ins_left[34] ;
 wire \ces_5_4_io_ins_left[35] ;
 wire \ces_5_4_io_ins_left[36] ;
 wire \ces_5_4_io_ins_left[37] ;
 wire \ces_5_4_io_ins_left[38] ;
 wire \ces_5_4_io_ins_left[39] ;
 wire \ces_5_4_io_ins_left[3] ;
 wire \ces_5_4_io_ins_left[40] ;
 wire \ces_5_4_io_ins_left[41] ;
 wire \ces_5_4_io_ins_left[42] ;
 wire \ces_5_4_io_ins_left[43] ;
 wire \ces_5_4_io_ins_left[44] ;
 wire \ces_5_4_io_ins_left[45] ;
 wire \ces_5_4_io_ins_left[46] ;
 wire \ces_5_4_io_ins_left[47] ;
 wire \ces_5_4_io_ins_left[48] ;
 wire \ces_5_4_io_ins_left[49] ;
 wire \ces_5_4_io_ins_left[4] ;
 wire \ces_5_4_io_ins_left[50] ;
 wire \ces_5_4_io_ins_left[51] ;
 wire \ces_5_4_io_ins_left[52] ;
 wire \ces_5_4_io_ins_left[53] ;
 wire \ces_5_4_io_ins_left[54] ;
 wire \ces_5_4_io_ins_left[55] ;
 wire \ces_5_4_io_ins_left[56] ;
 wire \ces_5_4_io_ins_left[57] ;
 wire \ces_5_4_io_ins_left[58] ;
 wire \ces_5_4_io_ins_left[59] ;
 wire \ces_5_4_io_ins_left[5] ;
 wire \ces_5_4_io_ins_left[60] ;
 wire \ces_5_4_io_ins_left[61] ;
 wire \ces_5_4_io_ins_left[62] ;
 wire \ces_5_4_io_ins_left[63] ;
 wire \ces_5_4_io_ins_left[6] ;
 wire \ces_5_4_io_ins_left[7] ;
 wire \ces_5_4_io_ins_left[8] ;
 wire \ces_5_4_io_ins_left[9] ;
 wire ces_5_4_io_lsbOuts_0;
 wire ces_5_4_io_lsbOuts_1;
 wire ces_5_4_io_lsbOuts_2;
 wire ces_5_4_io_lsbOuts_3;
 wire ces_5_4_io_lsbOuts_4;
 wire ces_5_4_io_lsbOuts_5;
 wire ces_5_4_io_lsbOuts_6;
 wire ces_5_4_io_lsbOuts_7;
 wire \ces_5_4_io_outs_right[0] ;
 wire \ces_5_4_io_outs_right[10] ;
 wire \ces_5_4_io_outs_right[11] ;
 wire \ces_5_4_io_outs_right[12] ;
 wire \ces_5_4_io_outs_right[13] ;
 wire \ces_5_4_io_outs_right[14] ;
 wire \ces_5_4_io_outs_right[15] ;
 wire \ces_5_4_io_outs_right[16] ;
 wire \ces_5_4_io_outs_right[17] ;
 wire \ces_5_4_io_outs_right[18] ;
 wire \ces_5_4_io_outs_right[19] ;
 wire \ces_5_4_io_outs_right[1] ;
 wire \ces_5_4_io_outs_right[20] ;
 wire \ces_5_4_io_outs_right[21] ;
 wire \ces_5_4_io_outs_right[22] ;
 wire \ces_5_4_io_outs_right[23] ;
 wire \ces_5_4_io_outs_right[24] ;
 wire \ces_5_4_io_outs_right[25] ;
 wire \ces_5_4_io_outs_right[26] ;
 wire \ces_5_4_io_outs_right[27] ;
 wire \ces_5_4_io_outs_right[28] ;
 wire \ces_5_4_io_outs_right[29] ;
 wire \ces_5_4_io_outs_right[2] ;
 wire \ces_5_4_io_outs_right[30] ;
 wire \ces_5_4_io_outs_right[31] ;
 wire \ces_5_4_io_outs_right[32] ;
 wire \ces_5_4_io_outs_right[33] ;
 wire \ces_5_4_io_outs_right[34] ;
 wire \ces_5_4_io_outs_right[35] ;
 wire \ces_5_4_io_outs_right[36] ;
 wire \ces_5_4_io_outs_right[37] ;
 wire \ces_5_4_io_outs_right[38] ;
 wire \ces_5_4_io_outs_right[39] ;
 wire \ces_5_4_io_outs_right[3] ;
 wire \ces_5_4_io_outs_right[40] ;
 wire \ces_5_4_io_outs_right[41] ;
 wire \ces_5_4_io_outs_right[42] ;
 wire \ces_5_4_io_outs_right[43] ;
 wire \ces_5_4_io_outs_right[44] ;
 wire \ces_5_4_io_outs_right[45] ;
 wire \ces_5_4_io_outs_right[46] ;
 wire \ces_5_4_io_outs_right[47] ;
 wire \ces_5_4_io_outs_right[48] ;
 wire \ces_5_4_io_outs_right[49] ;
 wire \ces_5_4_io_outs_right[4] ;
 wire \ces_5_4_io_outs_right[50] ;
 wire \ces_5_4_io_outs_right[51] ;
 wire \ces_5_4_io_outs_right[52] ;
 wire \ces_5_4_io_outs_right[53] ;
 wire \ces_5_4_io_outs_right[54] ;
 wire \ces_5_4_io_outs_right[55] ;
 wire \ces_5_4_io_outs_right[56] ;
 wire \ces_5_4_io_outs_right[57] ;
 wire \ces_5_4_io_outs_right[58] ;
 wire \ces_5_4_io_outs_right[59] ;
 wire \ces_5_4_io_outs_right[5] ;
 wire \ces_5_4_io_outs_right[60] ;
 wire \ces_5_4_io_outs_right[61] ;
 wire \ces_5_4_io_outs_right[62] ;
 wire \ces_5_4_io_outs_right[63] ;
 wire \ces_5_4_io_outs_right[6] ;
 wire \ces_5_4_io_outs_right[7] ;
 wire \ces_5_4_io_outs_right[8] ;
 wire \ces_5_4_io_outs_right[9] ;
 wire \ces_5_4_io_outs_up[0] ;
 wire \ces_5_4_io_outs_up[10] ;
 wire \ces_5_4_io_outs_up[11] ;
 wire \ces_5_4_io_outs_up[12] ;
 wire \ces_5_4_io_outs_up[13] ;
 wire \ces_5_4_io_outs_up[14] ;
 wire \ces_5_4_io_outs_up[15] ;
 wire \ces_5_4_io_outs_up[16] ;
 wire \ces_5_4_io_outs_up[17] ;
 wire \ces_5_4_io_outs_up[18] ;
 wire \ces_5_4_io_outs_up[19] ;
 wire \ces_5_4_io_outs_up[1] ;
 wire \ces_5_4_io_outs_up[20] ;
 wire \ces_5_4_io_outs_up[21] ;
 wire \ces_5_4_io_outs_up[22] ;
 wire \ces_5_4_io_outs_up[23] ;
 wire \ces_5_4_io_outs_up[24] ;
 wire \ces_5_4_io_outs_up[25] ;
 wire \ces_5_4_io_outs_up[26] ;
 wire \ces_5_4_io_outs_up[27] ;
 wire \ces_5_4_io_outs_up[28] ;
 wire \ces_5_4_io_outs_up[29] ;
 wire \ces_5_4_io_outs_up[2] ;
 wire \ces_5_4_io_outs_up[30] ;
 wire \ces_5_4_io_outs_up[31] ;
 wire \ces_5_4_io_outs_up[32] ;
 wire \ces_5_4_io_outs_up[33] ;
 wire \ces_5_4_io_outs_up[34] ;
 wire \ces_5_4_io_outs_up[35] ;
 wire \ces_5_4_io_outs_up[36] ;
 wire \ces_5_4_io_outs_up[37] ;
 wire \ces_5_4_io_outs_up[38] ;
 wire \ces_5_4_io_outs_up[39] ;
 wire \ces_5_4_io_outs_up[3] ;
 wire \ces_5_4_io_outs_up[40] ;
 wire \ces_5_4_io_outs_up[41] ;
 wire \ces_5_4_io_outs_up[42] ;
 wire \ces_5_4_io_outs_up[43] ;
 wire \ces_5_4_io_outs_up[44] ;
 wire \ces_5_4_io_outs_up[45] ;
 wire \ces_5_4_io_outs_up[46] ;
 wire \ces_5_4_io_outs_up[47] ;
 wire \ces_5_4_io_outs_up[48] ;
 wire \ces_5_4_io_outs_up[49] ;
 wire \ces_5_4_io_outs_up[4] ;
 wire \ces_5_4_io_outs_up[50] ;
 wire \ces_5_4_io_outs_up[51] ;
 wire \ces_5_4_io_outs_up[52] ;
 wire \ces_5_4_io_outs_up[53] ;
 wire \ces_5_4_io_outs_up[54] ;
 wire \ces_5_4_io_outs_up[55] ;
 wire \ces_5_4_io_outs_up[56] ;
 wire \ces_5_4_io_outs_up[57] ;
 wire \ces_5_4_io_outs_up[58] ;
 wire \ces_5_4_io_outs_up[59] ;
 wire \ces_5_4_io_outs_up[5] ;
 wire \ces_5_4_io_outs_up[60] ;
 wire \ces_5_4_io_outs_up[61] ;
 wire \ces_5_4_io_outs_up[62] ;
 wire \ces_5_4_io_outs_up[63] ;
 wire \ces_5_4_io_outs_up[6] ;
 wire \ces_5_4_io_outs_up[7] ;
 wire \ces_5_4_io_outs_up[8] ;
 wire \ces_5_4_io_outs_up[9] ;
 wire \ces_5_5_io_ins_down[0] ;
 wire \ces_5_5_io_ins_down[10] ;
 wire \ces_5_5_io_ins_down[11] ;
 wire \ces_5_5_io_ins_down[12] ;
 wire \ces_5_5_io_ins_down[13] ;
 wire \ces_5_5_io_ins_down[14] ;
 wire \ces_5_5_io_ins_down[15] ;
 wire \ces_5_5_io_ins_down[16] ;
 wire \ces_5_5_io_ins_down[17] ;
 wire \ces_5_5_io_ins_down[18] ;
 wire \ces_5_5_io_ins_down[19] ;
 wire \ces_5_5_io_ins_down[1] ;
 wire \ces_5_5_io_ins_down[20] ;
 wire \ces_5_5_io_ins_down[21] ;
 wire \ces_5_5_io_ins_down[22] ;
 wire \ces_5_5_io_ins_down[23] ;
 wire \ces_5_5_io_ins_down[24] ;
 wire \ces_5_5_io_ins_down[25] ;
 wire \ces_5_5_io_ins_down[26] ;
 wire \ces_5_5_io_ins_down[27] ;
 wire \ces_5_5_io_ins_down[28] ;
 wire \ces_5_5_io_ins_down[29] ;
 wire \ces_5_5_io_ins_down[2] ;
 wire \ces_5_5_io_ins_down[30] ;
 wire \ces_5_5_io_ins_down[31] ;
 wire \ces_5_5_io_ins_down[32] ;
 wire \ces_5_5_io_ins_down[33] ;
 wire \ces_5_5_io_ins_down[34] ;
 wire \ces_5_5_io_ins_down[35] ;
 wire \ces_5_5_io_ins_down[36] ;
 wire \ces_5_5_io_ins_down[37] ;
 wire \ces_5_5_io_ins_down[38] ;
 wire \ces_5_5_io_ins_down[39] ;
 wire \ces_5_5_io_ins_down[3] ;
 wire \ces_5_5_io_ins_down[40] ;
 wire \ces_5_5_io_ins_down[41] ;
 wire \ces_5_5_io_ins_down[42] ;
 wire \ces_5_5_io_ins_down[43] ;
 wire \ces_5_5_io_ins_down[44] ;
 wire \ces_5_5_io_ins_down[45] ;
 wire \ces_5_5_io_ins_down[46] ;
 wire \ces_5_5_io_ins_down[47] ;
 wire \ces_5_5_io_ins_down[48] ;
 wire \ces_5_5_io_ins_down[49] ;
 wire \ces_5_5_io_ins_down[4] ;
 wire \ces_5_5_io_ins_down[50] ;
 wire \ces_5_5_io_ins_down[51] ;
 wire \ces_5_5_io_ins_down[52] ;
 wire \ces_5_5_io_ins_down[53] ;
 wire \ces_5_5_io_ins_down[54] ;
 wire \ces_5_5_io_ins_down[55] ;
 wire \ces_5_5_io_ins_down[56] ;
 wire \ces_5_5_io_ins_down[57] ;
 wire \ces_5_5_io_ins_down[58] ;
 wire \ces_5_5_io_ins_down[59] ;
 wire \ces_5_5_io_ins_down[5] ;
 wire \ces_5_5_io_ins_down[60] ;
 wire \ces_5_5_io_ins_down[61] ;
 wire \ces_5_5_io_ins_down[62] ;
 wire \ces_5_5_io_ins_down[63] ;
 wire \ces_5_5_io_ins_down[6] ;
 wire \ces_5_5_io_ins_down[7] ;
 wire \ces_5_5_io_ins_down[8] ;
 wire \ces_5_5_io_ins_down[9] ;
 wire \ces_5_5_io_ins_left[0] ;
 wire \ces_5_5_io_ins_left[10] ;
 wire \ces_5_5_io_ins_left[11] ;
 wire \ces_5_5_io_ins_left[12] ;
 wire \ces_5_5_io_ins_left[13] ;
 wire \ces_5_5_io_ins_left[14] ;
 wire \ces_5_5_io_ins_left[15] ;
 wire \ces_5_5_io_ins_left[16] ;
 wire \ces_5_5_io_ins_left[17] ;
 wire \ces_5_5_io_ins_left[18] ;
 wire \ces_5_5_io_ins_left[19] ;
 wire \ces_5_5_io_ins_left[1] ;
 wire \ces_5_5_io_ins_left[20] ;
 wire \ces_5_5_io_ins_left[21] ;
 wire \ces_5_5_io_ins_left[22] ;
 wire \ces_5_5_io_ins_left[23] ;
 wire \ces_5_5_io_ins_left[24] ;
 wire \ces_5_5_io_ins_left[25] ;
 wire \ces_5_5_io_ins_left[26] ;
 wire \ces_5_5_io_ins_left[27] ;
 wire \ces_5_5_io_ins_left[28] ;
 wire \ces_5_5_io_ins_left[29] ;
 wire \ces_5_5_io_ins_left[2] ;
 wire \ces_5_5_io_ins_left[30] ;
 wire \ces_5_5_io_ins_left[31] ;
 wire \ces_5_5_io_ins_left[32] ;
 wire \ces_5_5_io_ins_left[33] ;
 wire \ces_5_5_io_ins_left[34] ;
 wire \ces_5_5_io_ins_left[35] ;
 wire \ces_5_5_io_ins_left[36] ;
 wire \ces_5_5_io_ins_left[37] ;
 wire \ces_5_5_io_ins_left[38] ;
 wire \ces_5_5_io_ins_left[39] ;
 wire \ces_5_5_io_ins_left[3] ;
 wire \ces_5_5_io_ins_left[40] ;
 wire \ces_5_5_io_ins_left[41] ;
 wire \ces_5_5_io_ins_left[42] ;
 wire \ces_5_5_io_ins_left[43] ;
 wire \ces_5_5_io_ins_left[44] ;
 wire \ces_5_5_io_ins_left[45] ;
 wire \ces_5_5_io_ins_left[46] ;
 wire \ces_5_5_io_ins_left[47] ;
 wire \ces_5_5_io_ins_left[48] ;
 wire \ces_5_5_io_ins_left[49] ;
 wire \ces_5_5_io_ins_left[4] ;
 wire \ces_5_5_io_ins_left[50] ;
 wire \ces_5_5_io_ins_left[51] ;
 wire \ces_5_5_io_ins_left[52] ;
 wire \ces_5_5_io_ins_left[53] ;
 wire \ces_5_5_io_ins_left[54] ;
 wire \ces_5_5_io_ins_left[55] ;
 wire \ces_5_5_io_ins_left[56] ;
 wire \ces_5_5_io_ins_left[57] ;
 wire \ces_5_5_io_ins_left[58] ;
 wire \ces_5_5_io_ins_left[59] ;
 wire \ces_5_5_io_ins_left[5] ;
 wire \ces_5_5_io_ins_left[60] ;
 wire \ces_5_5_io_ins_left[61] ;
 wire \ces_5_5_io_ins_left[62] ;
 wire \ces_5_5_io_ins_left[63] ;
 wire \ces_5_5_io_ins_left[6] ;
 wire \ces_5_5_io_ins_left[7] ;
 wire \ces_5_5_io_ins_left[8] ;
 wire \ces_5_5_io_ins_left[9] ;
 wire ces_5_5_io_lsbOuts_0;
 wire ces_5_5_io_lsbOuts_1;
 wire ces_5_5_io_lsbOuts_2;
 wire ces_5_5_io_lsbOuts_3;
 wire ces_5_5_io_lsbOuts_4;
 wire ces_5_5_io_lsbOuts_5;
 wire ces_5_5_io_lsbOuts_6;
 wire ces_5_5_io_lsbOuts_7;
 wire \ces_5_5_io_outs_right[0] ;
 wire \ces_5_5_io_outs_right[10] ;
 wire \ces_5_5_io_outs_right[11] ;
 wire \ces_5_5_io_outs_right[12] ;
 wire \ces_5_5_io_outs_right[13] ;
 wire \ces_5_5_io_outs_right[14] ;
 wire \ces_5_5_io_outs_right[15] ;
 wire \ces_5_5_io_outs_right[16] ;
 wire \ces_5_5_io_outs_right[17] ;
 wire \ces_5_5_io_outs_right[18] ;
 wire \ces_5_5_io_outs_right[19] ;
 wire \ces_5_5_io_outs_right[1] ;
 wire \ces_5_5_io_outs_right[20] ;
 wire \ces_5_5_io_outs_right[21] ;
 wire \ces_5_5_io_outs_right[22] ;
 wire \ces_5_5_io_outs_right[23] ;
 wire \ces_5_5_io_outs_right[24] ;
 wire \ces_5_5_io_outs_right[25] ;
 wire \ces_5_5_io_outs_right[26] ;
 wire \ces_5_5_io_outs_right[27] ;
 wire \ces_5_5_io_outs_right[28] ;
 wire \ces_5_5_io_outs_right[29] ;
 wire \ces_5_5_io_outs_right[2] ;
 wire \ces_5_5_io_outs_right[30] ;
 wire \ces_5_5_io_outs_right[31] ;
 wire \ces_5_5_io_outs_right[32] ;
 wire \ces_5_5_io_outs_right[33] ;
 wire \ces_5_5_io_outs_right[34] ;
 wire \ces_5_5_io_outs_right[35] ;
 wire \ces_5_5_io_outs_right[36] ;
 wire \ces_5_5_io_outs_right[37] ;
 wire \ces_5_5_io_outs_right[38] ;
 wire \ces_5_5_io_outs_right[39] ;
 wire \ces_5_5_io_outs_right[3] ;
 wire \ces_5_5_io_outs_right[40] ;
 wire \ces_5_5_io_outs_right[41] ;
 wire \ces_5_5_io_outs_right[42] ;
 wire \ces_5_5_io_outs_right[43] ;
 wire \ces_5_5_io_outs_right[44] ;
 wire \ces_5_5_io_outs_right[45] ;
 wire \ces_5_5_io_outs_right[46] ;
 wire \ces_5_5_io_outs_right[47] ;
 wire \ces_5_5_io_outs_right[48] ;
 wire \ces_5_5_io_outs_right[49] ;
 wire \ces_5_5_io_outs_right[4] ;
 wire \ces_5_5_io_outs_right[50] ;
 wire \ces_5_5_io_outs_right[51] ;
 wire \ces_5_5_io_outs_right[52] ;
 wire \ces_5_5_io_outs_right[53] ;
 wire \ces_5_5_io_outs_right[54] ;
 wire \ces_5_5_io_outs_right[55] ;
 wire \ces_5_5_io_outs_right[56] ;
 wire \ces_5_5_io_outs_right[57] ;
 wire \ces_5_5_io_outs_right[58] ;
 wire \ces_5_5_io_outs_right[59] ;
 wire \ces_5_5_io_outs_right[5] ;
 wire \ces_5_5_io_outs_right[60] ;
 wire \ces_5_5_io_outs_right[61] ;
 wire \ces_5_5_io_outs_right[62] ;
 wire \ces_5_5_io_outs_right[63] ;
 wire \ces_5_5_io_outs_right[6] ;
 wire \ces_5_5_io_outs_right[7] ;
 wire \ces_5_5_io_outs_right[8] ;
 wire \ces_5_5_io_outs_right[9] ;
 wire \ces_5_5_io_outs_up[0] ;
 wire \ces_5_5_io_outs_up[10] ;
 wire \ces_5_5_io_outs_up[11] ;
 wire \ces_5_5_io_outs_up[12] ;
 wire \ces_5_5_io_outs_up[13] ;
 wire \ces_5_5_io_outs_up[14] ;
 wire \ces_5_5_io_outs_up[15] ;
 wire \ces_5_5_io_outs_up[16] ;
 wire \ces_5_5_io_outs_up[17] ;
 wire \ces_5_5_io_outs_up[18] ;
 wire \ces_5_5_io_outs_up[19] ;
 wire \ces_5_5_io_outs_up[1] ;
 wire \ces_5_5_io_outs_up[20] ;
 wire \ces_5_5_io_outs_up[21] ;
 wire \ces_5_5_io_outs_up[22] ;
 wire \ces_5_5_io_outs_up[23] ;
 wire \ces_5_5_io_outs_up[24] ;
 wire \ces_5_5_io_outs_up[25] ;
 wire \ces_5_5_io_outs_up[26] ;
 wire \ces_5_5_io_outs_up[27] ;
 wire \ces_5_5_io_outs_up[28] ;
 wire \ces_5_5_io_outs_up[29] ;
 wire \ces_5_5_io_outs_up[2] ;
 wire \ces_5_5_io_outs_up[30] ;
 wire \ces_5_5_io_outs_up[31] ;
 wire \ces_5_5_io_outs_up[32] ;
 wire \ces_5_5_io_outs_up[33] ;
 wire \ces_5_5_io_outs_up[34] ;
 wire \ces_5_5_io_outs_up[35] ;
 wire \ces_5_5_io_outs_up[36] ;
 wire \ces_5_5_io_outs_up[37] ;
 wire \ces_5_5_io_outs_up[38] ;
 wire \ces_5_5_io_outs_up[39] ;
 wire \ces_5_5_io_outs_up[3] ;
 wire \ces_5_5_io_outs_up[40] ;
 wire \ces_5_5_io_outs_up[41] ;
 wire \ces_5_5_io_outs_up[42] ;
 wire \ces_5_5_io_outs_up[43] ;
 wire \ces_5_5_io_outs_up[44] ;
 wire \ces_5_5_io_outs_up[45] ;
 wire \ces_5_5_io_outs_up[46] ;
 wire \ces_5_5_io_outs_up[47] ;
 wire \ces_5_5_io_outs_up[48] ;
 wire \ces_5_5_io_outs_up[49] ;
 wire \ces_5_5_io_outs_up[4] ;
 wire \ces_5_5_io_outs_up[50] ;
 wire \ces_5_5_io_outs_up[51] ;
 wire \ces_5_5_io_outs_up[52] ;
 wire \ces_5_5_io_outs_up[53] ;
 wire \ces_5_5_io_outs_up[54] ;
 wire \ces_5_5_io_outs_up[55] ;
 wire \ces_5_5_io_outs_up[56] ;
 wire \ces_5_5_io_outs_up[57] ;
 wire \ces_5_5_io_outs_up[58] ;
 wire \ces_5_5_io_outs_up[59] ;
 wire \ces_5_5_io_outs_up[5] ;
 wire \ces_5_5_io_outs_up[60] ;
 wire \ces_5_5_io_outs_up[61] ;
 wire \ces_5_5_io_outs_up[62] ;
 wire \ces_5_5_io_outs_up[63] ;
 wire \ces_5_5_io_outs_up[6] ;
 wire \ces_5_5_io_outs_up[7] ;
 wire \ces_5_5_io_outs_up[8] ;
 wire \ces_5_5_io_outs_up[9] ;
 wire \ces_5_6_io_ins_down[0] ;
 wire \ces_5_6_io_ins_down[10] ;
 wire \ces_5_6_io_ins_down[11] ;
 wire \ces_5_6_io_ins_down[12] ;
 wire \ces_5_6_io_ins_down[13] ;
 wire \ces_5_6_io_ins_down[14] ;
 wire \ces_5_6_io_ins_down[15] ;
 wire \ces_5_6_io_ins_down[16] ;
 wire \ces_5_6_io_ins_down[17] ;
 wire \ces_5_6_io_ins_down[18] ;
 wire \ces_5_6_io_ins_down[19] ;
 wire \ces_5_6_io_ins_down[1] ;
 wire \ces_5_6_io_ins_down[20] ;
 wire \ces_5_6_io_ins_down[21] ;
 wire \ces_5_6_io_ins_down[22] ;
 wire \ces_5_6_io_ins_down[23] ;
 wire \ces_5_6_io_ins_down[24] ;
 wire \ces_5_6_io_ins_down[25] ;
 wire \ces_5_6_io_ins_down[26] ;
 wire \ces_5_6_io_ins_down[27] ;
 wire \ces_5_6_io_ins_down[28] ;
 wire \ces_5_6_io_ins_down[29] ;
 wire \ces_5_6_io_ins_down[2] ;
 wire \ces_5_6_io_ins_down[30] ;
 wire \ces_5_6_io_ins_down[31] ;
 wire \ces_5_6_io_ins_down[32] ;
 wire \ces_5_6_io_ins_down[33] ;
 wire \ces_5_6_io_ins_down[34] ;
 wire \ces_5_6_io_ins_down[35] ;
 wire \ces_5_6_io_ins_down[36] ;
 wire \ces_5_6_io_ins_down[37] ;
 wire \ces_5_6_io_ins_down[38] ;
 wire \ces_5_6_io_ins_down[39] ;
 wire \ces_5_6_io_ins_down[3] ;
 wire \ces_5_6_io_ins_down[40] ;
 wire \ces_5_6_io_ins_down[41] ;
 wire \ces_5_6_io_ins_down[42] ;
 wire \ces_5_6_io_ins_down[43] ;
 wire \ces_5_6_io_ins_down[44] ;
 wire \ces_5_6_io_ins_down[45] ;
 wire \ces_5_6_io_ins_down[46] ;
 wire \ces_5_6_io_ins_down[47] ;
 wire \ces_5_6_io_ins_down[48] ;
 wire \ces_5_6_io_ins_down[49] ;
 wire \ces_5_6_io_ins_down[4] ;
 wire \ces_5_6_io_ins_down[50] ;
 wire \ces_5_6_io_ins_down[51] ;
 wire \ces_5_6_io_ins_down[52] ;
 wire \ces_5_6_io_ins_down[53] ;
 wire \ces_5_6_io_ins_down[54] ;
 wire \ces_5_6_io_ins_down[55] ;
 wire \ces_5_6_io_ins_down[56] ;
 wire \ces_5_6_io_ins_down[57] ;
 wire \ces_5_6_io_ins_down[58] ;
 wire \ces_5_6_io_ins_down[59] ;
 wire \ces_5_6_io_ins_down[5] ;
 wire \ces_5_6_io_ins_down[60] ;
 wire \ces_5_6_io_ins_down[61] ;
 wire \ces_5_6_io_ins_down[62] ;
 wire \ces_5_6_io_ins_down[63] ;
 wire \ces_5_6_io_ins_down[6] ;
 wire \ces_5_6_io_ins_down[7] ;
 wire \ces_5_6_io_ins_down[8] ;
 wire \ces_5_6_io_ins_down[9] ;
 wire \ces_5_6_io_ins_left[0] ;
 wire \ces_5_6_io_ins_left[10] ;
 wire \ces_5_6_io_ins_left[11] ;
 wire \ces_5_6_io_ins_left[12] ;
 wire \ces_5_6_io_ins_left[13] ;
 wire \ces_5_6_io_ins_left[14] ;
 wire \ces_5_6_io_ins_left[15] ;
 wire \ces_5_6_io_ins_left[16] ;
 wire \ces_5_6_io_ins_left[17] ;
 wire \ces_5_6_io_ins_left[18] ;
 wire \ces_5_6_io_ins_left[19] ;
 wire \ces_5_6_io_ins_left[1] ;
 wire \ces_5_6_io_ins_left[20] ;
 wire \ces_5_6_io_ins_left[21] ;
 wire \ces_5_6_io_ins_left[22] ;
 wire \ces_5_6_io_ins_left[23] ;
 wire \ces_5_6_io_ins_left[24] ;
 wire \ces_5_6_io_ins_left[25] ;
 wire \ces_5_6_io_ins_left[26] ;
 wire \ces_5_6_io_ins_left[27] ;
 wire \ces_5_6_io_ins_left[28] ;
 wire \ces_5_6_io_ins_left[29] ;
 wire \ces_5_6_io_ins_left[2] ;
 wire \ces_5_6_io_ins_left[30] ;
 wire \ces_5_6_io_ins_left[31] ;
 wire \ces_5_6_io_ins_left[32] ;
 wire \ces_5_6_io_ins_left[33] ;
 wire \ces_5_6_io_ins_left[34] ;
 wire \ces_5_6_io_ins_left[35] ;
 wire \ces_5_6_io_ins_left[36] ;
 wire \ces_5_6_io_ins_left[37] ;
 wire \ces_5_6_io_ins_left[38] ;
 wire \ces_5_6_io_ins_left[39] ;
 wire \ces_5_6_io_ins_left[3] ;
 wire \ces_5_6_io_ins_left[40] ;
 wire \ces_5_6_io_ins_left[41] ;
 wire \ces_5_6_io_ins_left[42] ;
 wire \ces_5_6_io_ins_left[43] ;
 wire \ces_5_6_io_ins_left[44] ;
 wire \ces_5_6_io_ins_left[45] ;
 wire \ces_5_6_io_ins_left[46] ;
 wire \ces_5_6_io_ins_left[47] ;
 wire \ces_5_6_io_ins_left[48] ;
 wire \ces_5_6_io_ins_left[49] ;
 wire \ces_5_6_io_ins_left[4] ;
 wire \ces_5_6_io_ins_left[50] ;
 wire \ces_5_6_io_ins_left[51] ;
 wire \ces_5_6_io_ins_left[52] ;
 wire \ces_5_6_io_ins_left[53] ;
 wire \ces_5_6_io_ins_left[54] ;
 wire \ces_5_6_io_ins_left[55] ;
 wire \ces_5_6_io_ins_left[56] ;
 wire \ces_5_6_io_ins_left[57] ;
 wire \ces_5_6_io_ins_left[58] ;
 wire \ces_5_6_io_ins_left[59] ;
 wire \ces_5_6_io_ins_left[5] ;
 wire \ces_5_6_io_ins_left[60] ;
 wire \ces_5_6_io_ins_left[61] ;
 wire \ces_5_6_io_ins_left[62] ;
 wire \ces_5_6_io_ins_left[63] ;
 wire \ces_5_6_io_ins_left[6] ;
 wire \ces_5_6_io_ins_left[7] ;
 wire \ces_5_6_io_ins_left[8] ;
 wire \ces_5_6_io_ins_left[9] ;
 wire ces_5_6_io_lsbOuts_0;
 wire ces_5_6_io_lsbOuts_1;
 wire ces_5_6_io_lsbOuts_2;
 wire ces_5_6_io_lsbOuts_3;
 wire ces_5_6_io_lsbOuts_4;
 wire ces_5_6_io_lsbOuts_5;
 wire ces_5_6_io_lsbOuts_6;
 wire ces_5_6_io_lsbOuts_7;
 wire \ces_5_6_io_outs_right[0] ;
 wire \ces_5_6_io_outs_right[10] ;
 wire \ces_5_6_io_outs_right[11] ;
 wire \ces_5_6_io_outs_right[12] ;
 wire \ces_5_6_io_outs_right[13] ;
 wire \ces_5_6_io_outs_right[14] ;
 wire \ces_5_6_io_outs_right[15] ;
 wire \ces_5_6_io_outs_right[16] ;
 wire \ces_5_6_io_outs_right[17] ;
 wire \ces_5_6_io_outs_right[18] ;
 wire \ces_5_6_io_outs_right[19] ;
 wire \ces_5_6_io_outs_right[1] ;
 wire \ces_5_6_io_outs_right[20] ;
 wire \ces_5_6_io_outs_right[21] ;
 wire \ces_5_6_io_outs_right[22] ;
 wire \ces_5_6_io_outs_right[23] ;
 wire \ces_5_6_io_outs_right[24] ;
 wire \ces_5_6_io_outs_right[25] ;
 wire \ces_5_6_io_outs_right[26] ;
 wire \ces_5_6_io_outs_right[27] ;
 wire \ces_5_6_io_outs_right[28] ;
 wire \ces_5_6_io_outs_right[29] ;
 wire \ces_5_6_io_outs_right[2] ;
 wire \ces_5_6_io_outs_right[30] ;
 wire \ces_5_6_io_outs_right[31] ;
 wire \ces_5_6_io_outs_right[32] ;
 wire \ces_5_6_io_outs_right[33] ;
 wire \ces_5_6_io_outs_right[34] ;
 wire \ces_5_6_io_outs_right[35] ;
 wire \ces_5_6_io_outs_right[36] ;
 wire \ces_5_6_io_outs_right[37] ;
 wire \ces_5_6_io_outs_right[38] ;
 wire \ces_5_6_io_outs_right[39] ;
 wire \ces_5_6_io_outs_right[3] ;
 wire \ces_5_6_io_outs_right[40] ;
 wire \ces_5_6_io_outs_right[41] ;
 wire \ces_5_6_io_outs_right[42] ;
 wire \ces_5_6_io_outs_right[43] ;
 wire \ces_5_6_io_outs_right[44] ;
 wire \ces_5_6_io_outs_right[45] ;
 wire \ces_5_6_io_outs_right[46] ;
 wire \ces_5_6_io_outs_right[47] ;
 wire \ces_5_6_io_outs_right[48] ;
 wire \ces_5_6_io_outs_right[49] ;
 wire \ces_5_6_io_outs_right[4] ;
 wire \ces_5_6_io_outs_right[50] ;
 wire \ces_5_6_io_outs_right[51] ;
 wire \ces_5_6_io_outs_right[52] ;
 wire \ces_5_6_io_outs_right[53] ;
 wire \ces_5_6_io_outs_right[54] ;
 wire \ces_5_6_io_outs_right[55] ;
 wire \ces_5_6_io_outs_right[56] ;
 wire \ces_5_6_io_outs_right[57] ;
 wire \ces_5_6_io_outs_right[58] ;
 wire \ces_5_6_io_outs_right[59] ;
 wire \ces_5_6_io_outs_right[5] ;
 wire \ces_5_6_io_outs_right[60] ;
 wire \ces_5_6_io_outs_right[61] ;
 wire \ces_5_6_io_outs_right[62] ;
 wire \ces_5_6_io_outs_right[63] ;
 wire \ces_5_6_io_outs_right[6] ;
 wire \ces_5_6_io_outs_right[7] ;
 wire \ces_5_6_io_outs_right[8] ;
 wire \ces_5_6_io_outs_right[9] ;
 wire \ces_5_6_io_outs_up[0] ;
 wire \ces_5_6_io_outs_up[10] ;
 wire \ces_5_6_io_outs_up[11] ;
 wire \ces_5_6_io_outs_up[12] ;
 wire \ces_5_6_io_outs_up[13] ;
 wire \ces_5_6_io_outs_up[14] ;
 wire \ces_5_6_io_outs_up[15] ;
 wire \ces_5_6_io_outs_up[16] ;
 wire \ces_5_6_io_outs_up[17] ;
 wire \ces_5_6_io_outs_up[18] ;
 wire \ces_5_6_io_outs_up[19] ;
 wire \ces_5_6_io_outs_up[1] ;
 wire \ces_5_6_io_outs_up[20] ;
 wire \ces_5_6_io_outs_up[21] ;
 wire \ces_5_6_io_outs_up[22] ;
 wire \ces_5_6_io_outs_up[23] ;
 wire \ces_5_6_io_outs_up[24] ;
 wire \ces_5_6_io_outs_up[25] ;
 wire \ces_5_6_io_outs_up[26] ;
 wire \ces_5_6_io_outs_up[27] ;
 wire \ces_5_6_io_outs_up[28] ;
 wire \ces_5_6_io_outs_up[29] ;
 wire \ces_5_6_io_outs_up[2] ;
 wire \ces_5_6_io_outs_up[30] ;
 wire \ces_5_6_io_outs_up[31] ;
 wire \ces_5_6_io_outs_up[32] ;
 wire \ces_5_6_io_outs_up[33] ;
 wire \ces_5_6_io_outs_up[34] ;
 wire \ces_5_6_io_outs_up[35] ;
 wire \ces_5_6_io_outs_up[36] ;
 wire \ces_5_6_io_outs_up[37] ;
 wire \ces_5_6_io_outs_up[38] ;
 wire \ces_5_6_io_outs_up[39] ;
 wire \ces_5_6_io_outs_up[3] ;
 wire \ces_5_6_io_outs_up[40] ;
 wire \ces_5_6_io_outs_up[41] ;
 wire \ces_5_6_io_outs_up[42] ;
 wire \ces_5_6_io_outs_up[43] ;
 wire \ces_5_6_io_outs_up[44] ;
 wire \ces_5_6_io_outs_up[45] ;
 wire \ces_5_6_io_outs_up[46] ;
 wire \ces_5_6_io_outs_up[47] ;
 wire \ces_5_6_io_outs_up[48] ;
 wire \ces_5_6_io_outs_up[49] ;
 wire \ces_5_6_io_outs_up[4] ;
 wire \ces_5_6_io_outs_up[50] ;
 wire \ces_5_6_io_outs_up[51] ;
 wire \ces_5_6_io_outs_up[52] ;
 wire \ces_5_6_io_outs_up[53] ;
 wire \ces_5_6_io_outs_up[54] ;
 wire \ces_5_6_io_outs_up[55] ;
 wire \ces_5_6_io_outs_up[56] ;
 wire \ces_5_6_io_outs_up[57] ;
 wire \ces_5_6_io_outs_up[58] ;
 wire \ces_5_6_io_outs_up[59] ;
 wire \ces_5_6_io_outs_up[5] ;
 wire \ces_5_6_io_outs_up[60] ;
 wire \ces_5_6_io_outs_up[61] ;
 wire \ces_5_6_io_outs_up[62] ;
 wire \ces_5_6_io_outs_up[63] ;
 wire \ces_5_6_io_outs_up[6] ;
 wire \ces_5_6_io_outs_up[7] ;
 wire \ces_5_6_io_outs_up[8] ;
 wire \ces_5_6_io_outs_up[9] ;
 wire \ces_5_7_io_ins_down[0] ;
 wire \ces_5_7_io_ins_down[10] ;
 wire \ces_5_7_io_ins_down[11] ;
 wire \ces_5_7_io_ins_down[12] ;
 wire \ces_5_7_io_ins_down[13] ;
 wire \ces_5_7_io_ins_down[14] ;
 wire \ces_5_7_io_ins_down[15] ;
 wire \ces_5_7_io_ins_down[16] ;
 wire \ces_5_7_io_ins_down[17] ;
 wire \ces_5_7_io_ins_down[18] ;
 wire \ces_5_7_io_ins_down[19] ;
 wire \ces_5_7_io_ins_down[1] ;
 wire \ces_5_7_io_ins_down[20] ;
 wire \ces_5_7_io_ins_down[21] ;
 wire \ces_5_7_io_ins_down[22] ;
 wire \ces_5_7_io_ins_down[23] ;
 wire \ces_5_7_io_ins_down[24] ;
 wire \ces_5_7_io_ins_down[25] ;
 wire \ces_5_7_io_ins_down[26] ;
 wire \ces_5_7_io_ins_down[27] ;
 wire \ces_5_7_io_ins_down[28] ;
 wire \ces_5_7_io_ins_down[29] ;
 wire \ces_5_7_io_ins_down[2] ;
 wire \ces_5_7_io_ins_down[30] ;
 wire \ces_5_7_io_ins_down[31] ;
 wire \ces_5_7_io_ins_down[32] ;
 wire \ces_5_7_io_ins_down[33] ;
 wire \ces_5_7_io_ins_down[34] ;
 wire \ces_5_7_io_ins_down[35] ;
 wire \ces_5_7_io_ins_down[36] ;
 wire \ces_5_7_io_ins_down[37] ;
 wire \ces_5_7_io_ins_down[38] ;
 wire \ces_5_7_io_ins_down[39] ;
 wire \ces_5_7_io_ins_down[3] ;
 wire \ces_5_7_io_ins_down[40] ;
 wire \ces_5_7_io_ins_down[41] ;
 wire \ces_5_7_io_ins_down[42] ;
 wire \ces_5_7_io_ins_down[43] ;
 wire \ces_5_7_io_ins_down[44] ;
 wire \ces_5_7_io_ins_down[45] ;
 wire \ces_5_7_io_ins_down[46] ;
 wire \ces_5_7_io_ins_down[47] ;
 wire \ces_5_7_io_ins_down[48] ;
 wire \ces_5_7_io_ins_down[49] ;
 wire \ces_5_7_io_ins_down[4] ;
 wire \ces_5_7_io_ins_down[50] ;
 wire \ces_5_7_io_ins_down[51] ;
 wire \ces_5_7_io_ins_down[52] ;
 wire \ces_5_7_io_ins_down[53] ;
 wire \ces_5_7_io_ins_down[54] ;
 wire \ces_5_7_io_ins_down[55] ;
 wire \ces_5_7_io_ins_down[56] ;
 wire \ces_5_7_io_ins_down[57] ;
 wire \ces_5_7_io_ins_down[58] ;
 wire \ces_5_7_io_ins_down[59] ;
 wire \ces_5_7_io_ins_down[5] ;
 wire \ces_5_7_io_ins_down[60] ;
 wire \ces_5_7_io_ins_down[61] ;
 wire \ces_5_7_io_ins_down[62] ;
 wire \ces_5_7_io_ins_down[63] ;
 wire \ces_5_7_io_ins_down[6] ;
 wire \ces_5_7_io_ins_down[7] ;
 wire \ces_5_7_io_ins_down[8] ;
 wire \ces_5_7_io_ins_down[9] ;
 wire ces_5_7_io_lsbOuts_0;
 wire ces_5_7_io_lsbOuts_1;
 wire ces_5_7_io_lsbOuts_2;
 wire ces_5_7_io_lsbOuts_3;
 wire ces_5_7_io_lsbOuts_4;
 wire ces_5_7_io_lsbOuts_5;
 wire ces_5_7_io_lsbOuts_6;
 wire ces_5_7_io_lsbOuts_7;
 wire \ces_5_7_io_outs_up[0] ;
 wire \ces_5_7_io_outs_up[10] ;
 wire \ces_5_7_io_outs_up[11] ;
 wire \ces_5_7_io_outs_up[12] ;
 wire \ces_5_7_io_outs_up[13] ;
 wire \ces_5_7_io_outs_up[14] ;
 wire \ces_5_7_io_outs_up[15] ;
 wire \ces_5_7_io_outs_up[16] ;
 wire \ces_5_7_io_outs_up[17] ;
 wire \ces_5_7_io_outs_up[18] ;
 wire \ces_5_7_io_outs_up[19] ;
 wire \ces_5_7_io_outs_up[1] ;
 wire \ces_5_7_io_outs_up[20] ;
 wire \ces_5_7_io_outs_up[21] ;
 wire \ces_5_7_io_outs_up[22] ;
 wire \ces_5_7_io_outs_up[23] ;
 wire \ces_5_7_io_outs_up[24] ;
 wire \ces_5_7_io_outs_up[25] ;
 wire \ces_5_7_io_outs_up[26] ;
 wire \ces_5_7_io_outs_up[27] ;
 wire \ces_5_7_io_outs_up[28] ;
 wire \ces_5_7_io_outs_up[29] ;
 wire \ces_5_7_io_outs_up[2] ;
 wire \ces_5_7_io_outs_up[30] ;
 wire \ces_5_7_io_outs_up[31] ;
 wire \ces_5_7_io_outs_up[32] ;
 wire \ces_5_7_io_outs_up[33] ;
 wire \ces_5_7_io_outs_up[34] ;
 wire \ces_5_7_io_outs_up[35] ;
 wire \ces_5_7_io_outs_up[36] ;
 wire \ces_5_7_io_outs_up[37] ;
 wire \ces_5_7_io_outs_up[38] ;
 wire \ces_5_7_io_outs_up[39] ;
 wire \ces_5_7_io_outs_up[3] ;
 wire \ces_5_7_io_outs_up[40] ;
 wire \ces_5_7_io_outs_up[41] ;
 wire \ces_5_7_io_outs_up[42] ;
 wire \ces_5_7_io_outs_up[43] ;
 wire \ces_5_7_io_outs_up[44] ;
 wire \ces_5_7_io_outs_up[45] ;
 wire \ces_5_7_io_outs_up[46] ;
 wire \ces_5_7_io_outs_up[47] ;
 wire \ces_5_7_io_outs_up[48] ;
 wire \ces_5_7_io_outs_up[49] ;
 wire \ces_5_7_io_outs_up[4] ;
 wire \ces_5_7_io_outs_up[50] ;
 wire \ces_5_7_io_outs_up[51] ;
 wire \ces_5_7_io_outs_up[52] ;
 wire \ces_5_7_io_outs_up[53] ;
 wire \ces_5_7_io_outs_up[54] ;
 wire \ces_5_7_io_outs_up[55] ;
 wire \ces_5_7_io_outs_up[56] ;
 wire \ces_5_7_io_outs_up[57] ;
 wire \ces_5_7_io_outs_up[58] ;
 wire \ces_5_7_io_outs_up[59] ;
 wire \ces_5_7_io_outs_up[5] ;
 wire \ces_5_7_io_outs_up[60] ;
 wire \ces_5_7_io_outs_up[61] ;
 wire \ces_5_7_io_outs_up[62] ;
 wire \ces_5_7_io_outs_up[63] ;
 wire \ces_5_7_io_outs_up[6] ;
 wire \ces_5_7_io_outs_up[7] ;
 wire \ces_5_7_io_outs_up[8] ;
 wire \ces_5_7_io_outs_up[9] ;
 wire \ces_6_0_io_ins_down[0] ;
 wire \ces_6_0_io_ins_down[10] ;
 wire \ces_6_0_io_ins_down[11] ;
 wire \ces_6_0_io_ins_down[12] ;
 wire \ces_6_0_io_ins_down[13] ;
 wire \ces_6_0_io_ins_down[14] ;
 wire \ces_6_0_io_ins_down[15] ;
 wire \ces_6_0_io_ins_down[16] ;
 wire \ces_6_0_io_ins_down[17] ;
 wire \ces_6_0_io_ins_down[18] ;
 wire \ces_6_0_io_ins_down[19] ;
 wire \ces_6_0_io_ins_down[1] ;
 wire \ces_6_0_io_ins_down[20] ;
 wire \ces_6_0_io_ins_down[21] ;
 wire \ces_6_0_io_ins_down[22] ;
 wire \ces_6_0_io_ins_down[23] ;
 wire \ces_6_0_io_ins_down[24] ;
 wire \ces_6_0_io_ins_down[25] ;
 wire \ces_6_0_io_ins_down[26] ;
 wire \ces_6_0_io_ins_down[27] ;
 wire \ces_6_0_io_ins_down[28] ;
 wire \ces_6_0_io_ins_down[29] ;
 wire \ces_6_0_io_ins_down[2] ;
 wire \ces_6_0_io_ins_down[30] ;
 wire \ces_6_0_io_ins_down[31] ;
 wire \ces_6_0_io_ins_down[32] ;
 wire \ces_6_0_io_ins_down[33] ;
 wire \ces_6_0_io_ins_down[34] ;
 wire \ces_6_0_io_ins_down[35] ;
 wire \ces_6_0_io_ins_down[36] ;
 wire \ces_6_0_io_ins_down[37] ;
 wire \ces_6_0_io_ins_down[38] ;
 wire \ces_6_0_io_ins_down[39] ;
 wire \ces_6_0_io_ins_down[3] ;
 wire \ces_6_0_io_ins_down[40] ;
 wire \ces_6_0_io_ins_down[41] ;
 wire \ces_6_0_io_ins_down[42] ;
 wire \ces_6_0_io_ins_down[43] ;
 wire \ces_6_0_io_ins_down[44] ;
 wire \ces_6_0_io_ins_down[45] ;
 wire \ces_6_0_io_ins_down[46] ;
 wire \ces_6_0_io_ins_down[47] ;
 wire \ces_6_0_io_ins_down[48] ;
 wire \ces_6_0_io_ins_down[49] ;
 wire \ces_6_0_io_ins_down[4] ;
 wire \ces_6_0_io_ins_down[50] ;
 wire \ces_6_0_io_ins_down[51] ;
 wire \ces_6_0_io_ins_down[52] ;
 wire \ces_6_0_io_ins_down[53] ;
 wire \ces_6_0_io_ins_down[54] ;
 wire \ces_6_0_io_ins_down[55] ;
 wire \ces_6_0_io_ins_down[56] ;
 wire \ces_6_0_io_ins_down[57] ;
 wire \ces_6_0_io_ins_down[58] ;
 wire \ces_6_0_io_ins_down[59] ;
 wire \ces_6_0_io_ins_down[5] ;
 wire \ces_6_0_io_ins_down[60] ;
 wire \ces_6_0_io_ins_down[61] ;
 wire \ces_6_0_io_ins_down[62] ;
 wire \ces_6_0_io_ins_down[63] ;
 wire \ces_6_0_io_ins_down[6] ;
 wire \ces_6_0_io_ins_down[7] ;
 wire \ces_6_0_io_ins_down[8] ;
 wire \ces_6_0_io_ins_down[9] ;
 wire \ces_6_0_io_ins_left[0] ;
 wire \ces_6_0_io_ins_left[10] ;
 wire \ces_6_0_io_ins_left[11] ;
 wire \ces_6_0_io_ins_left[12] ;
 wire \ces_6_0_io_ins_left[13] ;
 wire \ces_6_0_io_ins_left[14] ;
 wire \ces_6_0_io_ins_left[15] ;
 wire \ces_6_0_io_ins_left[16] ;
 wire \ces_6_0_io_ins_left[17] ;
 wire \ces_6_0_io_ins_left[18] ;
 wire \ces_6_0_io_ins_left[19] ;
 wire \ces_6_0_io_ins_left[1] ;
 wire \ces_6_0_io_ins_left[20] ;
 wire \ces_6_0_io_ins_left[21] ;
 wire \ces_6_0_io_ins_left[22] ;
 wire \ces_6_0_io_ins_left[23] ;
 wire \ces_6_0_io_ins_left[24] ;
 wire \ces_6_0_io_ins_left[25] ;
 wire \ces_6_0_io_ins_left[26] ;
 wire \ces_6_0_io_ins_left[27] ;
 wire \ces_6_0_io_ins_left[28] ;
 wire \ces_6_0_io_ins_left[29] ;
 wire \ces_6_0_io_ins_left[2] ;
 wire \ces_6_0_io_ins_left[30] ;
 wire \ces_6_0_io_ins_left[31] ;
 wire \ces_6_0_io_ins_left[32] ;
 wire \ces_6_0_io_ins_left[33] ;
 wire \ces_6_0_io_ins_left[34] ;
 wire \ces_6_0_io_ins_left[35] ;
 wire \ces_6_0_io_ins_left[36] ;
 wire \ces_6_0_io_ins_left[37] ;
 wire \ces_6_0_io_ins_left[38] ;
 wire \ces_6_0_io_ins_left[39] ;
 wire \ces_6_0_io_ins_left[3] ;
 wire \ces_6_0_io_ins_left[40] ;
 wire \ces_6_0_io_ins_left[41] ;
 wire \ces_6_0_io_ins_left[42] ;
 wire \ces_6_0_io_ins_left[43] ;
 wire \ces_6_0_io_ins_left[44] ;
 wire \ces_6_0_io_ins_left[45] ;
 wire \ces_6_0_io_ins_left[46] ;
 wire \ces_6_0_io_ins_left[47] ;
 wire \ces_6_0_io_ins_left[48] ;
 wire \ces_6_0_io_ins_left[49] ;
 wire \ces_6_0_io_ins_left[4] ;
 wire \ces_6_0_io_ins_left[50] ;
 wire \ces_6_0_io_ins_left[51] ;
 wire \ces_6_0_io_ins_left[52] ;
 wire \ces_6_0_io_ins_left[53] ;
 wire \ces_6_0_io_ins_left[54] ;
 wire \ces_6_0_io_ins_left[55] ;
 wire \ces_6_0_io_ins_left[56] ;
 wire \ces_6_0_io_ins_left[57] ;
 wire \ces_6_0_io_ins_left[58] ;
 wire \ces_6_0_io_ins_left[59] ;
 wire \ces_6_0_io_ins_left[5] ;
 wire \ces_6_0_io_ins_left[60] ;
 wire \ces_6_0_io_ins_left[61] ;
 wire \ces_6_0_io_ins_left[62] ;
 wire \ces_6_0_io_ins_left[63] ;
 wire \ces_6_0_io_ins_left[6] ;
 wire \ces_6_0_io_ins_left[7] ;
 wire \ces_6_0_io_ins_left[8] ;
 wire \ces_6_0_io_ins_left[9] ;
 wire ces_6_0_io_lsbOuts_0;
 wire ces_6_0_io_lsbOuts_1;
 wire ces_6_0_io_lsbOuts_2;
 wire ces_6_0_io_lsbOuts_3;
 wire ces_6_0_io_lsbOuts_4;
 wire ces_6_0_io_lsbOuts_5;
 wire ces_6_0_io_lsbOuts_6;
 wire ces_6_0_io_lsbOuts_7;
 wire \ces_6_0_io_outs_right[0] ;
 wire \ces_6_0_io_outs_right[10] ;
 wire \ces_6_0_io_outs_right[11] ;
 wire \ces_6_0_io_outs_right[12] ;
 wire \ces_6_0_io_outs_right[13] ;
 wire \ces_6_0_io_outs_right[14] ;
 wire \ces_6_0_io_outs_right[15] ;
 wire \ces_6_0_io_outs_right[16] ;
 wire \ces_6_0_io_outs_right[17] ;
 wire \ces_6_0_io_outs_right[18] ;
 wire \ces_6_0_io_outs_right[19] ;
 wire \ces_6_0_io_outs_right[1] ;
 wire \ces_6_0_io_outs_right[20] ;
 wire \ces_6_0_io_outs_right[21] ;
 wire \ces_6_0_io_outs_right[22] ;
 wire \ces_6_0_io_outs_right[23] ;
 wire \ces_6_0_io_outs_right[24] ;
 wire \ces_6_0_io_outs_right[25] ;
 wire \ces_6_0_io_outs_right[26] ;
 wire \ces_6_0_io_outs_right[27] ;
 wire \ces_6_0_io_outs_right[28] ;
 wire \ces_6_0_io_outs_right[29] ;
 wire \ces_6_0_io_outs_right[2] ;
 wire \ces_6_0_io_outs_right[30] ;
 wire \ces_6_0_io_outs_right[31] ;
 wire \ces_6_0_io_outs_right[32] ;
 wire \ces_6_0_io_outs_right[33] ;
 wire \ces_6_0_io_outs_right[34] ;
 wire \ces_6_0_io_outs_right[35] ;
 wire \ces_6_0_io_outs_right[36] ;
 wire \ces_6_0_io_outs_right[37] ;
 wire \ces_6_0_io_outs_right[38] ;
 wire \ces_6_0_io_outs_right[39] ;
 wire \ces_6_0_io_outs_right[3] ;
 wire \ces_6_0_io_outs_right[40] ;
 wire \ces_6_0_io_outs_right[41] ;
 wire \ces_6_0_io_outs_right[42] ;
 wire \ces_6_0_io_outs_right[43] ;
 wire \ces_6_0_io_outs_right[44] ;
 wire \ces_6_0_io_outs_right[45] ;
 wire \ces_6_0_io_outs_right[46] ;
 wire \ces_6_0_io_outs_right[47] ;
 wire \ces_6_0_io_outs_right[48] ;
 wire \ces_6_0_io_outs_right[49] ;
 wire \ces_6_0_io_outs_right[4] ;
 wire \ces_6_0_io_outs_right[50] ;
 wire \ces_6_0_io_outs_right[51] ;
 wire \ces_6_0_io_outs_right[52] ;
 wire \ces_6_0_io_outs_right[53] ;
 wire \ces_6_0_io_outs_right[54] ;
 wire \ces_6_0_io_outs_right[55] ;
 wire \ces_6_0_io_outs_right[56] ;
 wire \ces_6_0_io_outs_right[57] ;
 wire \ces_6_0_io_outs_right[58] ;
 wire \ces_6_0_io_outs_right[59] ;
 wire \ces_6_0_io_outs_right[5] ;
 wire \ces_6_0_io_outs_right[60] ;
 wire \ces_6_0_io_outs_right[61] ;
 wire \ces_6_0_io_outs_right[62] ;
 wire \ces_6_0_io_outs_right[63] ;
 wire \ces_6_0_io_outs_right[6] ;
 wire \ces_6_0_io_outs_right[7] ;
 wire \ces_6_0_io_outs_right[8] ;
 wire \ces_6_0_io_outs_right[9] ;
 wire \ces_6_0_io_outs_up[0] ;
 wire \ces_6_0_io_outs_up[10] ;
 wire \ces_6_0_io_outs_up[11] ;
 wire \ces_6_0_io_outs_up[12] ;
 wire \ces_6_0_io_outs_up[13] ;
 wire \ces_6_0_io_outs_up[14] ;
 wire \ces_6_0_io_outs_up[15] ;
 wire \ces_6_0_io_outs_up[16] ;
 wire \ces_6_0_io_outs_up[17] ;
 wire \ces_6_0_io_outs_up[18] ;
 wire \ces_6_0_io_outs_up[19] ;
 wire \ces_6_0_io_outs_up[1] ;
 wire \ces_6_0_io_outs_up[20] ;
 wire \ces_6_0_io_outs_up[21] ;
 wire \ces_6_0_io_outs_up[22] ;
 wire \ces_6_0_io_outs_up[23] ;
 wire \ces_6_0_io_outs_up[24] ;
 wire \ces_6_0_io_outs_up[25] ;
 wire \ces_6_0_io_outs_up[26] ;
 wire \ces_6_0_io_outs_up[27] ;
 wire \ces_6_0_io_outs_up[28] ;
 wire \ces_6_0_io_outs_up[29] ;
 wire \ces_6_0_io_outs_up[2] ;
 wire \ces_6_0_io_outs_up[30] ;
 wire \ces_6_0_io_outs_up[31] ;
 wire \ces_6_0_io_outs_up[32] ;
 wire \ces_6_0_io_outs_up[33] ;
 wire \ces_6_0_io_outs_up[34] ;
 wire \ces_6_0_io_outs_up[35] ;
 wire \ces_6_0_io_outs_up[36] ;
 wire \ces_6_0_io_outs_up[37] ;
 wire \ces_6_0_io_outs_up[38] ;
 wire \ces_6_0_io_outs_up[39] ;
 wire \ces_6_0_io_outs_up[3] ;
 wire \ces_6_0_io_outs_up[40] ;
 wire \ces_6_0_io_outs_up[41] ;
 wire \ces_6_0_io_outs_up[42] ;
 wire \ces_6_0_io_outs_up[43] ;
 wire \ces_6_0_io_outs_up[44] ;
 wire \ces_6_0_io_outs_up[45] ;
 wire \ces_6_0_io_outs_up[46] ;
 wire \ces_6_0_io_outs_up[47] ;
 wire \ces_6_0_io_outs_up[48] ;
 wire \ces_6_0_io_outs_up[49] ;
 wire \ces_6_0_io_outs_up[4] ;
 wire \ces_6_0_io_outs_up[50] ;
 wire \ces_6_0_io_outs_up[51] ;
 wire \ces_6_0_io_outs_up[52] ;
 wire \ces_6_0_io_outs_up[53] ;
 wire \ces_6_0_io_outs_up[54] ;
 wire \ces_6_0_io_outs_up[55] ;
 wire \ces_6_0_io_outs_up[56] ;
 wire \ces_6_0_io_outs_up[57] ;
 wire \ces_6_0_io_outs_up[58] ;
 wire \ces_6_0_io_outs_up[59] ;
 wire \ces_6_0_io_outs_up[5] ;
 wire \ces_6_0_io_outs_up[60] ;
 wire \ces_6_0_io_outs_up[61] ;
 wire \ces_6_0_io_outs_up[62] ;
 wire \ces_6_0_io_outs_up[63] ;
 wire \ces_6_0_io_outs_up[6] ;
 wire \ces_6_0_io_outs_up[7] ;
 wire \ces_6_0_io_outs_up[8] ;
 wire \ces_6_0_io_outs_up[9] ;
 wire \ces_6_1_io_ins_down[0] ;
 wire \ces_6_1_io_ins_down[10] ;
 wire \ces_6_1_io_ins_down[11] ;
 wire \ces_6_1_io_ins_down[12] ;
 wire \ces_6_1_io_ins_down[13] ;
 wire \ces_6_1_io_ins_down[14] ;
 wire \ces_6_1_io_ins_down[15] ;
 wire \ces_6_1_io_ins_down[16] ;
 wire \ces_6_1_io_ins_down[17] ;
 wire \ces_6_1_io_ins_down[18] ;
 wire \ces_6_1_io_ins_down[19] ;
 wire \ces_6_1_io_ins_down[1] ;
 wire \ces_6_1_io_ins_down[20] ;
 wire \ces_6_1_io_ins_down[21] ;
 wire \ces_6_1_io_ins_down[22] ;
 wire \ces_6_1_io_ins_down[23] ;
 wire \ces_6_1_io_ins_down[24] ;
 wire \ces_6_1_io_ins_down[25] ;
 wire \ces_6_1_io_ins_down[26] ;
 wire \ces_6_1_io_ins_down[27] ;
 wire \ces_6_1_io_ins_down[28] ;
 wire \ces_6_1_io_ins_down[29] ;
 wire \ces_6_1_io_ins_down[2] ;
 wire \ces_6_1_io_ins_down[30] ;
 wire \ces_6_1_io_ins_down[31] ;
 wire \ces_6_1_io_ins_down[32] ;
 wire \ces_6_1_io_ins_down[33] ;
 wire \ces_6_1_io_ins_down[34] ;
 wire \ces_6_1_io_ins_down[35] ;
 wire \ces_6_1_io_ins_down[36] ;
 wire \ces_6_1_io_ins_down[37] ;
 wire \ces_6_1_io_ins_down[38] ;
 wire \ces_6_1_io_ins_down[39] ;
 wire \ces_6_1_io_ins_down[3] ;
 wire \ces_6_1_io_ins_down[40] ;
 wire \ces_6_1_io_ins_down[41] ;
 wire \ces_6_1_io_ins_down[42] ;
 wire \ces_6_1_io_ins_down[43] ;
 wire \ces_6_1_io_ins_down[44] ;
 wire \ces_6_1_io_ins_down[45] ;
 wire \ces_6_1_io_ins_down[46] ;
 wire \ces_6_1_io_ins_down[47] ;
 wire \ces_6_1_io_ins_down[48] ;
 wire \ces_6_1_io_ins_down[49] ;
 wire \ces_6_1_io_ins_down[4] ;
 wire \ces_6_1_io_ins_down[50] ;
 wire \ces_6_1_io_ins_down[51] ;
 wire \ces_6_1_io_ins_down[52] ;
 wire \ces_6_1_io_ins_down[53] ;
 wire \ces_6_1_io_ins_down[54] ;
 wire \ces_6_1_io_ins_down[55] ;
 wire \ces_6_1_io_ins_down[56] ;
 wire \ces_6_1_io_ins_down[57] ;
 wire \ces_6_1_io_ins_down[58] ;
 wire \ces_6_1_io_ins_down[59] ;
 wire \ces_6_1_io_ins_down[5] ;
 wire \ces_6_1_io_ins_down[60] ;
 wire \ces_6_1_io_ins_down[61] ;
 wire \ces_6_1_io_ins_down[62] ;
 wire \ces_6_1_io_ins_down[63] ;
 wire \ces_6_1_io_ins_down[6] ;
 wire \ces_6_1_io_ins_down[7] ;
 wire \ces_6_1_io_ins_down[8] ;
 wire \ces_6_1_io_ins_down[9] ;
 wire \ces_6_1_io_ins_left[0] ;
 wire \ces_6_1_io_ins_left[10] ;
 wire \ces_6_1_io_ins_left[11] ;
 wire \ces_6_1_io_ins_left[12] ;
 wire \ces_6_1_io_ins_left[13] ;
 wire \ces_6_1_io_ins_left[14] ;
 wire \ces_6_1_io_ins_left[15] ;
 wire \ces_6_1_io_ins_left[16] ;
 wire \ces_6_1_io_ins_left[17] ;
 wire \ces_6_1_io_ins_left[18] ;
 wire \ces_6_1_io_ins_left[19] ;
 wire \ces_6_1_io_ins_left[1] ;
 wire \ces_6_1_io_ins_left[20] ;
 wire \ces_6_1_io_ins_left[21] ;
 wire \ces_6_1_io_ins_left[22] ;
 wire \ces_6_1_io_ins_left[23] ;
 wire \ces_6_1_io_ins_left[24] ;
 wire \ces_6_1_io_ins_left[25] ;
 wire \ces_6_1_io_ins_left[26] ;
 wire \ces_6_1_io_ins_left[27] ;
 wire \ces_6_1_io_ins_left[28] ;
 wire \ces_6_1_io_ins_left[29] ;
 wire \ces_6_1_io_ins_left[2] ;
 wire \ces_6_1_io_ins_left[30] ;
 wire \ces_6_1_io_ins_left[31] ;
 wire \ces_6_1_io_ins_left[32] ;
 wire \ces_6_1_io_ins_left[33] ;
 wire \ces_6_1_io_ins_left[34] ;
 wire \ces_6_1_io_ins_left[35] ;
 wire \ces_6_1_io_ins_left[36] ;
 wire \ces_6_1_io_ins_left[37] ;
 wire \ces_6_1_io_ins_left[38] ;
 wire \ces_6_1_io_ins_left[39] ;
 wire \ces_6_1_io_ins_left[3] ;
 wire \ces_6_1_io_ins_left[40] ;
 wire \ces_6_1_io_ins_left[41] ;
 wire \ces_6_1_io_ins_left[42] ;
 wire \ces_6_1_io_ins_left[43] ;
 wire \ces_6_1_io_ins_left[44] ;
 wire \ces_6_1_io_ins_left[45] ;
 wire \ces_6_1_io_ins_left[46] ;
 wire \ces_6_1_io_ins_left[47] ;
 wire \ces_6_1_io_ins_left[48] ;
 wire \ces_6_1_io_ins_left[49] ;
 wire \ces_6_1_io_ins_left[4] ;
 wire \ces_6_1_io_ins_left[50] ;
 wire \ces_6_1_io_ins_left[51] ;
 wire \ces_6_1_io_ins_left[52] ;
 wire \ces_6_1_io_ins_left[53] ;
 wire \ces_6_1_io_ins_left[54] ;
 wire \ces_6_1_io_ins_left[55] ;
 wire \ces_6_1_io_ins_left[56] ;
 wire \ces_6_1_io_ins_left[57] ;
 wire \ces_6_1_io_ins_left[58] ;
 wire \ces_6_1_io_ins_left[59] ;
 wire \ces_6_1_io_ins_left[5] ;
 wire \ces_6_1_io_ins_left[60] ;
 wire \ces_6_1_io_ins_left[61] ;
 wire \ces_6_1_io_ins_left[62] ;
 wire \ces_6_1_io_ins_left[63] ;
 wire \ces_6_1_io_ins_left[6] ;
 wire \ces_6_1_io_ins_left[7] ;
 wire \ces_6_1_io_ins_left[8] ;
 wire \ces_6_1_io_ins_left[9] ;
 wire ces_6_1_io_lsbOuts_0;
 wire ces_6_1_io_lsbOuts_1;
 wire ces_6_1_io_lsbOuts_2;
 wire ces_6_1_io_lsbOuts_3;
 wire ces_6_1_io_lsbOuts_4;
 wire ces_6_1_io_lsbOuts_5;
 wire ces_6_1_io_lsbOuts_6;
 wire ces_6_1_io_lsbOuts_7;
 wire \ces_6_1_io_outs_right[0] ;
 wire \ces_6_1_io_outs_right[10] ;
 wire \ces_6_1_io_outs_right[11] ;
 wire \ces_6_1_io_outs_right[12] ;
 wire \ces_6_1_io_outs_right[13] ;
 wire \ces_6_1_io_outs_right[14] ;
 wire \ces_6_1_io_outs_right[15] ;
 wire \ces_6_1_io_outs_right[16] ;
 wire \ces_6_1_io_outs_right[17] ;
 wire \ces_6_1_io_outs_right[18] ;
 wire \ces_6_1_io_outs_right[19] ;
 wire \ces_6_1_io_outs_right[1] ;
 wire \ces_6_1_io_outs_right[20] ;
 wire \ces_6_1_io_outs_right[21] ;
 wire \ces_6_1_io_outs_right[22] ;
 wire \ces_6_1_io_outs_right[23] ;
 wire \ces_6_1_io_outs_right[24] ;
 wire \ces_6_1_io_outs_right[25] ;
 wire \ces_6_1_io_outs_right[26] ;
 wire \ces_6_1_io_outs_right[27] ;
 wire \ces_6_1_io_outs_right[28] ;
 wire \ces_6_1_io_outs_right[29] ;
 wire \ces_6_1_io_outs_right[2] ;
 wire \ces_6_1_io_outs_right[30] ;
 wire \ces_6_1_io_outs_right[31] ;
 wire \ces_6_1_io_outs_right[32] ;
 wire \ces_6_1_io_outs_right[33] ;
 wire \ces_6_1_io_outs_right[34] ;
 wire \ces_6_1_io_outs_right[35] ;
 wire \ces_6_1_io_outs_right[36] ;
 wire \ces_6_1_io_outs_right[37] ;
 wire \ces_6_1_io_outs_right[38] ;
 wire \ces_6_1_io_outs_right[39] ;
 wire \ces_6_1_io_outs_right[3] ;
 wire \ces_6_1_io_outs_right[40] ;
 wire \ces_6_1_io_outs_right[41] ;
 wire \ces_6_1_io_outs_right[42] ;
 wire \ces_6_1_io_outs_right[43] ;
 wire \ces_6_1_io_outs_right[44] ;
 wire \ces_6_1_io_outs_right[45] ;
 wire \ces_6_1_io_outs_right[46] ;
 wire \ces_6_1_io_outs_right[47] ;
 wire \ces_6_1_io_outs_right[48] ;
 wire \ces_6_1_io_outs_right[49] ;
 wire \ces_6_1_io_outs_right[4] ;
 wire \ces_6_1_io_outs_right[50] ;
 wire \ces_6_1_io_outs_right[51] ;
 wire \ces_6_1_io_outs_right[52] ;
 wire \ces_6_1_io_outs_right[53] ;
 wire \ces_6_1_io_outs_right[54] ;
 wire \ces_6_1_io_outs_right[55] ;
 wire \ces_6_1_io_outs_right[56] ;
 wire \ces_6_1_io_outs_right[57] ;
 wire \ces_6_1_io_outs_right[58] ;
 wire \ces_6_1_io_outs_right[59] ;
 wire \ces_6_1_io_outs_right[5] ;
 wire \ces_6_1_io_outs_right[60] ;
 wire \ces_6_1_io_outs_right[61] ;
 wire \ces_6_1_io_outs_right[62] ;
 wire \ces_6_1_io_outs_right[63] ;
 wire \ces_6_1_io_outs_right[6] ;
 wire \ces_6_1_io_outs_right[7] ;
 wire \ces_6_1_io_outs_right[8] ;
 wire \ces_6_1_io_outs_right[9] ;
 wire \ces_6_1_io_outs_up[0] ;
 wire \ces_6_1_io_outs_up[10] ;
 wire \ces_6_1_io_outs_up[11] ;
 wire \ces_6_1_io_outs_up[12] ;
 wire \ces_6_1_io_outs_up[13] ;
 wire \ces_6_1_io_outs_up[14] ;
 wire \ces_6_1_io_outs_up[15] ;
 wire \ces_6_1_io_outs_up[16] ;
 wire \ces_6_1_io_outs_up[17] ;
 wire \ces_6_1_io_outs_up[18] ;
 wire \ces_6_1_io_outs_up[19] ;
 wire \ces_6_1_io_outs_up[1] ;
 wire \ces_6_1_io_outs_up[20] ;
 wire \ces_6_1_io_outs_up[21] ;
 wire \ces_6_1_io_outs_up[22] ;
 wire \ces_6_1_io_outs_up[23] ;
 wire \ces_6_1_io_outs_up[24] ;
 wire \ces_6_1_io_outs_up[25] ;
 wire \ces_6_1_io_outs_up[26] ;
 wire \ces_6_1_io_outs_up[27] ;
 wire \ces_6_1_io_outs_up[28] ;
 wire \ces_6_1_io_outs_up[29] ;
 wire \ces_6_1_io_outs_up[2] ;
 wire \ces_6_1_io_outs_up[30] ;
 wire \ces_6_1_io_outs_up[31] ;
 wire \ces_6_1_io_outs_up[32] ;
 wire \ces_6_1_io_outs_up[33] ;
 wire \ces_6_1_io_outs_up[34] ;
 wire \ces_6_1_io_outs_up[35] ;
 wire \ces_6_1_io_outs_up[36] ;
 wire \ces_6_1_io_outs_up[37] ;
 wire \ces_6_1_io_outs_up[38] ;
 wire \ces_6_1_io_outs_up[39] ;
 wire \ces_6_1_io_outs_up[3] ;
 wire \ces_6_1_io_outs_up[40] ;
 wire \ces_6_1_io_outs_up[41] ;
 wire \ces_6_1_io_outs_up[42] ;
 wire \ces_6_1_io_outs_up[43] ;
 wire \ces_6_1_io_outs_up[44] ;
 wire \ces_6_1_io_outs_up[45] ;
 wire \ces_6_1_io_outs_up[46] ;
 wire \ces_6_1_io_outs_up[47] ;
 wire \ces_6_1_io_outs_up[48] ;
 wire \ces_6_1_io_outs_up[49] ;
 wire \ces_6_1_io_outs_up[4] ;
 wire \ces_6_1_io_outs_up[50] ;
 wire \ces_6_1_io_outs_up[51] ;
 wire \ces_6_1_io_outs_up[52] ;
 wire \ces_6_1_io_outs_up[53] ;
 wire \ces_6_1_io_outs_up[54] ;
 wire \ces_6_1_io_outs_up[55] ;
 wire \ces_6_1_io_outs_up[56] ;
 wire \ces_6_1_io_outs_up[57] ;
 wire \ces_6_1_io_outs_up[58] ;
 wire \ces_6_1_io_outs_up[59] ;
 wire \ces_6_1_io_outs_up[5] ;
 wire \ces_6_1_io_outs_up[60] ;
 wire \ces_6_1_io_outs_up[61] ;
 wire \ces_6_1_io_outs_up[62] ;
 wire \ces_6_1_io_outs_up[63] ;
 wire \ces_6_1_io_outs_up[6] ;
 wire \ces_6_1_io_outs_up[7] ;
 wire \ces_6_1_io_outs_up[8] ;
 wire \ces_6_1_io_outs_up[9] ;
 wire \ces_6_2_io_ins_down[0] ;
 wire \ces_6_2_io_ins_down[10] ;
 wire \ces_6_2_io_ins_down[11] ;
 wire \ces_6_2_io_ins_down[12] ;
 wire \ces_6_2_io_ins_down[13] ;
 wire \ces_6_2_io_ins_down[14] ;
 wire \ces_6_2_io_ins_down[15] ;
 wire \ces_6_2_io_ins_down[16] ;
 wire \ces_6_2_io_ins_down[17] ;
 wire \ces_6_2_io_ins_down[18] ;
 wire \ces_6_2_io_ins_down[19] ;
 wire \ces_6_2_io_ins_down[1] ;
 wire \ces_6_2_io_ins_down[20] ;
 wire \ces_6_2_io_ins_down[21] ;
 wire \ces_6_2_io_ins_down[22] ;
 wire \ces_6_2_io_ins_down[23] ;
 wire \ces_6_2_io_ins_down[24] ;
 wire \ces_6_2_io_ins_down[25] ;
 wire \ces_6_2_io_ins_down[26] ;
 wire \ces_6_2_io_ins_down[27] ;
 wire \ces_6_2_io_ins_down[28] ;
 wire \ces_6_2_io_ins_down[29] ;
 wire \ces_6_2_io_ins_down[2] ;
 wire \ces_6_2_io_ins_down[30] ;
 wire \ces_6_2_io_ins_down[31] ;
 wire \ces_6_2_io_ins_down[32] ;
 wire \ces_6_2_io_ins_down[33] ;
 wire \ces_6_2_io_ins_down[34] ;
 wire \ces_6_2_io_ins_down[35] ;
 wire \ces_6_2_io_ins_down[36] ;
 wire \ces_6_2_io_ins_down[37] ;
 wire \ces_6_2_io_ins_down[38] ;
 wire \ces_6_2_io_ins_down[39] ;
 wire \ces_6_2_io_ins_down[3] ;
 wire \ces_6_2_io_ins_down[40] ;
 wire \ces_6_2_io_ins_down[41] ;
 wire \ces_6_2_io_ins_down[42] ;
 wire \ces_6_2_io_ins_down[43] ;
 wire \ces_6_2_io_ins_down[44] ;
 wire \ces_6_2_io_ins_down[45] ;
 wire \ces_6_2_io_ins_down[46] ;
 wire \ces_6_2_io_ins_down[47] ;
 wire \ces_6_2_io_ins_down[48] ;
 wire \ces_6_2_io_ins_down[49] ;
 wire \ces_6_2_io_ins_down[4] ;
 wire \ces_6_2_io_ins_down[50] ;
 wire \ces_6_2_io_ins_down[51] ;
 wire \ces_6_2_io_ins_down[52] ;
 wire \ces_6_2_io_ins_down[53] ;
 wire \ces_6_2_io_ins_down[54] ;
 wire \ces_6_2_io_ins_down[55] ;
 wire \ces_6_2_io_ins_down[56] ;
 wire \ces_6_2_io_ins_down[57] ;
 wire \ces_6_2_io_ins_down[58] ;
 wire \ces_6_2_io_ins_down[59] ;
 wire \ces_6_2_io_ins_down[5] ;
 wire \ces_6_2_io_ins_down[60] ;
 wire \ces_6_2_io_ins_down[61] ;
 wire \ces_6_2_io_ins_down[62] ;
 wire \ces_6_2_io_ins_down[63] ;
 wire \ces_6_2_io_ins_down[6] ;
 wire \ces_6_2_io_ins_down[7] ;
 wire \ces_6_2_io_ins_down[8] ;
 wire \ces_6_2_io_ins_down[9] ;
 wire \ces_6_2_io_ins_left[0] ;
 wire \ces_6_2_io_ins_left[10] ;
 wire \ces_6_2_io_ins_left[11] ;
 wire \ces_6_2_io_ins_left[12] ;
 wire \ces_6_2_io_ins_left[13] ;
 wire \ces_6_2_io_ins_left[14] ;
 wire \ces_6_2_io_ins_left[15] ;
 wire \ces_6_2_io_ins_left[16] ;
 wire \ces_6_2_io_ins_left[17] ;
 wire \ces_6_2_io_ins_left[18] ;
 wire \ces_6_2_io_ins_left[19] ;
 wire \ces_6_2_io_ins_left[1] ;
 wire \ces_6_2_io_ins_left[20] ;
 wire \ces_6_2_io_ins_left[21] ;
 wire \ces_6_2_io_ins_left[22] ;
 wire \ces_6_2_io_ins_left[23] ;
 wire \ces_6_2_io_ins_left[24] ;
 wire \ces_6_2_io_ins_left[25] ;
 wire \ces_6_2_io_ins_left[26] ;
 wire \ces_6_2_io_ins_left[27] ;
 wire \ces_6_2_io_ins_left[28] ;
 wire \ces_6_2_io_ins_left[29] ;
 wire \ces_6_2_io_ins_left[2] ;
 wire \ces_6_2_io_ins_left[30] ;
 wire \ces_6_2_io_ins_left[31] ;
 wire \ces_6_2_io_ins_left[32] ;
 wire \ces_6_2_io_ins_left[33] ;
 wire \ces_6_2_io_ins_left[34] ;
 wire \ces_6_2_io_ins_left[35] ;
 wire \ces_6_2_io_ins_left[36] ;
 wire \ces_6_2_io_ins_left[37] ;
 wire \ces_6_2_io_ins_left[38] ;
 wire \ces_6_2_io_ins_left[39] ;
 wire \ces_6_2_io_ins_left[3] ;
 wire \ces_6_2_io_ins_left[40] ;
 wire \ces_6_2_io_ins_left[41] ;
 wire \ces_6_2_io_ins_left[42] ;
 wire \ces_6_2_io_ins_left[43] ;
 wire \ces_6_2_io_ins_left[44] ;
 wire \ces_6_2_io_ins_left[45] ;
 wire \ces_6_2_io_ins_left[46] ;
 wire \ces_6_2_io_ins_left[47] ;
 wire \ces_6_2_io_ins_left[48] ;
 wire \ces_6_2_io_ins_left[49] ;
 wire \ces_6_2_io_ins_left[4] ;
 wire \ces_6_2_io_ins_left[50] ;
 wire \ces_6_2_io_ins_left[51] ;
 wire \ces_6_2_io_ins_left[52] ;
 wire \ces_6_2_io_ins_left[53] ;
 wire \ces_6_2_io_ins_left[54] ;
 wire \ces_6_2_io_ins_left[55] ;
 wire \ces_6_2_io_ins_left[56] ;
 wire \ces_6_2_io_ins_left[57] ;
 wire \ces_6_2_io_ins_left[58] ;
 wire \ces_6_2_io_ins_left[59] ;
 wire \ces_6_2_io_ins_left[5] ;
 wire \ces_6_2_io_ins_left[60] ;
 wire \ces_6_2_io_ins_left[61] ;
 wire \ces_6_2_io_ins_left[62] ;
 wire \ces_6_2_io_ins_left[63] ;
 wire \ces_6_2_io_ins_left[6] ;
 wire \ces_6_2_io_ins_left[7] ;
 wire \ces_6_2_io_ins_left[8] ;
 wire \ces_6_2_io_ins_left[9] ;
 wire ces_6_2_io_lsbOuts_0;
 wire ces_6_2_io_lsbOuts_1;
 wire ces_6_2_io_lsbOuts_2;
 wire ces_6_2_io_lsbOuts_3;
 wire ces_6_2_io_lsbOuts_4;
 wire ces_6_2_io_lsbOuts_5;
 wire ces_6_2_io_lsbOuts_6;
 wire ces_6_2_io_lsbOuts_7;
 wire \ces_6_2_io_outs_right[0] ;
 wire \ces_6_2_io_outs_right[10] ;
 wire \ces_6_2_io_outs_right[11] ;
 wire \ces_6_2_io_outs_right[12] ;
 wire \ces_6_2_io_outs_right[13] ;
 wire \ces_6_2_io_outs_right[14] ;
 wire \ces_6_2_io_outs_right[15] ;
 wire \ces_6_2_io_outs_right[16] ;
 wire \ces_6_2_io_outs_right[17] ;
 wire \ces_6_2_io_outs_right[18] ;
 wire \ces_6_2_io_outs_right[19] ;
 wire \ces_6_2_io_outs_right[1] ;
 wire \ces_6_2_io_outs_right[20] ;
 wire \ces_6_2_io_outs_right[21] ;
 wire \ces_6_2_io_outs_right[22] ;
 wire \ces_6_2_io_outs_right[23] ;
 wire \ces_6_2_io_outs_right[24] ;
 wire \ces_6_2_io_outs_right[25] ;
 wire \ces_6_2_io_outs_right[26] ;
 wire \ces_6_2_io_outs_right[27] ;
 wire \ces_6_2_io_outs_right[28] ;
 wire \ces_6_2_io_outs_right[29] ;
 wire \ces_6_2_io_outs_right[2] ;
 wire \ces_6_2_io_outs_right[30] ;
 wire \ces_6_2_io_outs_right[31] ;
 wire \ces_6_2_io_outs_right[32] ;
 wire \ces_6_2_io_outs_right[33] ;
 wire \ces_6_2_io_outs_right[34] ;
 wire \ces_6_2_io_outs_right[35] ;
 wire \ces_6_2_io_outs_right[36] ;
 wire \ces_6_2_io_outs_right[37] ;
 wire \ces_6_2_io_outs_right[38] ;
 wire \ces_6_2_io_outs_right[39] ;
 wire \ces_6_2_io_outs_right[3] ;
 wire \ces_6_2_io_outs_right[40] ;
 wire \ces_6_2_io_outs_right[41] ;
 wire \ces_6_2_io_outs_right[42] ;
 wire \ces_6_2_io_outs_right[43] ;
 wire \ces_6_2_io_outs_right[44] ;
 wire \ces_6_2_io_outs_right[45] ;
 wire \ces_6_2_io_outs_right[46] ;
 wire \ces_6_2_io_outs_right[47] ;
 wire \ces_6_2_io_outs_right[48] ;
 wire \ces_6_2_io_outs_right[49] ;
 wire \ces_6_2_io_outs_right[4] ;
 wire \ces_6_2_io_outs_right[50] ;
 wire \ces_6_2_io_outs_right[51] ;
 wire \ces_6_2_io_outs_right[52] ;
 wire \ces_6_2_io_outs_right[53] ;
 wire \ces_6_2_io_outs_right[54] ;
 wire \ces_6_2_io_outs_right[55] ;
 wire \ces_6_2_io_outs_right[56] ;
 wire \ces_6_2_io_outs_right[57] ;
 wire \ces_6_2_io_outs_right[58] ;
 wire \ces_6_2_io_outs_right[59] ;
 wire \ces_6_2_io_outs_right[5] ;
 wire \ces_6_2_io_outs_right[60] ;
 wire \ces_6_2_io_outs_right[61] ;
 wire \ces_6_2_io_outs_right[62] ;
 wire \ces_6_2_io_outs_right[63] ;
 wire \ces_6_2_io_outs_right[6] ;
 wire \ces_6_2_io_outs_right[7] ;
 wire \ces_6_2_io_outs_right[8] ;
 wire \ces_6_2_io_outs_right[9] ;
 wire \ces_6_2_io_outs_up[0] ;
 wire \ces_6_2_io_outs_up[10] ;
 wire \ces_6_2_io_outs_up[11] ;
 wire \ces_6_2_io_outs_up[12] ;
 wire \ces_6_2_io_outs_up[13] ;
 wire \ces_6_2_io_outs_up[14] ;
 wire \ces_6_2_io_outs_up[15] ;
 wire \ces_6_2_io_outs_up[16] ;
 wire \ces_6_2_io_outs_up[17] ;
 wire \ces_6_2_io_outs_up[18] ;
 wire \ces_6_2_io_outs_up[19] ;
 wire \ces_6_2_io_outs_up[1] ;
 wire \ces_6_2_io_outs_up[20] ;
 wire \ces_6_2_io_outs_up[21] ;
 wire \ces_6_2_io_outs_up[22] ;
 wire \ces_6_2_io_outs_up[23] ;
 wire \ces_6_2_io_outs_up[24] ;
 wire \ces_6_2_io_outs_up[25] ;
 wire \ces_6_2_io_outs_up[26] ;
 wire \ces_6_2_io_outs_up[27] ;
 wire \ces_6_2_io_outs_up[28] ;
 wire \ces_6_2_io_outs_up[29] ;
 wire \ces_6_2_io_outs_up[2] ;
 wire \ces_6_2_io_outs_up[30] ;
 wire \ces_6_2_io_outs_up[31] ;
 wire \ces_6_2_io_outs_up[32] ;
 wire \ces_6_2_io_outs_up[33] ;
 wire \ces_6_2_io_outs_up[34] ;
 wire \ces_6_2_io_outs_up[35] ;
 wire \ces_6_2_io_outs_up[36] ;
 wire \ces_6_2_io_outs_up[37] ;
 wire \ces_6_2_io_outs_up[38] ;
 wire \ces_6_2_io_outs_up[39] ;
 wire \ces_6_2_io_outs_up[3] ;
 wire \ces_6_2_io_outs_up[40] ;
 wire \ces_6_2_io_outs_up[41] ;
 wire \ces_6_2_io_outs_up[42] ;
 wire \ces_6_2_io_outs_up[43] ;
 wire \ces_6_2_io_outs_up[44] ;
 wire \ces_6_2_io_outs_up[45] ;
 wire \ces_6_2_io_outs_up[46] ;
 wire \ces_6_2_io_outs_up[47] ;
 wire \ces_6_2_io_outs_up[48] ;
 wire \ces_6_2_io_outs_up[49] ;
 wire \ces_6_2_io_outs_up[4] ;
 wire \ces_6_2_io_outs_up[50] ;
 wire \ces_6_2_io_outs_up[51] ;
 wire \ces_6_2_io_outs_up[52] ;
 wire \ces_6_2_io_outs_up[53] ;
 wire \ces_6_2_io_outs_up[54] ;
 wire \ces_6_2_io_outs_up[55] ;
 wire \ces_6_2_io_outs_up[56] ;
 wire \ces_6_2_io_outs_up[57] ;
 wire \ces_6_2_io_outs_up[58] ;
 wire \ces_6_2_io_outs_up[59] ;
 wire \ces_6_2_io_outs_up[5] ;
 wire \ces_6_2_io_outs_up[60] ;
 wire \ces_6_2_io_outs_up[61] ;
 wire \ces_6_2_io_outs_up[62] ;
 wire \ces_6_2_io_outs_up[63] ;
 wire \ces_6_2_io_outs_up[6] ;
 wire \ces_6_2_io_outs_up[7] ;
 wire \ces_6_2_io_outs_up[8] ;
 wire \ces_6_2_io_outs_up[9] ;
 wire \ces_6_3_io_ins_down[0] ;
 wire \ces_6_3_io_ins_down[10] ;
 wire \ces_6_3_io_ins_down[11] ;
 wire \ces_6_3_io_ins_down[12] ;
 wire \ces_6_3_io_ins_down[13] ;
 wire \ces_6_3_io_ins_down[14] ;
 wire \ces_6_3_io_ins_down[15] ;
 wire \ces_6_3_io_ins_down[16] ;
 wire \ces_6_3_io_ins_down[17] ;
 wire \ces_6_3_io_ins_down[18] ;
 wire \ces_6_3_io_ins_down[19] ;
 wire \ces_6_3_io_ins_down[1] ;
 wire \ces_6_3_io_ins_down[20] ;
 wire \ces_6_3_io_ins_down[21] ;
 wire \ces_6_3_io_ins_down[22] ;
 wire \ces_6_3_io_ins_down[23] ;
 wire \ces_6_3_io_ins_down[24] ;
 wire \ces_6_3_io_ins_down[25] ;
 wire \ces_6_3_io_ins_down[26] ;
 wire \ces_6_3_io_ins_down[27] ;
 wire \ces_6_3_io_ins_down[28] ;
 wire \ces_6_3_io_ins_down[29] ;
 wire \ces_6_3_io_ins_down[2] ;
 wire \ces_6_3_io_ins_down[30] ;
 wire \ces_6_3_io_ins_down[31] ;
 wire \ces_6_3_io_ins_down[32] ;
 wire \ces_6_3_io_ins_down[33] ;
 wire \ces_6_3_io_ins_down[34] ;
 wire \ces_6_3_io_ins_down[35] ;
 wire \ces_6_3_io_ins_down[36] ;
 wire \ces_6_3_io_ins_down[37] ;
 wire \ces_6_3_io_ins_down[38] ;
 wire \ces_6_3_io_ins_down[39] ;
 wire \ces_6_3_io_ins_down[3] ;
 wire \ces_6_3_io_ins_down[40] ;
 wire \ces_6_3_io_ins_down[41] ;
 wire \ces_6_3_io_ins_down[42] ;
 wire \ces_6_3_io_ins_down[43] ;
 wire \ces_6_3_io_ins_down[44] ;
 wire \ces_6_3_io_ins_down[45] ;
 wire \ces_6_3_io_ins_down[46] ;
 wire \ces_6_3_io_ins_down[47] ;
 wire \ces_6_3_io_ins_down[48] ;
 wire \ces_6_3_io_ins_down[49] ;
 wire \ces_6_3_io_ins_down[4] ;
 wire \ces_6_3_io_ins_down[50] ;
 wire \ces_6_3_io_ins_down[51] ;
 wire \ces_6_3_io_ins_down[52] ;
 wire \ces_6_3_io_ins_down[53] ;
 wire \ces_6_3_io_ins_down[54] ;
 wire \ces_6_3_io_ins_down[55] ;
 wire \ces_6_3_io_ins_down[56] ;
 wire \ces_6_3_io_ins_down[57] ;
 wire \ces_6_3_io_ins_down[58] ;
 wire \ces_6_3_io_ins_down[59] ;
 wire \ces_6_3_io_ins_down[5] ;
 wire \ces_6_3_io_ins_down[60] ;
 wire \ces_6_3_io_ins_down[61] ;
 wire \ces_6_3_io_ins_down[62] ;
 wire \ces_6_3_io_ins_down[63] ;
 wire \ces_6_3_io_ins_down[6] ;
 wire \ces_6_3_io_ins_down[7] ;
 wire \ces_6_3_io_ins_down[8] ;
 wire \ces_6_3_io_ins_down[9] ;
 wire \ces_6_3_io_ins_left[0] ;
 wire \ces_6_3_io_ins_left[10] ;
 wire \ces_6_3_io_ins_left[11] ;
 wire \ces_6_3_io_ins_left[12] ;
 wire \ces_6_3_io_ins_left[13] ;
 wire \ces_6_3_io_ins_left[14] ;
 wire \ces_6_3_io_ins_left[15] ;
 wire \ces_6_3_io_ins_left[16] ;
 wire \ces_6_3_io_ins_left[17] ;
 wire \ces_6_3_io_ins_left[18] ;
 wire \ces_6_3_io_ins_left[19] ;
 wire \ces_6_3_io_ins_left[1] ;
 wire \ces_6_3_io_ins_left[20] ;
 wire \ces_6_3_io_ins_left[21] ;
 wire \ces_6_3_io_ins_left[22] ;
 wire \ces_6_3_io_ins_left[23] ;
 wire \ces_6_3_io_ins_left[24] ;
 wire \ces_6_3_io_ins_left[25] ;
 wire \ces_6_3_io_ins_left[26] ;
 wire \ces_6_3_io_ins_left[27] ;
 wire \ces_6_3_io_ins_left[28] ;
 wire \ces_6_3_io_ins_left[29] ;
 wire \ces_6_3_io_ins_left[2] ;
 wire \ces_6_3_io_ins_left[30] ;
 wire \ces_6_3_io_ins_left[31] ;
 wire \ces_6_3_io_ins_left[32] ;
 wire \ces_6_3_io_ins_left[33] ;
 wire \ces_6_3_io_ins_left[34] ;
 wire \ces_6_3_io_ins_left[35] ;
 wire \ces_6_3_io_ins_left[36] ;
 wire \ces_6_3_io_ins_left[37] ;
 wire \ces_6_3_io_ins_left[38] ;
 wire \ces_6_3_io_ins_left[39] ;
 wire \ces_6_3_io_ins_left[3] ;
 wire \ces_6_3_io_ins_left[40] ;
 wire \ces_6_3_io_ins_left[41] ;
 wire \ces_6_3_io_ins_left[42] ;
 wire \ces_6_3_io_ins_left[43] ;
 wire \ces_6_3_io_ins_left[44] ;
 wire \ces_6_3_io_ins_left[45] ;
 wire \ces_6_3_io_ins_left[46] ;
 wire \ces_6_3_io_ins_left[47] ;
 wire \ces_6_3_io_ins_left[48] ;
 wire \ces_6_3_io_ins_left[49] ;
 wire \ces_6_3_io_ins_left[4] ;
 wire \ces_6_3_io_ins_left[50] ;
 wire \ces_6_3_io_ins_left[51] ;
 wire \ces_6_3_io_ins_left[52] ;
 wire \ces_6_3_io_ins_left[53] ;
 wire \ces_6_3_io_ins_left[54] ;
 wire \ces_6_3_io_ins_left[55] ;
 wire \ces_6_3_io_ins_left[56] ;
 wire \ces_6_3_io_ins_left[57] ;
 wire \ces_6_3_io_ins_left[58] ;
 wire \ces_6_3_io_ins_left[59] ;
 wire \ces_6_3_io_ins_left[5] ;
 wire \ces_6_3_io_ins_left[60] ;
 wire \ces_6_3_io_ins_left[61] ;
 wire \ces_6_3_io_ins_left[62] ;
 wire \ces_6_3_io_ins_left[63] ;
 wire \ces_6_3_io_ins_left[6] ;
 wire \ces_6_3_io_ins_left[7] ;
 wire \ces_6_3_io_ins_left[8] ;
 wire \ces_6_3_io_ins_left[9] ;
 wire ces_6_3_io_lsbOuts_0;
 wire ces_6_3_io_lsbOuts_1;
 wire ces_6_3_io_lsbOuts_2;
 wire ces_6_3_io_lsbOuts_3;
 wire ces_6_3_io_lsbOuts_4;
 wire ces_6_3_io_lsbOuts_5;
 wire ces_6_3_io_lsbOuts_6;
 wire ces_6_3_io_lsbOuts_7;
 wire \ces_6_3_io_outs_right[0] ;
 wire \ces_6_3_io_outs_right[10] ;
 wire \ces_6_3_io_outs_right[11] ;
 wire \ces_6_3_io_outs_right[12] ;
 wire \ces_6_3_io_outs_right[13] ;
 wire \ces_6_3_io_outs_right[14] ;
 wire \ces_6_3_io_outs_right[15] ;
 wire \ces_6_3_io_outs_right[16] ;
 wire \ces_6_3_io_outs_right[17] ;
 wire \ces_6_3_io_outs_right[18] ;
 wire \ces_6_3_io_outs_right[19] ;
 wire \ces_6_3_io_outs_right[1] ;
 wire \ces_6_3_io_outs_right[20] ;
 wire \ces_6_3_io_outs_right[21] ;
 wire \ces_6_3_io_outs_right[22] ;
 wire \ces_6_3_io_outs_right[23] ;
 wire \ces_6_3_io_outs_right[24] ;
 wire \ces_6_3_io_outs_right[25] ;
 wire \ces_6_3_io_outs_right[26] ;
 wire \ces_6_3_io_outs_right[27] ;
 wire \ces_6_3_io_outs_right[28] ;
 wire \ces_6_3_io_outs_right[29] ;
 wire \ces_6_3_io_outs_right[2] ;
 wire \ces_6_3_io_outs_right[30] ;
 wire \ces_6_3_io_outs_right[31] ;
 wire \ces_6_3_io_outs_right[32] ;
 wire \ces_6_3_io_outs_right[33] ;
 wire \ces_6_3_io_outs_right[34] ;
 wire \ces_6_3_io_outs_right[35] ;
 wire \ces_6_3_io_outs_right[36] ;
 wire \ces_6_3_io_outs_right[37] ;
 wire \ces_6_3_io_outs_right[38] ;
 wire \ces_6_3_io_outs_right[39] ;
 wire \ces_6_3_io_outs_right[3] ;
 wire \ces_6_3_io_outs_right[40] ;
 wire \ces_6_3_io_outs_right[41] ;
 wire \ces_6_3_io_outs_right[42] ;
 wire \ces_6_3_io_outs_right[43] ;
 wire \ces_6_3_io_outs_right[44] ;
 wire \ces_6_3_io_outs_right[45] ;
 wire \ces_6_3_io_outs_right[46] ;
 wire \ces_6_3_io_outs_right[47] ;
 wire \ces_6_3_io_outs_right[48] ;
 wire \ces_6_3_io_outs_right[49] ;
 wire \ces_6_3_io_outs_right[4] ;
 wire \ces_6_3_io_outs_right[50] ;
 wire \ces_6_3_io_outs_right[51] ;
 wire \ces_6_3_io_outs_right[52] ;
 wire \ces_6_3_io_outs_right[53] ;
 wire \ces_6_3_io_outs_right[54] ;
 wire \ces_6_3_io_outs_right[55] ;
 wire \ces_6_3_io_outs_right[56] ;
 wire \ces_6_3_io_outs_right[57] ;
 wire \ces_6_3_io_outs_right[58] ;
 wire \ces_6_3_io_outs_right[59] ;
 wire \ces_6_3_io_outs_right[5] ;
 wire \ces_6_3_io_outs_right[60] ;
 wire \ces_6_3_io_outs_right[61] ;
 wire \ces_6_3_io_outs_right[62] ;
 wire \ces_6_3_io_outs_right[63] ;
 wire \ces_6_3_io_outs_right[6] ;
 wire \ces_6_3_io_outs_right[7] ;
 wire \ces_6_3_io_outs_right[8] ;
 wire \ces_6_3_io_outs_right[9] ;
 wire \ces_6_3_io_outs_up[0] ;
 wire \ces_6_3_io_outs_up[10] ;
 wire \ces_6_3_io_outs_up[11] ;
 wire \ces_6_3_io_outs_up[12] ;
 wire \ces_6_3_io_outs_up[13] ;
 wire \ces_6_3_io_outs_up[14] ;
 wire \ces_6_3_io_outs_up[15] ;
 wire \ces_6_3_io_outs_up[16] ;
 wire \ces_6_3_io_outs_up[17] ;
 wire \ces_6_3_io_outs_up[18] ;
 wire \ces_6_3_io_outs_up[19] ;
 wire \ces_6_3_io_outs_up[1] ;
 wire \ces_6_3_io_outs_up[20] ;
 wire \ces_6_3_io_outs_up[21] ;
 wire \ces_6_3_io_outs_up[22] ;
 wire \ces_6_3_io_outs_up[23] ;
 wire \ces_6_3_io_outs_up[24] ;
 wire \ces_6_3_io_outs_up[25] ;
 wire \ces_6_3_io_outs_up[26] ;
 wire \ces_6_3_io_outs_up[27] ;
 wire \ces_6_3_io_outs_up[28] ;
 wire \ces_6_3_io_outs_up[29] ;
 wire \ces_6_3_io_outs_up[2] ;
 wire \ces_6_3_io_outs_up[30] ;
 wire \ces_6_3_io_outs_up[31] ;
 wire \ces_6_3_io_outs_up[32] ;
 wire \ces_6_3_io_outs_up[33] ;
 wire \ces_6_3_io_outs_up[34] ;
 wire \ces_6_3_io_outs_up[35] ;
 wire \ces_6_3_io_outs_up[36] ;
 wire \ces_6_3_io_outs_up[37] ;
 wire \ces_6_3_io_outs_up[38] ;
 wire \ces_6_3_io_outs_up[39] ;
 wire \ces_6_3_io_outs_up[3] ;
 wire \ces_6_3_io_outs_up[40] ;
 wire \ces_6_3_io_outs_up[41] ;
 wire \ces_6_3_io_outs_up[42] ;
 wire \ces_6_3_io_outs_up[43] ;
 wire \ces_6_3_io_outs_up[44] ;
 wire \ces_6_3_io_outs_up[45] ;
 wire \ces_6_3_io_outs_up[46] ;
 wire \ces_6_3_io_outs_up[47] ;
 wire \ces_6_3_io_outs_up[48] ;
 wire \ces_6_3_io_outs_up[49] ;
 wire \ces_6_3_io_outs_up[4] ;
 wire \ces_6_3_io_outs_up[50] ;
 wire \ces_6_3_io_outs_up[51] ;
 wire \ces_6_3_io_outs_up[52] ;
 wire \ces_6_3_io_outs_up[53] ;
 wire \ces_6_3_io_outs_up[54] ;
 wire \ces_6_3_io_outs_up[55] ;
 wire \ces_6_3_io_outs_up[56] ;
 wire \ces_6_3_io_outs_up[57] ;
 wire \ces_6_3_io_outs_up[58] ;
 wire \ces_6_3_io_outs_up[59] ;
 wire \ces_6_3_io_outs_up[5] ;
 wire \ces_6_3_io_outs_up[60] ;
 wire \ces_6_3_io_outs_up[61] ;
 wire \ces_6_3_io_outs_up[62] ;
 wire \ces_6_3_io_outs_up[63] ;
 wire \ces_6_3_io_outs_up[6] ;
 wire \ces_6_3_io_outs_up[7] ;
 wire \ces_6_3_io_outs_up[8] ;
 wire \ces_6_3_io_outs_up[9] ;
 wire \ces_6_4_io_ins_down[0] ;
 wire \ces_6_4_io_ins_down[10] ;
 wire \ces_6_4_io_ins_down[11] ;
 wire \ces_6_4_io_ins_down[12] ;
 wire \ces_6_4_io_ins_down[13] ;
 wire \ces_6_4_io_ins_down[14] ;
 wire \ces_6_4_io_ins_down[15] ;
 wire \ces_6_4_io_ins_down[16] ;
 wire \ces_6_4_io_ins_down[17] ;
 wire \ces_6_4_io_ins_down[18] ;
 wire \ces_6_4_io_ins_down[19] ;
 wire \ces_6_4_io_ins_down[1] ;
 wire \ces_6_4_io_ins_down[20] ;
 wire \ces_6_4_io_ins_down[21] ;
 wire \ces_6_4_io_ins_down[22] ;
 wire \ces_6_4_io_ins_down[23] ;
 wire \ces_6_4_io_ins_down[24] ;
 wire \ces_6_4_io_ins_down[25] ;
 wire \ces_6_4_io_ins_down[26] ;
 wire \ces_6_4_io_ins_down[27] ;
 wire \ces_6_4_io_ins_down[28] ;
 wire \ces_6_4_io_ins_down[29] ;
 wire \ces_6_4_io_ins_down[2] ;
 wire \ces_6_4_io_ins_down[30] ;
 wire \ces_6_4_io_ins_down[31] ;
 wire \ces_6_4_io_ins_down[32] ;
 wire \ces_6_4_io_ins_down[33] ;
 wire \ces_6_4_io_ins_down[34] ;
 wire \ces_6_4_io_ins_down[35] ;
 wire \ces_6_4_io_ins_down[36] ;
 wire \ces_6_4_io_ins_down[37] ;
 wire \ces_6_4_io_ins_down[38] ;
 wire \ces_6_4_io_ins_down[39] ;
 wire \ces_6_4_io_ins_down[3] ;
 wire \ces_6_4_io_ins_down[40] ;
 wire \ces_6_4_io_ins_down[41] ;
 wire \ces_6_4_io_ins_down[42] ;
 wire \ces_6_4_io_ins_down[43] ;
 wire \ces_6_4_io_ins_down[44] ;
 wire \ces_6_4_io_ins_down[45] ;
 wire \ces_6_4_io_ins_down[46] ;
 wire \ces_6_4_io_ins_down[47] ;
 wire \ces_6_4_io_ins_down[48] ;
 wire \ces_6_4_io_ins_down[49] ;
 wire \ces_6_4_io_ins_down[4] ;
 wire \ces_6_4_io_ins_down[50] ;
 wire \ces_6_4_io_ins_down[51] ;
 wire \ces_6_4_io_ins_down[52] ;
 wire \ces_6_4_io_ins_down[53] ;
 wire \ces_6_4_io_ins_down[54] ;
 wire \ces_6_4_io_ins_down[55] ;
 wire \ces_6_4_io_ins_down[56] ;
 wire \ces_6_4_io_ins_down[57] ;
 wire \ces_6_4_io_ins_down[58] ;
 wire \ces_6_4_io_ins_down[59] ;
 wire \ces_6_4_io_ins_down[5] ;
 wire \ces_6_4_io_ins_down[60] ;
 wire \ces_6_4_io_ins_down[61] ;
 wire \ces_6_4_io_ins_down[62] ;
 wire \ces_6_4_io_ins_down[63] ;
 wire \ces_6_4_io_ins_down[6] ;
 wire \ces_6_4_io_ins_down[7] ;
 wire \ces_6_4_io_ins_down[8] ;
 wire \ces_6_4_io_ins_down[9] ;
 wire \ces_6_4_io_ins_left[0] ;
 wire \ces_6_4_io_ins_left[10] ;
 wire \ces_6_4_io_ins_left[11] ;
 wire \ces_6_4_io_ins_left[12] ;
 wire \ces_6_4_io_ins_left[13] ;
 wire \ces_6_4_io_ins_left[14] ;
 wire \ces_6_4_io_ins_left[15] ;
 wire \ces_6_4_io_ins_left[16] ;
 wire \ces_6_4_io_ins_left[17] ;
 wire \ces_6_4_io_ins_left[18] ;
 wire \ces_6_4_io_ins_left[19] ;
 wire \ces_6_4_io_ins_left[1] ;
 wire \ces_6_4_io_ins_left[20] ;
 wire \ces_6_4_io_ins_left[21] ;
 wire \ces_6_4_io_ins_left[22] ;
 wire \ces_6_4_io_ins_left[23] ;
 wire \ces_6_4_io_ins_left[24] ;
 wire \ces_6_4_io_ins_left[25] ;
 wire \ces_6_4_io_ins_left[26] ;
 wire \ces_6_4_io_ins_left[27] ;
 wire \ces_6_4_io_ins_left[28] ;
 wire \ces_6_4_io_ins_left[29] ;
 wire \ces_6_4_io_ins_left[2] ;
 wire \ces_6_4_io_ins_left[30] ;
 wire \ces_6_4_io_ins_left[31] ;
 wire \ces_6_4_io_ins_left[32] ;
 wire \ces_6_4_io_ins_left[33] ;
 wire \ces_6_4_io_ins_left[34] ;
 wire \ces_6_4_io_ins_left[35] ;
 wire \ces_6_4_io_ins_left[36] ;
 wire \ces_6_4_io_ins_left[37] ;
 wire \ces_6_4_io_ins_left[38] ;
 wire \ces_6_4_io_ins_left[39] ;
 wire \ces_6_4_io_ins_left[3] ;
 wire \ces_6_4_io_ins_left[40] ;
 wire \ces_6_4_io_ins_left[41] ;
 wire \ces_6_4_io_ins_left[42] ;
 wire \ces_6_4_io_ins_left[43] ;
 wire \ces_6_4_io_ins_left[44] ;
 wire \ces_6_4_io_ins_left[45] ;
 wire \ces_6_4_io_ins_left[46] ;
 wire \ces_6_4_io_ins_left[47] ;
 wire \ces_6_4_io_ins_left[48] ;
 wire \ces_6_4_io_ins_left[49] ;
 wire \ces_6_4_io_ins_left[4] ;
 wire \ces_6_4_io_ins_left[50] ;
 wire \ces_6_4_io_ins_left[51] ;
 wire \ces_6_4_io_ins_left[52] ;
 wire \ces_6_4_io_ins_left[53] ;
 wire \ces_6_4_io_ins_left[54] ;
 wire \ces_6_4_io_ins_left[55] ;
 wire \ces_6_4_io_ins_left[56] ;
 wire \ces_6_4_io_ins_left[57] ;
 wire \ces_6_4_io_ins_left[58] ;
 wire \ces_6_4_io_ins_left[59] ;
 wire \ces_6_4_io_ins_left[5] ;
 wire \ces_6_4_io_ins_left[60] ;
 wire \ces_6_4_io_ins_left[61] ;
 wire \ces_6_4_io_ins_left[62] ;
 wire \ces_6_4_io_ins_left[63] ;
 wire \ces_6_4_io_ins_left[6] ;
 wire \ces_6_4_io_ins_left[7] ;
 wire \ces_6_4_io_ins_left[8] ;
 wire \ces_6_4_io_ins_left[9] ;
 wire ces_6_4_io_lsbOuts_0;
 wire ces_6_4_io_lsbOuts_1;
 wire ces_6_4_io_lsbOuts_2;
 wire ces_6_4_io_lsbOuts_3;
 wire ces_6_4_io_lsbOuts_4;
 wire ces_6_4_io_lsbOuts_5;
 wire ces_6_4_io_lsbOuts_6;
 wire ces_6_4_io_lsbOuts_7;
 wire \ces_6_4_io_outs_right[0] ;
 wire \ces_6_4_io_outs_right[10] ;
 wire \ces_6_4_io_outs_right[11] ;
 wire \ces_6_4_io_outs_right[12] ;
 wire \ces_6_4_io_outs_right[13] ;
 wire \ces_6_4_io_outs_right[14] ;
 wire \ces_6_4_io_outs_right[15] ;
 wire \ces_6_4_io_outs_right[16] ;
 wire \ces_6_4_io_outs_right[17] ;
 wire \ces_6_4_io_outs_right[18] ;
 wire \ces_6_4_io_outs_right[19] ;
 wire \ces_6_4_io_outs_right[1] ;
 wire \ces_6_4_io_outs_right[20] ;
 wire \ces_6_4_io_outs_right[21] ;
 wire \ces_6_4_io_outs_right[22] ;
 wire \ces_6_4_io_outs_right[23] ;
 wire \ces_6_4_io_outs_right[24] ;
 wire \ces_6_4_io_outs_right[25] ;
 wire \ces_6_4_io_outs_right[26] ;
 wire \ces_6_4_io_outs_right[27] ;
 wire \ces_6_4_io_outs_right[28] ;
 wire \ces_6_4_io_outs_right[29] ;
 wire \ces_6_4_io_outs_right[2] ;
 wire \ces_6_4_io_outs_right[30] ;
 wire \ces_6_4_io_outs_right[31] ;
 wire \ces_6_4_io_outs_right[32] ;
 wire \ces_6_4_io_outs_right[33] ;
 wire \ces_6_4_io_outs_right[34] ;
 wire \ces_6_4_io_outs_right[35] ;
 wire \ces_6_4_io_outs_right[36] ;
 wire \ces_6_4_io_outs_right[37] ;
 wire \ces_6_4_io_outs_right[38] ;
 wire \ces_6_4_io_outs_right[39] ;
 wire \ces_6_4_io_outs_right[3] ;
 wire \ces_6_4_io_outs_right[40] ;
 wire \ces_6_4_io_outs_right[41] ;
 wire \ces_6_4_io_outs_right[42] ;
 wire \ces_6_4_io_outs_right[43] ;
 wire \ces_6_4_io_outs_right[44] ;
 wire \ces_6_4_io_outs_right[45] ;
 wire \ces_6_4_io_outs_right[46] ;
 wire \ces_6_4_io_outs_right[47] ;
 wire \ces_6_4_io_outs_right[48] ;
 wire \ces_6_4_io_outs_right[49] ;
 wire \ces_6_4_io_outs_right[4] ;
 wire \ces_6_4_io_outs_right[50] ;
 wire \ces_6_4_io_outs_right[51] ;
 wire \ces_6_4_io_outs_right[52] ;
 wire \ces_6_4_io_outs_right[53] ;
 wire \ces_6_4_io_outs_right[54] ;
 wire \ces_6_4_io_outs_right[55] ;
 wire \ces_6_4_io_outs_right[56] ;
 wire \ces_6_4_io_outs_right[57] ;
 wire \ces_6_4_io_outs_right[58] ;
 wire \ces_6_4_io_outs_right[59] ;
 wire \ces_6_4_io_outs_right[5] ;
 wire \ces_6_4_io_outs_right[60] ;
 wire \ces_6_4_io_outs_right[61] ;
 wire \ces_6_4_io_outs_right[62] ;
 wire \ces_6_4_io_outs_right[63] ;
 wire \ces_6_4_io_outs_right[6] ;
 wire \ces_6_4_io_outs_right[7] ;
 wire \ces_6_4_io_outs_right[8] ;
 wire \ces_6_4_io_outs_right[9] ;
 wire \ces_6_4_io_outs_up[0] ;
 wire \ces_6_4_io_outs_up[10] ;
 wire \ces_6_4_io_outs_up[11] ;
 wire \ces_6_4_io_outs_up[12] ;
 wire \ces_6_4_io_outs_up[13] ;
 wire \ces_6_4_io_outs_up[14] ;
 wire \ces_6_4_io_outs_up[15] ;
 wire \ces_6_4_io_outs_up[16] ;
 wire \ces_6_4_io_outs_up[17] ;
 wire \ces_6_4_io_outs_up[18] ;
 wire \ces_6_4_io_outs_up[19] ;
 wire \ces_6_4_io_outs_up[1] ;
 wire \ces_6_4_io_outs_up[20] ;
 wire \ces_6_4_io_outs_up[21] ;
 wire \ces_6_4_io_outs_up[22] ;
 wire \ces_6_4_io_outs_up[23] ;
 wire \ces_6_4_io_outs_up[24] ;
 wire \ces_6_4_io_outs_up[25] ;
 wire \ces_6_4_io_outs_up[26] ;
 wire \ces_6_4_io_outs_up[27] ;
 wire \ces_6_4_io_outs_up[28] ;
 wire \ces_6_4_io_outs_up[29] ;
 wire \ces_6_4_io_outs_up[2] ;
 wire \ces_6_4_io_outs_up[30] ;
 wire \ces_6_4_io_outs_up[31] ;
 wire \ces_6_4_io_outs_up[32] ;
 wire \ces_6_4_io_outs_up[33] ;
 wire \ces_6_4_io_outs_up[34] ;
 wire \ces_6_4_io_outs_up[35] ;
 wire \ces_6_4_io_outs_up[36] ;
 wire \ces_6_4_io_outs_up[37] ;
 wire \ces_6_4_io_outs_up[38] ;
 wire \ces_6_4_io_outs_up[39] ;
 wire \ces_6_4_io_outs_up[3] ;
 wire \ces_6_4_io_outs_up[40] ;
 wire \ces_6_4_io_outs_up[41] ;
 wire \ces_6_4_io_outs_up[42] ;
 wire \ces_6_4_io_outs_up[43] ;
 wire \ces_6_4_io_outs_up[44] ;
 wire \ces_6_4_io_outs_up[45] ;
 wire \ces_6_4_io_outs_up[46] ;
 wire \ces_6_4_io_outs_up[47] ;
 wire \ces_6_4_io_outs_up[48] ;
 wire \ces_6_4_io_outs_up[49] ;
 wire \ces_6_4_io_outs_up[4] ;
 wire \ces_6_4_io_outs_up[50] ;
 wire \ces_6_4_io_outs_up[51] ;
 wire \ces_6_4_io_outs_up[52] ;
 wire \ces_6_4_io_outs_up[53] ;
 wire \ces_6_4_io_outs_up[54] ;
 wire \ces_6_4_io_outs_up[55] ;
 wire \ces_6_4_io_outs_up[56] ;
 wire \ces_6_4_io_outs_up[57] ;
 wire \ces_6_4_io_outs_up[58] ;
 wire \ces_6_4_io_outs_up[59] ;
 wire \ces_6_4_io_outs_up[5] ;
 wire \ces_6_4_io_outs_up[60] ;
 wire \ces_6_4_io_outs_up[61] ;
 wire \ces_6_4_io_outs_up[62] ;
 wire \ces_6_4_io_outs_up[63] ;
 wire \ces_6_4_io_outs_up[6] ;
 wire \ces_6_4_io_outs_up[7] ;
 wire \ces_6_4_io_outs_up[8] ;
 wire \ces_6_4_io_outs_up[9] ;
 wire \ces_6_5_io_ins_down[0] ;
 wire \ces_6_5_io_ins_down[10] ;
 wire \ces_6_5_io_ins_down[11] ;
 wire \ces_6_5_io_ins_down[12] ;
 wire \ces_6_5_io_ins_down[13] ;
 wire \ces_6_5_io_ins_down[14] ;
 wire \ces_6_5_io_ins_down[15] ;
 wire \ces_6_5_io_ins_down[16] ;
 wire \ces_6_5_io_ins_down[17] ;
 wire \ces_6_5_io_ins_down[18] ;
 wire \ces_6_5_io_ins_down[19] ;
 wire \ces_6_5_io_ins_down[1] ;
 wire \ces_6_5_io_ins_down[20] ;
 wire \ces_6_5_io_ins_down[21] ;
 wire \ces_6_5_io_ins_down[22] ;
 wire \ces_6_5_io_ins_down[23] ;
 wire \ces_6_5_io_ins_down[24] ;
 wire \ces_6_5_io_ins_down[25] ;
 wire \ces_6_5_io_ins_down[26] ;
 wire \ces_6_5_io_ins_down[27] ;
 wire \ces_6_5_io_ins_down[28] ;
 wire \ces_6_5_io_ins_down[29] ;
 wire \ces_6_5_io_ins_down[2] ;
 wire \ces_6_5_io_ins_down[30] ;
 wire \ces_6_5_io_ins_down[31] ;
 wire \ces_6_5_io_ins_down[32] ;
 wire \ces_6_5_io_ins_down[33] ;
 wire \ces_6_5_io_ins_down[34] ;
 wire \ces_6_5_io_ins_down[35] ;
 wire \ces_6_5_io_ins_down[36] ;
 wire \ces_6_5_io_ins_down[37] ;
 wire \ces_6_5_io_ins_down[38] ;
 wire \ces_6_5_io_ins_down[39] ;
 wire \ces_6_5_io_ins_down[3] ;
 wire \ces_6_5_io_ins_down[40] ;
 wire \ces_6_5_io_ins_down[41] ;
 wire \ces_6_5_io_ins_down[42] ;
 wire \ces_6_5_io_ins_down[43] ;
 wire \ces_6_5_io_ins_down[44] ;
 wire \ces_6_5_io_ins_down[45] ;
 wire \ces_6_5_io_ins_down[46] ;
 wire \ces_6_5_io_ins_down[47] ;
 wire \ces_6_5_io_ins_down[48] ;
 wire \ces_6_5_io_ins_down[49] ;
 wire \ces_6_5_io_ins_down[4] ;
 wire \ces_6_5_io_ins_down[50] ;
 wire \ces_6_5_io_ins_down[51] ;
 wire \ces_6_5_io_ins_down[52] ;
 wire \ces_6_5_io_ins_down[53] ;
 wire \ces_6_5_io_ins_down[54] ;
 wire \ces_6_5_io_ins_down[55] ;
 wire \ces_6_5_io_ins_down[56] ;
 wire \ces_6_5_io_ins_down[57] ;
 wire \ces_6_5_io_ins_down[58] ;
 wire \ces_6_5_io_ins_down[59] ;
 wire \ces_6_5_io_ins_down[5] ;
 wire \ces_6_5_io_ins_down[60] ;
 wire \ces_6_5_io_ins_down[61] ;
 wire \ces_6_5_io_ins_down[62] ;
 wire \ces_6_5_io_ins_down[63] ;
 wire \ces_6_5_io_ins_down[6] ;
 wire \ces_6_5_io_ins_down[7] ;
 wire \ces_6_5_io_ins_down[8] ;
 wire \ces_6_5_io_ins_down[9] ;
 wire \ces_6_5_io_ins_left[0] ;
 wire \ces_6_5_io_ins_left[10] ;
 wire \ces_6_5_io_ins_left[11] ;
 wire \ces_6_5_io_ins_left[12] ;
 wire \ces_6_5_io_ins_left[13] ;
 wire \ces_6_5_io_ins_left[14] ;
 wire \ces_6_5_io_ins_left[15] ;
 wire \ces_6_5_io_ins_left[16] ;
 wire \ces_6_5_io_ins_left[17] ;
 wire \ces_6_5_io_ins_left[18] ;
 wire \ces_6_5_io_ins_left[19] ;
 wire \ces_6_5_io_ins_left[1] ;
 wire \ces_6_5_io_ins_left[20] ;
 wire \ces_6_5_io_ins_left[21] ;
 wire \ces_6_5_io_ins_left[22] ;
 wire \ces_6_5_io_ins_left[23] ;
 wire \ces_6_5_io_ins_left[24] ;
 wire \ces_6_5_io_ins_left[25] ;
 wire \ces_6_5_io_ins_left[26] ;
 wire \ces_6_5_io_ins_left[27] ;
 wire \ces_6_5_io_ins_left[28] ;
 wire \ces_6_5_io_ins_left[29] ;
 wire \ces_6_5_io_ins_left[2] ;
 wire \ces_6_5_io_ins_left[30] ;
 wire \ces_6_5_io_ins_left[31] ;
 wire \ces_6_5_io_ins_left[32] ;
 wire \ces_6_5_io_ins_left[33] ;
 wire \ces_6_5_io_ins_left[34] ;
 wire \ces_6_5_io_ins_left[35] ;
 wire \ces_6_5_io_ins_left[36] ;
 wire \ces_6_5_io_ins_left[37] ;
 wire \ces_6_5_io_ins_left[38] ;
 wire \ces_6_5_io_ins_left[39] ;
 wire \ces_6_5_io_ins_left[3] ;
 wire \ces_6_5_io_ins_left[40] ;
 wire \ces_6_5_io_ins_left[41] ;
 wire \ces_6_5_io_ins_left[42] ;
 wire \ces_6_5_io_ins_left[43] ;
 wire \ces_6_5_io_ins_left[44] ;
 wire \ces_6_5_io_ins_left[45] ;
 wire \ces_6_5_io_ins_left[46] ;
 wire \ces_6_5_io_ins_left[47] ;
 wire \ces_6_5_io_ins_left[48] ;
 wire \ces_6_5_io_ins_left[49] ;
 wire \ces_6_5_io_ins_left[4] ;
 wire \ces_6_5_io_ins_left[50] ;
 wire \ces_6_5_io_ins_left[51] ;
 wire \ces_6_5_io_ins_left[52] ;
 wire \ces_6_5_io_ins_left[53] ;
 wire \ces_6_5_io_ins_left[54] ;
 wire \ces_6_5_io_ins_left[55] ;
 wire \ces_6_5_io_ins_left[56] ;
 wire \ces_6_5_io_ins_left[57] ;
 wire \ces_6_5_io_ins_left[58] ;
 wire \ces_6_5_io_ins_left[59] ;
 wire \ces_6_5_io_ins_left[5] ;
 wire \ces_6_5_io_ins_left[60] ;
 wire \ces_6_5_io_ins_left[61] ;
 wire \ces_6_5_io_ins_left[62] ;
 wire \ces_6_5_io_ins_left[63] ;
 wire \ces_6_5_io_ins_left[6] ;
 wire \ces_6_5_io_ins_left[7] ;
 wire \ces_6_5_io_ins_left[8] ;
 wire \ces_6_5_io_ins_left[9] ;
 wire ces_6_5_io_lsbOuts_0;
 wire ces_6_5_io_lsbOuts_1;
 wire ces_6_5_io_lsbOuts_2;
 wire ces_6_5_io_lsbOuts_3;
 wire ces_6_5_io_lsbOuts_4;
 wire ces_6_5_io_lsbOuts_5;
 wire ces_6_5_io_lsbOuts_6;
 wire ces_6_5_io_lsbOuts_7;
 wire \ces_6_5_io_outs_right[0] ;
 wire \ces_6_5_io_outs_right[10] ;
 wire \ces_6_5_io_outs_right[11] ;
 wire \ces_6_5_io_outs_right[12] ;
 wire \ces_6_5_io_outs_right[13] ;
 wire \ces_6_5_io_outs_right[14] ;
 wire \ces_6_5_io_outs_right[15] ;
 wire \ces_6_5_io_outs_right[16] ;
 wire \ces_6_5_io_outs_right[17] ;
 wire \ces_6_5_io_outs_right[18] ;
 wire \ces_6_5_io_outs_right[19] ;
 wire \ces_6_5_io_outs_right[1] ;
 wire \ces_6_5_io_outs_right[20] ;
 wire \ces_6_5_io_outs_right[21] ;
 wire \ces_6_5_io_outs_right[22] ;
 wire \ces_6_5_io_outs_right[23] ;
 wire \ces_6_5_io_outs_right[24] ;
 wire \ces_6_5_io_outs_right[25] ;
 wire \ces_6_5_io_outs_right[26] ;
 wire \ces_6_5_io_outs_right[27] ;
 wire \ces_6_5_io_outs_right[28] ;
 wire \ces_6_5_io_outs_right[29] ;
 wire \ces_6_5_io_outs_right[2] ;
 wire \ces_6_5_io_outs_right[30] ;
 wire \ces_6_5_io_outs_right[31] ;
 wire \ces_6_5_io_outs_right[32] ;
 wire \ces_6_5_io_outs_right[33] ;
 wire \ces_6_5_io_outs_right[34] ;
 wire \ces_6_5_io_outs_right[35] ;
 wire \ces_6_5_io_outs_right[36] ;
 wire \ces_6_5_io_outs_right[37] ;
 wire \ces_6_5_io_outs_right[38] ;
 wire \ces_6_5_io_outs_right[39] ;
 wire \ces_6_5_io_outs_right[3] ;
 wire \ces_6_5_io_outs_right[40] ;
 wire \ces_6_5_io_outs_right[41] ;
 wire \ces_6_5_io_outs_right[42] ;
 wire \ces_6_5_io_outs_right[43] ;
 wire \ces_6_5_io_outs_right[44] ;
 wire \ces_6_5_io_outs_right[45] ;
 wire \ces_6_5_io_outs_right[46] ;
 wire \ces_6_5_io_outs_right[47] ;
 wire \ces_6_5_io_outs_right[48] ;
 wire \ces_6_5_io_outs_right[49] ;
 wire \ces_6_5_io_outs_right[4] ;
 wire \ces_6_5_io_outs_right[50] ;
 wire \ces_6_5_io_outs_right[51] ;
 wire \ces_6_5_io_outs_right[52] ;
 wire \ces_6_5_io_outs_right[53] ;
 wire \ces_6_5_io_outs_right[54] ;
 wire \ces_6_5_io_outs_right[55] ;
 wire \ces_6_5_io_outs_right[56] ;
 wire \ces_6_5_io_outs_right[57] ;
 wire \ces_6_5_io_outs_right[58] ;
 wire \ces_6_5_io_outs_right[59] ;
 wire \ces_6_5_io_outs_right[5] ;
 wire \ces_6_5_io_outs_right[60] ;
 wire \ces_6_5_io_outs_right[61] ;
 wire \ces_6_5_io_outs_right[62] ;
 wire \ces_6_5_io_outs_right[63] ;
 wire \ces_6_5_io_outs_right[6] ;
 wire \ces_6_5_io_outs_right[7] ;
 wire \ces_6_5_io_outs_right[8] ;
 wire \ces_6_5_io_outs_right[9] ;
 wire \ces_6_5_io_outs_up[0] ;
 wire \ces_6_5_io_outs_up[10] ;
 wire \ces_6_5_io_outs_up[11] ;
 wire \ces_6_5_io_outs_up[12] ;
 wire \ces_6_5_io_outs_up[13] ;
 wire \ces_6_5_io_outs_up[14] ;
 wire \ces_6_5_io_outs_up[15] ;
 wire \ces_6_5_io_outs_up[16] ;
 wire \ces_6_5_io_outs_up[17] ;
 wire \ces_6_5_io_outs_up[18] ;
 wire \ces_6_5_io_outs_up[19] ;
 wire \ces_6_5_io_outs_up[1] ;
 wire \ces_6_5_io_outs_up[20] ;
 wire \ces_6_5_io_outs_up[21] ;
 wire \ces_6_5_io_outs_up[22] ;
 wire \ces_6_5_io_outs_up[23] ;
 wire \ces_6_5_io_outs_up[24] ;
 wire \ces_6_5_io_outs_up[25] ;
 wire \ces_6_5_io_outs_up[26] ;
 wire \ces_6_5_io_outs_up[27] ;
 wire \ces_6_5_io_outs_up[28] ;
 wire \ces_6_5_io_outs_up[29] ;
 wire \ces_6_5_io_outs_up[2] ;
 wire \ces_6_5_io_outs_up[30] ;
 wire \ces_6_5_io_outs_up[31] ;
 wire \ces_6_5_io_outs_up[32] ;
 wire \ces_6_5_io_outs_up[33] ;
 wire \ces_6_5_io_outs_up[34] ;
 wire \ces_6_5_io_outs_up[35] ;
 wire \ces_6_5_io_outs_up[36] ;
 wire \ces_6_5_io_outs_up[37] ;
 wire \ces_6_5_io_outs_up[38] ;
 wire \ces_6_5_io_outs_up[39] ;
 wire \ces_6_5_io_outs_up[3] ;
 wire \ces_6_5_io_outs_up[40] ;
 wire \ces_6_5_io_outs_up[41] ;
 wire \ces_6_5_io_outs_up[42] ;
 wire \ces_6_5_io_outs_up[43] ;
 wire \ces_6_5_io_outs_up[44] ;
 wire \ces_6_5_io_outs_up[45] ;
 wire \ces_6_5_io_outs_up[46] ;
 wire \ces_6_5_io_outs_up[47] ;
 wire \ces_6_5_io_outs_up[48] ;
 wire \ces_6_5_io_outs_up[49] ;
 wire \ces_6_5_io_outs_up[4] ;
 wire \ces_6_5_io_outs_up[50] ;
 wire \ces_6_5_io_outs_up[51] ;
 wire \ces_6_5_io_outs_up[52] ;
 wire \ces_6_5_io_outs_up[53] ;
 wire \ces_6_5_io_outs_up[54] ;
 wire \ces_6_5_io_outs_up[55] ;
 wire \ces_6_5_io_outs_up[56] ;
 wire \ces_6_5_io_outs_up[57] ;
 wire \ces_6_5_io_outs_up[58] ;
 wire \ces_6_5_io_outs_up[59] ;
 wire \ces_6_5_io_outs_up[5] ;
 wire \ces_6_5_io_outs_up[60] ;
 wire \ces_6_5_io_outs_up[61] ;
 wire \ces_6_5_io_outs_up[62] ;
 wire \ces_6_5_io_outs_up[63] ;
 wire \ces_6_5_io_outs_up[6] ;
 wire \ces_6_5_io_outs_up[7] ;
 wire \ces_6_5_io_outs_up[8] ;
 wire \ces_6_5_io_outs_up[9] ;
 wire \ces_6_6_io_ins_down[0] ;
 wire \ces_6_6_io_ins_down[10] ;
 wire \ces_6_6_io_ins_down[11] ;
 wire \ces_6_6_io_ins_down[12] ;
 wire \ces_6_6_io_ins_down[13] ;
 wire \ces_6_6_io_ins_down[14] ;
 wire \ces_6_6_io_ins_down[15] ;
 wire \ces_6_6_io_ins_down[16] ;
 wire \ces_6_6_io_ins_down[17] ;
 wire \ces_6_6_io_ins_down[18] ;
 wire \ces_6_6_io_ins_down[19] ;
 wire \ces_6_6_io_ins_down[1] ;
 wire \ces_6_6_io_ins_down[20] ;
 wire \ces_6_6_io_ins_down[21] ;
 wire \ces_6_6_io_ins_down[22] ;
 wire \ces_6_6_io_ins_down[23] ;
 wire \ces_6_6_io_ins_down[24] ;
 wire \ces_6_6_io_ins_down[25] ;
 wire \ces_6_6_io_ins_down[26] ;
 wire \ces_6_6_io_ins_down[27] ;
 wire \ces_6_6_io_ins_down[28] ;
 wire \ces_6_6_io_ins_down[29] ;
 wire \ces_6_6_io_ins_down[2] ;
 wire \ces_6_6_io_ins_down[30] ;
 wire \ces_6_6_io_ins_down[31] ;
 wire \ces_6_6_io_ins_down[32] ;
 wire \ces_6_6_io_ins_down[33] ;
 wire \ces_6_6_io_ins_down[34] ;
 wire \ces_6_6_io_ins_down[35] ;
 wire \ces_6_6_io_ins_down[36] ;
 wire \ces_6_6_io_ins_down[37] ;
 wire \ces_6_6_io_ins_down[38] ;
 wire \ces_6_6_io_ins_down[39] ;
 wire \ces_6_6_io_ins_down[3] ;
 wire \ces_6_6_io_ins_down[40] ;
 wire \ces_6_6_io_ins_down[41] ;
 wire \ces_6_6_io_ins_down[42] ;
 wire \ces_6_6_io_ins_down[43] ;
 wire \ces_6_6_io_ins_down[44] ;
 wire \ces_6_6_io_ins_down[45] ;
 wire \ces_6_6_io_ins_down[46] ;
 wire \ces_6_6_io_ins_down[47] ;
 wire \ces_6_6_io_ins_down[48] ;
 wire \ces_6_6_io_ins_down[49] ;
 wire \ces_6_6_io_ins_down[4] ;
 wire \ces_6_6_io_ins_down[50] ;
 wire \ces_6_6_io_ins_down[51] ;
 wire \ces_6_6_io_ins_down[52] ;
 wire \ces_6_6_io_ins_down[53] ;
 wire \ces_6_6_io_ins_down[54] ;
 wire \ces_6_6_io_ins_down[55] ;
 wire \ces_6_6_io_ins_down[56] ;
 wire \ces_6_6_io_ins_down[57] ;
 wire \ces_6_6_io_ins_down[58] ;
 wire \ces_6_6_io_ins_down[59] ;
 wire \ces_6_6_io_ins_down[5] ;
 wire \ces_6_6_io_ins_down[60] ;
 wire \ces_6_6_io_ins_down[61] ;
 wire \ces_6_6_io_ins_down[62] ;
 wire \ces_6_6_io_ins_down[63] ;
 wire \ces_6_6_io_ins_down[6] ;
 wire \ces_6_6_io_ins_down[7] ;
 wire \ces_6_6_io_ins_down[8] ;
 wire \ces_6_6_io_ins_down[9] ;
 wire \ces_6_6_io_ins_left[0] ;
 wire \ces_6_6_io_ins_left[10] ;
 wire \ces_6_6_io_ins_left[11] ;
 wire \ces_6_6_io_ins_left[12] ;
 wire \ces_6_6_io_ins_left[13] ;
 wire \ces_6_6_io_ins_left[14] ;
 wire \ces_6_6_io_ins_left[15] ;
 wire \ces_6_6_io_ins_left[16] ;
 wire \ces_6_6_io_ins_left[17] ;
 wire \ces_6_6_io_ins_left[18] ;
 wire \ces_6_6_io_ins_left[19] ;
 wire \ces_6_6_io_ins_left[1] ;
 wire \ces_6_6_io_ins_left[20] ;
 wire \ces_6_6_io_ins_left[21] ;
 wire \ces_6_6_io_ins_left[22] ;
 wire \ces_6_6_io_ins_left[23] ;
 wire \ces_6_6_io_ins_left[24] ;
 wire \ces_6_6_io_ins_left[25] ;
 wire \ces_6_6_io_ins_left[26] ;
 wire \ces_6_6_io_ins_left[27] ;
 wire \ces_6_6_io_ins_left[28] ;
 wire \ces_6_6_io_ins_left[29] ;
 wire \ces_6_6_io_ins_left[2] ;
 wire \ces_6_6_io_ins_left[30] ;
 wire \ces_6_6_io_ins_left[31] ;
 wire \ces_6_6_io_ins_left[32] ;
 wire \ces_6_6_io_ins_left[33] ;
 wire \ces_6_6_io_ins_left[34] ;
 wire \ces_6_6_io_ins_left[35] ;
 wire \ces_6_6_io_ins_left[36] ;
 wire \ces_6_6_io_ins_left[37] ;
 wire \ces_6_6_io_ins_left[38] ;
 wire \ces_6_6_io_ins_left[39] ;
 wire \ces_6_6_io_ins_left[3] ;
 wire \ces_6_6_io_ins_left[40] ;
 wire \ces_6_6_io_ins_left[41] ;
 wire \ces_6_6_io_ins_left[42] ;
 wire \ces_6_6_io_ins_left[43] ;
 wire \ces_6_6_io_ins_left[44] ;
 wire \ces_6_6_io_ins_left[45] ;
 wire \ces_6_6_io_ins_left[46] ;
 wire \ces_6_6_io_ins_left[47] ;
 wire \ces_6_6_io_ins_left[48] ;
 wire \ces_6_6_io_ins_left[49] ;
 wire \ces_6_6_io_ins_left[4] ;
 wire \ces_6_6_io_ins_left[50] ;
 wire \ces_6_6_io_ins_left[51] ;
 wire \ces_6_6_io_ins_left[52] ;
 wire \ces_6_6_io_ins_left[53] ;
 wire \ces_6_6_io_ins_left[54] ;
 wire \ces_6_6_io_ins_left[55] ;
 wire \ces_6_6_io_ins_left[56] ;
 wire \ces_6_6_io_ins_left[57] ;
 wire \ces_6_6_io_ins_left[58] ;
 wire \ces_6_6_io_ins_left[59] ;
 wire \ces_6_6_io_ins_left[5] ;
 wire \ces_6_6_io_ins_left[60] ;
 wire \ces_6_6_io_ins_left[61] ;
 wire \ces_6_6_io_ins_left[62] ;
 wire \ces_6_6_io_ins_left[63] ;
 wire \ces_6_6_io_ins_left[6] ;
 wire \ces_6_6_io_ins_left[7] ;
 wire \ces_6_6_io_ins_left[8] ;
 wire \ces_6_6_io_ins_left[9] ;
 wire ces_6_6_io_lsbOuts_0;
 wire ces_6_6_io_lsbOuts_1;
 wire ces_6_6_io_lsbOuts_2;
 wire ces_6_6_io_lsbOuts_3;
 wire ces_6_6_io_lsbOuts_4;
 wire ces_6_6_io_lsbOuts_5;
 wire ces_6_6_io_lsbOuts_6;
 wire ces_6_6_io_lsbOuts_7;
 wire \ces_6_6_io_outs_right[0] ;
 wire \ces_6_6_io_outs_right[10] ;
 wire \ces_6_6_io_outs_right[11] ;
 wire \ces_6_6_io_outs_right[12] ;
 wire \ces_6_6_io_outs_right[13] ;
 wire \ces_6_6_io_outs_right[14] ;
 wire \ces_6_6_io_outs_right[15] ;
 wire \ces_6_6_io_outs_right[16] ;
 wire \ces_6_6_io_outs_right[17] ;
 wire \ces_6_6_io_outs_right[18] ;
 wire \ces_6_6_io_outs_right[19] ;
 wire \ces_6_6_io_outs_right[1] ;
 wire \ces_6_6_io_outs_right[20] ;
 wire \ces_6_6_io_outs_right[21] ;
 wire \ces_6_6_io_outs_right[22] ;
 wire \ces_6_6_io_outs_right[23] ;
 wire \ces_6_6_io_outs_right[24] ;
 wire \ces_6_6_io_outs_right[25] ;
 wire \ces_6_6_io_outs_right[26] ;
 wire \ces_6_6_io_outs_right[27] ;
 wire \ces_6_6_io_outs_right[28] ;
 wire \ces_6_6_io_outs_right[29] ;
 wire \ces_6_6_io_outs_right[2] ;
 wire \ces_6_6_io_outs_right[30] ;
 wire \ces_6_6_io_outs_right[31] ;
 wire \ces_6_6_io_outs_right[32] ;
 wire \ces_6_6_io_outs_right[33] ;
 wire \ces_6_6_io_outs_right[34] ;
 wire \ces_6_6_io_outs_right[35] ;
 wire \ces_6_6_io_outs_right[36] ;
 wire \ces_6_6_io_outs_right[37] ;
 wire \ces_6_6_io_outs_right[38] ;
 wire \ces_6_6_io_outs_right[39] ;
 wire \ces_6_6_io_outs_right[3] ;
 wire \ces_6_6_io_outs_right[40] ;
 wire \ces_6_6_io_outs_right[41] ;
 wire \ces_6_6_io_outs_right[42] ;
 wire \ces_6_6_io_outs_right[43] ;
 wire \ces_6_6_io_outs_right[44] ;
 wire \ces_6_6_io_outs_right[45] ;
 wire \ces_6_6_io_outs_right[46] ;
 wire \ces_6_6_io_outs_right[47] ;
 wire \ces_6_6_io_outs_right[48] ;
 wire \ces_6_6_io_outs_right[49] ;
 wire \ces_6_6_io_outs_right[4] ;
 wire \ces_6_6_io_outs_right[50] ;
 wire \ces_6_6_io_outs_right[51] ;
 wire \ces_6_6_io_outs_right[52] ;
 wire \ces_6_6_io_outs_right[53] ;
 wire \ces_6_6_io_outs_right[54] ;
 wire \ces_6_6_io_outs_right[55] ;
 wire \ces_6_6_io_outs_right[56] ;
 wire \ces_6_6_io_outs_right[57] ;
 wire \ces_6_6_io_outs_right[58] ;
 wire \ces_6_6_io_outs_right[59] ;
 wire \ces_6_6_io_outs_right[5] ;
 wire \ces_6_6_io_outs_right[60] ;
 wire \ces_6_6_io_outs_right[61] ;
 wire \ces_6_6_io_outs_right[62] ;
 wire \ces_6_6_io_outs_right[63] ;
 wire \ces_6_6_io_outs_right[6] ;
 wire \ces_6_6_io_outs_right[7] ;
 wire \ces_6_6_io_outs_right[8] ;
 wire \ces_6_6_io_outs_right[9] ;
 wire \ces_6_6_io_outs_up[0] ;
 wire \ces_6_6_io_outs_up[10] ;
 wire \ces_6_6_io_outs_up[11] ;
 wire \ces_6_6_io_outs_up[12] ;
 wire \ces_6_6_io_outs_up[13] ;
 wire \ces_6_6_io_outs_up[14] ;
 wire \ces_6_6_io_outs_up[15] ;
 wire \ces_6_6_io_outs_up[16] ;
 wire \ces_6_6_io_outs_up[17] ;
 wire \ces_6_6_io_outs_up[18] ;
 wire \ces_6_6_io_outs_up[19] ;
 wire \ces_6_6_io_outs_up[1] ;
 wire \ces_6_6_io_outs_up[20] ;
 wire \ces_6_6_io_outs_up[21] ;
 wire \ces_6_6_io_outs_up[22] ;
 wire \ces_6_6_io_outs_up[23] ;
 wire \ces_6_6_io_outs_up[24] ;
 wire \ces_6_6_io_outs_up[25] ;
 wire \ces_6_6_io_outs_up[26] ;
 wire \ces_6_6_io_outs_up[27] ;
 wire \ces_6_6_io_outs_up[28] ;
 wire \ces_6_6_io_outs_up[29] ;
 wire \ces_6_6_io_outs_up[2] ;
 wire \ces_6_6_io_outs_up[30] ;
 wire \ces_6_6_io_outs_up[31] ;
 wire \ces_6_6_io_outs_up[32] ;
 wire \ces_6_6_io_outs_up[33] ;
 wire \ces_6_6_io_outs_up[34] ;
 wire \ces_6_6_io_outs_up[35] ;
 wire \ces_6_6_io_outs_up[36] ;
 wire \ces_6_6_io_outs_up[37] ;
 wire \ces_6_6_io_outs_up[38] ;
 wire \ces_6_6_io_outs_up[39] ;
 wire \ces_6_6_io_outs_up[3] ;
 wire \ces_6_6_io_outs_up[40] ;
 wire \ces_6_6_io_outs_up[41] ;
 wire \ces_6_6_io_outs_up[42] ;
 wire \ces_6_6_io_outs_up[43] ;
 wire \ces_6_6_io_outs_up[44] ;
 wire \ces_6_6_io_outs_up[45] ;
 wire \ces_6_6_io_outs_up[46] ;
 wire \ces_6_6_io_outs_up[47] ;
 wire \ces_6_6_io_outs_up[48] ;
 wire \ces_6_6_io_outs_up[49] ;
 wire \ces_6_6_io_outs_up[4] ;
 wire \ces_6_6_io_outs_up[50] ;
 wire \ces_6_6_io_outs_up[51] ;
 wire \ces_6_6_io_outs_up[52] ;
 wire \ces_6_6_io_outs_up[53] ;
 wire \ces_6_6_io_outs_up[54] ;
 wire \ces_6_6_io_outs_up[55] ;
 wire \ces_6_6_io_outs_up[56] ;
 wire \ces_6_6_io_outs_up[57] ;
 wire \ces_6_6_io_outs_up[58] ;
 wire \ces_6_6_io_outs_up[59] ;
 wire \ces_6_6_io_outs_up[5] ;
 wire \ces_6_6_io_outs_up[60] ;
 wire \ces_6_6_io_outs_up[61] ;
 wire \ces_6_6_io_outs_up[62] ;
 wire \ces_6_6_io_outs_up[63] ;
 wire \ces_6_6_io_outs_up[6] ;
 wire \ces_6_6_io_outs_up[7] ;
 wire \ces_6_6_io_outs_up[8] ;
 wire \ces_6_6_io_outs_up[9] ;
 wire \ces_6_7_io_ins_down[0] ;
 wire \ces_6_7_io_ins_down[10] ;
 wire \ces_6_7_io_ins_down[11] ;
 wire \ces_6_7_io_ins_down[12] ;
 wire \ces_6_7_io_ins_down[13] ;
 wire \ces_6_7_io_ins_down[14] ;
 wire \ces_6_7_io_ins_down[15] ;
 wire \ces_6_7_io_ins_down[16] ;
 wire \ces_6_7_io_ins_down[17] ;
 wire \ces_6_7_io_ins_down[18] ;
 wire \ces_6_7_io_ins_down[19] ;
 wire \ces_6_7_io_ins_down[1] ;
 wire \ces_6_7_io_ins_down[20] ;
 wire \ces_6_7_io_ins_down[21] ;
 wire \ces_6_7_io_ins_down[22] ;
 wire \ces_6_7_io_ins_down[23] ;
 wire \ces_6_7_io_ins_down[24] ;
 wire \ces_6_7_io_ins_down[25] ;
 wire \ces_6_7_io_ins_down[26] ;
 wire \ces_6_7_io_ins_down[27] ;
 wire \ces_6_7_io_ins_down[28] ;
 wire \ces_6_7_io_ins_down[29] ;
 wire \ces_6_7_io_ins_down[2] ;
 wire \ces_6_7_io_ins_down[30] ;
 wire \ces_6_7_io_ins_down[31] ;
 wire \ces_6_7_io_ins_down[32] ;
 wire \ces_6_7_io_ins_down[33] ;
 wire \ces_6_7_io_ins_down[34] ;
 wire \ces_6_7_io_ins_down[35] ;
 wire \ces_6_7_io_ins_down[36] ;
 wire \ces_6_7_io_ins_down[37] ;
 wire \ces_6_7_io_ins_down[38] ;
 wire \ces_6_7_io_ins_down[39] ;
 wire \ces_6_7_io_ins_down[3] ;
 wire \ces_6_7_io_ins_down[40] ;
 wire \ces_6_7_io_ins_down[41] ;
 wire \ces_6_7_io_ins_down[42] ;
 wire \ces_6_7_io_ins_down[43] ;
 wire \ces_6_7_io_ins_down[44] ;
 wire \ces_6_7_io_ins_down[45] ;
 wire \ces_6_7_io_ins_down[46] ;
 wire \ces_6_7_io_ins_down[47] ;
 wire \ces_6_7_io_ins_down[48] ;
 wire \ces_6_7_io_ins_down[49] ;
 wire \ces_6_7_io_ins_down[4] ;
 wire \ces_6_7_io_ins_down[50] ;
 wire \ces_6_7_io_ins_down[51] ;
 wire \ces_6_7_io_ins_down[52] ;
 wire \ces_6_7_io_ins_down[53] ;
 wire \ces_6_7_io_ins_down[54] ;
 wire \ces_6_7_io_ins_down[55] ;
 wire \ces_6_7_io_ins_down[56] ;
 wire \ces_6_7_io_ins_down[57] ;
 wire \ces_6_7_io_ins_down[58] ;
 wire \ces_6_7_io_ins_down[59] ;
 wire \ces_6_7_io_ins_down[5] ;
 wire \ces_6_7_io_ins_down[60] ;
 wire \ces_6_7_io_ins_down[61] ;
 wire \ces_6_7_io_ins_down[62] ;
 wire \ces_6_7_io_ins_down[63] ;
 wire \ces_6_7_io_ins_down[6] ;
 wire \ces_6_7_io_ins_down[7] ;
 wire \ces_6_7_io_ins_down[8] ;
 wire \ces_6_7_io_ins_down[9] ;
 wire ces_6_7_io_lsbOuts_0;
 wire ces_6_7_io_lsbOuts_1;
 wire ces_6_7_io_lsbOuts_2;
 wire ces_6_7_io_lsbOuts_3;
 wire ces_6_7_io_lsbOuts_4;
 wire ces_6_7_io_lsbOuts_5;
 wire ces_6_7_io_lsbOuts_6;
 wire ces_6_7_io_lsbOuts_7;
 wire \ces_6_7_io_outs_up[0] ;
 wire \ces_6_7_io_outs_up[10] ;
 wire \ces_6_7_io_outs_up[11] ;
 wire \ces_6_7_io_outs_up[12] ;
 wire \ces_6_7_io_outs_up[13] ;
 wire \ces_6_7_io_outs_up[14] ;
 wire \ces_6_7_io_outs_up[15] ;
 wire \ces_6_7_io_outs_up[16] ;
 wire \ces_6_7_io_outs_up[17] ;
 wire \ces_6_7_io_outs_up[18] ;
 wire \ces_6_7_io_outs_up[19] ;
 wire \ces_6_7_io_outs_up[1] ;
 wire \ces_6_7_io_outs_up[20] ;
 wire \ces_6_7_io_outs_up[21] ;
 wire \ces_6_7_io_outs_up[22] ;
 wire \ces_6_7_io_outs_up[23] ;
 wire \ces_6_7_io_outs_up[24] ;
 wire \ces_6_7_io_outs_up[25] ;
 wire \ces_6_7_io_outs_up[26] ;
 wire \ces_6_7_io_outs_up[27] ;
 wire \ces_6_7_io_outs_up[28] ;
 wire \ces_6_7_io_outs_up[29] ;
 wire \ces_6_7_io_outs_up[2] ;
 wire \ces_6_7_io_outs_up[30] ;
 wire \ces_6_7_io_outs_up[31] ;
 wire \ces_6_7_io_outs_up[32] ;
 wire \ces_6_7_io_outs_up[33] ;
 wire \ces_6_7_io_outs_up[34] ;
 wire \ces_6_7_io_outs_up[35] ;
 wire \ces_6_7_io_outs_up[36] ;
 wire \ces_6_7_io_outs_up[37] ;
 wire \ces_6_7_io_outs_up[38] ;
 wire \ces_6_7_io_outs_up[39] ;
 wire \ces_6_7_io_outs_up[3] ;
 wire \ces_6_7_io_outs_up[40] ;
 wire \ces_6_7_io_outs_up[41] ;
 wire \ces_6_7_io_outs_up[42] ;
 wire \ces_6_7_io_outs_up[43] ;
 wire \ces_6_7_io_outs_up[44] ;
 wire \ces_6_7_io_outs_up[45] ;
 wire \ces_6_7_io_outs_up[46] ;
 wire \ces_6_7_io_outs_up[47] ;
 wire \ces_6_7_io_outs_up[48] ;
 wire \ces_6_7_io_outs_up[49] ;
 wire \ces_6_7_io_outs_up[4] ;
 wire \ces_6_7_io_outs_up[50] ;
 wire \ces_6_7_io_outs_up[51] ;
 wire \ces_6_7_io_outs_up[52] ;
 wire \ces_6_7_io_outs_up[53] ;
 wire \ces_6_7_io_outs_up[54] ;
 wire \ces_6_7_io_outs_up[55] ;
 wire \ces_6_7_io_outs_up[56] ;
 wire \ces_6_7_io_outs_up[57] ;
 wire \ces_6_7_io_outs_up[58] ;
 wire \ces_6_7_io_outs_up[59] ;
 wire \ces_6_7_io_outs_up[5] ;
 wire \ces_6_7_io_outs_up[60] ;
 wire \ces_6_7_io_outs_up[61] ;
 wire \ces_6_7_io_outs_up[62] ;
 wire \ces_6_7_io_outs_up[63] ;
 wire \ces_6_7_io_outs_up[6] ;
 wire \ces_6_7_io_outs_up[7] ;
 wire \ces_6_7_io_outs_up[8] ;
 wire \ces_6_7_io_outs_up[9] ;
 wire \ces_7_0_io_ins_left[0] ;
 wire \ces_7_0_io_ins_left[10] ;
 wire \ces_7_0_io_ins_left[11] ;
 wire \ces_7_0_io_ins_left[12] ;
 wire \ces_7_0_io_ins_left[13] ;
 wire \ces_7_0_io_ins_left[14] ;
 wire \ces_7_0_io_ins_left[15] ;
 wire \ces_7_0_io_ins_left[16] ;
 wire \ces_7_0_io_ins_left[17] ;
 wire \ces_7_0_io_ins_left[18] ;
 wire \ces_7_0_io_ins_left[19] ;
 wire \ces_7_0_io_ins_left[1] ;
 wire \ces_7_0_io_ins_left[20] ;
 wire \ces_7_0_io_ins_left[21] ;
 wire \ces_7_0_io_ins_left[22] ;
 wire \ces_7_0_io_ins_left[23] ;
 wire \ces_7_0_io_ins_left[24] ;
 wire \ces_7_0_io_ins_left[25] ;
 wire \ces_7_0_io_ins_left[26] ;
 wire \ces_7_0_io_ins_left[27] ;
 wire \ces_7_0_io_ins_left[28] ;
 wire \ces_7_0_io_ins_left[29] ;
 wire \ces_7_0_io_ins_left[2] ;
 wire \ces_7_0_io_ins_left[30] ;
 wire \ces_7_0_io_ins_left[31] ;
 wire \ces_7_0_io_ins_left[32] ;
 wire \ces_7_0_io_ins_left[33] ;
 wire \ces_7_0_io_ins_left[34] ;
 wire \ces_7_0_io_ins_left[35] ;
 wire \ces_7_0_io_ins_left[36] ;
 wire \ces_7_0_io_ins_left[37] ;
 wire \ces_7_0_io_ins_left[38] ;
 wire \ces_7_0_io_ins_left[39] ;
 wire \ces_7_0_io_ins_left[3] ;
 wire \ces_7_0_io_ins_left[40] ;
 wire \ces_7_0_io_ins_left[41] ;
 wire \ces_7_0_io_ins_left[42] ;
 wire \ces_7_0_io_ins_left[43] ;
 wire \ces_7_0_io_ins_left[44] ;
 wire \ces_7_0_io_ins_left[45] ;
 wire \ces_7_0_io_ins_left[46] ;
 wire \ces_7_0_io_ins_left[47] ;
 wire \ces_7_0_io_ins_left[48] ;
 wire \ces_7_0_io_ins_left[49] ;
 wire \ces_7_0_io_ins_left[4] ;
 wire \ces_7_0_io_ins_left[50] ;
 wire \ces_7_0_io_ins_left[51] ;
 wire \ces_7_0_io_ins_left[52] ;
 wire \ces_7_0_io_ins_left[53] ;
 wire \ces_7_0_io_ins_left[54] ;
 wire \ces_7_0_io_ins_left[55] ;
 wire \ces_7_0_io_ins_left[56] ;
 wire \ces_7_0_io_ins_left[57] ;
 wire \ces_7_0_io_ins_left[58] ;
 wire \ces_7_0_io_ins_left[59] ;
 wire \ces_7_0_io_ins_left[5] ;
 wire \ces_7_0_io_ins_left[60] ;
 wire \ces_7_0_io_ins_left[61] ;
 wire \ces_7_0_io_ins_left[62] ;
 wire \ces_7_0_io_ins_left[63] ;
 wire \ces_7_0_io_ins_left[6] ;
 wire \ces_7_0_io_ins_left[7] ;
 wire \ces_7_0_io_ins_left[8] ;
 wire \ces_7_0_io_ins_left[9] ;
 wire ces_7_0_io_lsbOuts_0;
 wire ces_7_0_io_lsbOuts_1;
 wire ces_7_0_io_lsbOuts_2;
 wire ces_7_0_io_lsbOuts_3;
 wire ces_7_0_io_lsbOuts_4;
 wire ces_7_0_io_lsbOuts_5;
 wire ces_7_0_io_lsbOuts_6;
 wire ces_7_0_io_lsbOuts_7;
 wire \ces_7_0_io_outs_right[0] ;
 wire \ces_7_0_io_outs_right[10] ;
 wire \ces_7_0_io_outs_right[11] ;
 wire \ces_7_0_io_outs_right[12] ;
 wire \ces_7_0_io_outs_right[13] ;
 wire \ces_7_0_io_outs_right[14] ;
 wire \ces_7_0_io_outs_right[15] ;
 wire \ces_7_0_io_outs_right[16] ;
 wire \ces_7_0_io_outs_right[17] ;
 wire \ces_7_0_io_outs_right[18] ;
 wire \ces_7_0_io_outs_right[19] ;
 wire \ces_7_0_io_outs_right[1] ;
 wire \ces_7_0_io_outs_right[20] ;
 wire \ces_7_0_io_outs_right[21] ;
 wire \ces_7_0_io_outs_right[22] ;
 wire \ces_7_0_io_outs_right[23] ;
 wire \ces_7_0_io_outs_right[24] ;
 wire \ces_7_0_io_outs_right[25] ;
 wire \ces_7_0_io_outs_right[26] ;
 wire \ces_7_0_io_outs_right[27] ;
 wire \ces_7_0_io_outs_right[28] ;
 wire \ces_7_0_io_outs_right[29] ;
 wire \ces_7_0_io_outs_right[2] ;
 wire \ces_7_0_io_outs_right[30] ;
 wire \ces_7_0_io_outs_right[31] ;
 wire \ces_7_0_io_outs_right[32] ;
 wire \ces_7_0_io_outs_right[33] ;
 wire \ces_7_0_io_outs_right[34] ;
 wire \ces_7_0_io_outs_right[35] ;
 wire \ces_7_0_io_outs_right[36] ;
 wire \ces_7_0_io_outs_right[37] ;
 wire \ces_7_0_io_outs_right[38] ;
 wire \ces_7_0_io_outs_right[39] ;
 wire \ces_7_0_io_outs_right[3] ;
 wire \ces_7_0_io_outs_right[40] ;
 wire \ces_7_0_io_outs_right[41] ;
 wire \ces_7_0_io_outs_right[42] ;
 wire \ces_7_0_io_outs_right[43] ;
 wire \ces_7_0_io_outs_right[44] ;
 wire \ces_7_0_io_outs_right[45] ;
 wire \ces_7_0_io_outs_right[46] ;
 wire \ces_7_0_io_outs_right[47] ;
 wire \ces_7_0_io_outs_right[48] ;
 wire \ces_7_0_io_outs_right[49] ;
 wire \ces_7_0_io_outs_right[4] ;
 wire \ces_7_0_io_outs_right[50] ;
 wire \ces_7_0_io_outs_right[51] ;
 wire \ces_7_0_io_outs_right[52] ;
 wire \ces_7_0_io_outs_right[53] ;
 wire \ces_7_0_io_outs_right[54] ;
 wire \ces_7_0_io_outs_right[55] ;
 wire \ces_7_0_io_outs_right[56] ;
 wire \ces_7_0_io_outs_right[57] ;
 wire \ces_7_0_io_outs_right[58] ;
 wire \ces_7_0_io_outs_right[59] ;
 wire \ces_7_0_io_outs_right[5] ;
 wire \ces_7_0_io_outs_right[60] ;
 wire \ces_7_0_io_outs_right[61] ;
 wire \ces_7_0_io_outs_right[62] ;
 wire \ces_7_0_io_outs_right[63] ;
 wire \ces_7_0_io_outs_right[6] ;
 wire \ces_7_0_io_outs_right[7] ;
 wire \ces_7_0_io_outs_right[8] ;
 wire \ces_7_0_io_outs_right[9] ;
 wire \ces_7_1_io_ins_left[0] ;
 wire \ces_7_1_io_ins_left[10] ;
 wire \ces_7_1_io_ins_left[11] ;
 wire \ces_7_1_io_ins_left[12] ;
 wire \ces_7_1_io_ins_left[13] ;
 wire \ces_7_1_io_ins_left[14] ;
 wire \ces_7_1_io_ins_left[15] ;
 wire \ces_7_1_io_ins_left[16] ;
 wire \ces_7_1_io_ins_left[17] ;
 wire \ces_7_1_io_ins_left[18] ;
 wire \ces_7_1_io_ins_left[19] ;
 wire \ces_7_1_io_ins_left[1] ;
 wire \ces_7_1_io_ins_left[20] ;
 wire \ces_7_1_io_ins_left[21] ;
 wire \ces_7_1_io_ins_left[22] ;
 wire \ces_7_1_io_ins_left[23] ;
 wire \ces_7_1_io_ins_left[24] ;
 wire \ces_7_1_io_ins_left[25] ;
 wire \ces_7_1_io_ins_left[26] ;
 wire \ces_7_1_io_ins_left[27] ;
 wire \ces_7_1_io_ins_left[28] ;
 wire \ces_7_1_io_ins_left[29] ;
 wire \ces_7_1_io_ins_left[2] ;
 wire \ces_7_1_io_ins_left[30] ;
 wire \ces_7_1_io_ins_left[31] ;
 wire \ces_7_1_io_ins_left[32] ;
 wire \ces_7_1_io_ins_left[33] ;
 wire \ces_7_1_io_ins_left[34] ;
 wire \ces_7_1_io_ins_left[35] ;
 wire \ces_7_1_io_ins_left[36] ;
 wire \ces_7_1_io_ins_left[37] ;
 wire \ces_7_1_io_ins_left[38] ;
 wire \ces_7_1_io_ins_left[39] ;
 wire \ces_7_1_io_ins_left[3] ;
 wire \ces_7_1_io_ins_left[40] ;
 wire \ces_7_1_io_ins_left[41] ;
 wire \ces_7_1_io_ins_left[42] ;
 wire \ces_7_1_io_ins_left[43] ;
 wire \ces_7_1_io_ins_left[44] ;
 wire \ces_7_1_io_ins_left[45] ;
 wire \ces_7_1_io_ins_left[46] ;
 wire \ces_7_1_io_ins_left[47] ;
 wire \ces_7_1_io_ins_left[48] ;
 wire \ces_7_1_io_ins_left[49] ;
 wire \ces_7_1_io_ins_left[4] ;
 wire \ces_7_1_io_ins_left[50] ;
 wire \ces_7_1_io_ins_left[51] ;
 wire \ces_7_1_io_ins_left[52] ;
 wire \ces_7_1_io_ins_left[53] ;
 wire \ces_7_1_io_ins_left[54] ;
 wire \ces_7_1_io_ins_left[55] ;
 wire \ces_7_1_io_ins_left[56] ;
 wire \ces_7_1_io_ins_left[57] ;
 wire \ces_7_1_io_ins_left[58] ;
 wire \ces_7_1_io_ins_left[59] ;
 wire \ces_7_1_io_ins_left[5] ;
 wire \ces_7_1_io_ins_left[60] ;
 wire \ces_7_1_io_ins_left[61] ;
 wire \ces_7_1_io_ins_left[62] ;
 wire \ces_7_1_io_ins_left[63] ;
 wire \ces_7_1_io_ins_left[6] ;
 wire \ces_7_1_io_ins_left[7] ;
 wire \ces_7_1_io_ins_left[8] ;
 wire \ces_7_1_io_ins_left[9] ;
 wire ces_7_1_io_lsbOuts_0;
 wire ces_7_1_io_lsbOuts_1;
 wire ces_7_1_io_lsbOuts_2;
 wire ces_7_1_io_lsbOuts_3;
 wire ces_7_1_io_lsbOuts_4;
 wire ces_7_1_io_lsbOuts_5;
 wire ces_7_1_io_lsbOuts_6;
 wire ces_7_1_io_lsbOuts_7;
 wire \ces_7_1_io_outs_right[0] ;
 wire \ces_7_1_io_outs_right[10] ;
 wire \ces_7_1_io_outs_right[11] ;
 wire \ces_7_1_io_outs_right[12] ;
 wire \ces_7_1_io_outs_right[13] ;
 wire \ces_7_1_io_outs_right[14] ;
 wire \ces_7_1_io_outs_right[15] ;
 wire \ces_7_1_io_outs_right[16] ;
 wire \ces_7_1_io_outs_right[17] ;
 wire \ces_7_1_io_outs_right[18] ;
 wire \ces_7_1_io_outs_right[19] ;
 wire \ces_7_1_io_outs_right[1] ;
 wire \ces_7_1_io_outs_right[20] ;
 wire \ces_7_1_io_outs_right[21] ;
 wire \ces_7_1_io_outs_right[22] ;
 wire \ces_7_1_io_outs_right[23] ;
 wire \ces_7_1_io_outs_right[24] ;
 wire \ces_7_1_io_outs_right[25] ;
 wire \ces_7_1_io_outs_right[26] ;
 wire \ces_7_1_io_outs_right[27] ;
 wire \ces_7_1_io_outs_right[28] ;
 wire \ces_7_1_io_outs_right[29] ;
 wire \ces_7_1_io_outs_right[2] ;
 wire \ces_7_1_io_outs_right[30] ;
 wire \ces_7_1_io_outs_right[31] ;
 wire \ces_7_1_io_outs_right[32] ;
 wire \ces_7_1_io_outs_right[33] ;
 wire \ces_7_1_io_outs_right[34] ;
 wire \ces_7_1_io_outs_right[35] ;
 wire \ces_7_1_io_outs_right[36] ;
 wire \ces_7_1_io_outs_right[37] ;
 wire \ces_7_1_io_outs_right[38] ;
 wire \ces_7_1_io_outs_right[39] ;
 wire \ces_7_1_io_outs_right[3] ;
 wire \ces_7_1_io_outs_right[40] ;
 wire \ces_7_1_io_outs_right[41] ;
 wire \ces_7_1_io_outs_right[42] ;
 wire \ces_7_1_io_outs_right[43] ;
 wire \ces_7_1_io_outs_right[44] ;
 wire \ces_7_1_io_outs_right[45] ;
 wire \ces_7_1_io_outs_right[46] ;
 wire \ces_7_1_io_outs_right[47] ;
 wire \ces_7_1_io_outs_right[48] ;
 wire \ces_7_1_io_outs_right[49] ;
 wire \ces_7_1_io_outs_right[4] ;
 wire \ces_7_1_io_outs_right[50] ;
 wire \ces_7_1_io_outs_right[51] ;
 wire \ces_7_1_io_outs_right[52] ;
 wire \ces_7_1_io_outs_right[53] ;
 wire \ces_7_1_io_outs_right[54] ;
 wire \ces_7_1_io_outs_right[55] ;
 wire \ces_7_1_io_outs_right[56] ;
 wire \ces_7_1_io_outs_right[57] ;
 wire \ces_7_1_io_outs_right[58] ;
 wire \ces_7_1_io_outs_right[59] ;
 wire \ces_7_1_io_outs_right[5] ;
 wire \ces_7_1_io_outs_right[60] ;
 wire \ces_7_1_io_outs_right[61] ;
 wire \ces_7_1_io_outs_right[62] ;
 wire \ces_7_1_io_outs_right[63] ;
 wire \ces_7_1_io_outs_right[6] ;
 wire \ces_7_1_io_outs_right[7] ;
 wire \ces_7_1_io_outs_right[8] ;
 wire \ces_7_1_io_outs_right[9] ;
 wire \ces_7_2_io_ins_left[0] ;
 wire \ces_7_2_io_ins_left[10] ;
 wire \ces_7_2_io_ins_left[11] ;
 wire \ces_7_2_io_ins_left[12] ;
 wire \ces_7_2_io_ins_left[13] ;
 wire \ces_7_2_io_ins_left[14] ;
 wire \ces_7_2_io_ins_left[15] ;
 wire \ces_7_2_io_ins_left[16] ;
 wire \ces_7_2_io_ins_left[17] ;
 wire \ces_7_2_io_ins_left[18] ;
 wire \ces_7_2_io_ins_left[19] ;
 wire \ces_7_2_io_ins_left[1] ;
 wire \ces_7_2_io_ins_left[20] ;
 wire \ces_7_2_io_ins_left[21] ;
 wire \ces_7_2_io_ins_left[22] ;
 wire \ces_7_2_io_ins_left[23] ;
 wire \ces_7_2_io_ins_left[24] ;
 wire \ces_7_2_io_ins_left[25] ;
 wire \ces_7_2_io_ins_left[26] ;
 wire \ces_7_2_io_ins_left[27] ;
 wire \ces_7_2_io_ins_left[28] ;
 wire \ces_7_2_io_ins_left[29] ;
 wire \ces_7_2_io_ins_left[2] ;
 wire \ces_7_2_io_ins_left[30] ;
 wire \ces_7_2_io_ins_left[31] ;
 wire \ces_7_2_io_ins_left[32] ;
 wire \ces_7_2_io_ins_left[33] ;
 wire \ces_7_2_io_ins_left[34] ;
 wire \ces_7_2_io_ins_left[35] ;
 wire \ces_7_2_io_ins_left[36] ;
 wire \ces_7_2_io_ins_left[37] ;
 wire \ces_7_2_io_ins_left[38] ;
 wire \ces_7_2_io_ins_left[39] ;
 wire \ces_7_2_io_ins_left[3] ;
 wire \ces_7_2_io_ins_left[40] ;
 wire \ces_7_2_io_ins_left[41] ;
 wire \ces_7_2_io_ins_left[42] ;
 wire \ces_7_2_io_ins_left[43] ;
 wire \ces_7_2_io_ins_left[44] ;
 wire \ces_7_2_io_ins_left[45] ;
 wire \ces_7_2_io_ins_left[46] ;
 wire \ces_7_2_io_ins_left[47] ;
 wire \ces_7_2_io_ins_left[48] ;
 wire \ces_7_2_io_ins_left[49] ;
 wire \ces_7_2_io_ins_left[4] ;
 wire \ces_7_2_io_ins_left[50] ;
 wire \ces_7_2_io_ins_left[51] ;
 wire \ces_7_2_io_ins_left[52] ;
 wire \ces_7_2_io_ins_left[53] ;
 wire \ces_7_2_io_ins_left[54] ;
 wire \ces_7_2_io_ins_left[55] ;
 wire \ces_7_2_io_ins_left[56] ;
 wire \ces_7_2_io_ins_left[57] ;
 wire \ces_7_2_io_ins_left[58] ;
 wire \ces_7_2_io_ins_left[59] ;
 wire \ces_7_2_io_ins_left[5] ;
 wire \ces_7_2_io_ins_left[60] ;
 wire \ces_7_2_io_ins_left[61] ;
 wire \ces_7_2_io_ins_left[62] ;
 wire \ces_7_2_io_ins_left[63] ;
 wire \ces_7_2_io_ins_left[6] ;
 wire \ces_7_2_io_ins_left[7] ;
 wire \ces_7_2_io_ins_left[8] ;
 wire \ces_7_2_io_ins_left[9] ;
 wire ces_7_2_io_lsbOuts_0;
 wire ces_7_2_io_lsbOuts_1;
 wire ces_7_2_io_lsbOuts_2;
 wire ces_7_2_io_lsbOuts_3;
 wire ces_7_2_io_lsbOuts_4;
 wire ces_7_2_io_lsbOuts_5;
 wire ces_7_2_io_lsbOuts_6;
 wire ces_7_2_io_lsbOuts_7;
 wire \ces_7_2_io_outs_right[0] ;
 wire \ces_7_2_io_outs_right[10] ;
 wire \ces_7_2_io_outs_right[11] ;
 wire \ces_7_2_io_outs_right[12] ;
 wire \ces_7_2_io_outs_right[13] ;
 wire \ces_7_2_io_outs_right[14] ;
 wire \ces_7_2_io_outs_right[15] ;
 wire \ces_7_2_io_outs_right[16] ;
 wire \ces_7_2_io_outs_right[17] ;
 wire \ces_7_2_io_outs_right[18] ;
 wire \ces_7_2_io_outs_right[19] ;
 wire \ces_7_2_io_outs_right[1] ;
 wire \ces_7_2_io_outs_right[20] ;
 wire \ces_7_2_io_outs_right[21] ;
 wire \ces_7_2_io_outs_right[22] ;
 wire \ces_7_2_io_outs_right[23] ;
 wire \ces_7_2_io_outs_right[24] ;
 wire \ces_7_2_io_outs_right[25] ;
 wire \ces_7_2_io_outs_right[26] ;
 wire \ces_7_2_io_outs_right[27] ;
 wire \ces_7_2_io_outs_right[28] ;
 wire \ces_7_2_io_outs_right[29] ;
 wire \ces_7_2_io_outs_right[2] ;
 wire \ces_7_2_io_outs_right[30] ;
 wire \ces_7_2_io_outs_right[31] ;
 wire \ces_7_2_io_outs_right[32] ;
 wire \ces_7_2_io_outs_right[33] ;
 wire \ces_7_2_io_outs_right[34] ;
 wire \ces_7_2_io_outs_right[35] ;
 wire \ces_7_2_io_outs_right[36] ;
 wire \ces_7_2_io_outs_right[37] ;
 wire \ces_7_2_io_outs_right[38] ;
 wire \ces_7_2_io_outs_right[39] ;
 wire \ces_7_2_io_outs_right[3] ;
 wire \ces_7_2_io_outs_right[40] ;
 wire \ces_7_2_io_outs_right[41] ;
 wire \ces_7_2_io_outs_right[42] ;
 wire \ces_7_2_io_outs_right[43] ;
 wire \ces_7_2_io_outs_right[44] ;
 wire \ces_7_2_io_outs_right[45] ;
 wire \ces_7_2_io_outs_right[46] ;
 wire \ces_7_2_io_outs_right[47] ;
 wire \ces_7_2_io_outs_right[48] ;
 wire \ces_7_2_io_outs_right[49] ;
 wire \ces_7_2_io_outs_right[4] ;
 wire \ces_7_2_io_outs_right[50] ;
 wire \ces_7_2_io_outs_right[51] ;
 wire \ces_7_2_io_outs_right[52] ;
 wire \ces_7_2_io_outs_right[53] ;
 wire \ces_7_2_io_outs_right[54] ;
 wire \ces_7_2_io_outs_right[55] ;
 wire \ces_7_2_io_outs_right[56] ;
 wire \ces_7_2_io_outs_right[57] ;
 wire \ces_7_2_io_outs_right[58] ;
 wire \ces_7_2_io_outs_right[59] ;
 wire \ces_7_2_io_outs_right[5] ;
 wire \ces_7_2_io_outs_right[60] ;
 wire \ces_7_2_io_outs_right[61] ;
 wire \ces_7_2_io_outs_right[62] ;
 wire \ces_7_2_io_outs_right[63] ;
 wire \ces_7_2_io_outs_right[6] ;
 wire \ces_7_2_io_outs_right[7] ;
 wire \ces_7_2_io_outs_right[8] ;
 wire \ces_7_2_io_outs_right[9] ;
 wire \ces_7_3_io_ins_left[0] ;
 wire \ces_7_3_io_ins_left[10] ;
 wire \ces_7_3_io_ins_left[11] ;
 wire \ces_7_3_io_ins_left[12] ;
 wire \ces_7_3_io_ins_left[13] ;
 wire \ces_7_3_io_ins_left[14] ;
 wire \ces_7_3_io_ins_left[15] ;
 wire \ces_7_3_io_ins_left[16] ;
 wire \ces_7_3_io_ins_left[17] ;
 wire \ces_7_3_io_ins_left[18] ;
 wire \ces_7_3_io_ins_left[19] ;
 wire \ces_7_3_io_ins_left[1] ;
 wire \ces_7_3_io_ins_left[20] ;
 wire \ces_7_3_io_ins_left[21] ;
 wire \ces_7_3_io_ins_left[22] ;
 wire \ces_7_3_io_ins_left[23] ;
 wire \ces_7_3_io_ins_left[24] ;
 wire \ces_7_3_io_ins_left[25] ;
 wire \ces_7_3_io_ins_left[26] ;
 wire \ces_7_3_io_ins_left[27] ;
 wire \ces_7_3_io_ins_left[28] ;
 wire \ces_7_3_io_ins_left[29] ;
 wire \ces_7_3_io_ins_left[2] ;
 wire \ces_7_3_io_ins_left[30] ;
 wire \ces_7_3_io_ins_left[31] ;
 wire \ces_7_3_io_ins_left[32] ;
 wire \ces_7_3_io_ins_left[33] ;
 wire \ces_7_3_io_ins_left[34] ;
 wire \ces_7_3_io_ins_left[35] ;
 wire \ces_7_3_io_ins_left[36] ;
 wire \ces_7_3_io_ins_left[37] ;
 wire \ces_7_3_io_ins_left[38] ;
 wire \ces_7_3_io_ins_left[39] ;
 wire \ces_7_3_io_ins_left[3] ;
 wire \ces_7_3_io_ins_left[40] ;
 wire \ces_7_3_io_ins_left[41] ;
 wire \ces_7_3_io_ins_left[42] ;
 wire \ces_7_3_io_ins_left[43] ;
 wire \ces_7_3_io_ins_left[44] ;
 wire \ces_7_3_io_ins_left[45] ;
 wire \ces_7_3_io_ins_left[46] ;
 wire \ces_7_3_io_ins_left[47] ;
 wire \ces_7_3_io_ins_left[48] ;
 wire \ces_7_3_io_ins_left[49] ;
 wire \ces_7_3_io_ins_left[4] ;
 wire \ces_7_3_io_ins_left[50] ;
 wire \ces_7_3_io_ins_left[51] ;
 wire \ces_7_3_io_ins_left[52] ;
 wire \ces_7_3_io_ins_left[53] ;
 wire \ces_7_3_io_ins_left[54] ;
 wire \ces_7_3_io_ins_left[55] ;
 wire \ces_7_3_io_ins_left[56] ;
 wire \ces_7_3_io_ins_left[57] ;
 wire \ces_7_3_io_ins_left[58] ;
 wire \ces_7_3_io_ins_left[59] ;
 wire \ces_7_3_io_ins_left[5] ;
 wire \ces_7_3_io_ins_left[60] ;
 wire \ces_7_3_io_ins_left[61] ;
 wire \ces_7_3_io_ins_left[62] ;
 wire \ces_7_3_io_ins_left[63] ;
 wire \ces_7_3_io_ins_left[6] ;
 wire \ces_7_3_io_ins_left[7] ;
 wire \ces_7_3_io_ins_left[8] ;
 wire \ces_7_3_io_ins_left[9] ;
 wire ces_7_3_io_lsbOuts_0;
 wire ces_7_3_io_lsbOuts_1;
 wire ces_7_3_io_lsbOuts_2;
 wire ces_7_3_io_lsbOuts_3;
 wire ces_7_3_io_lsbOuts_4;
 wire ces_7_3_io_lsbOuts_5;
 wire ces_7_3_io_lsbOuts_6;
 wire ces_7_3_io_lsbOuts_7;
 wire \ces_7_3_io_outs_right[0] ;
 wire \ces_7_3_io_outs_right[10] ;
 wire \ces_7_3_io_outs_right[11] ;
 wire \ces_7_3_io_outs_right[12] ;
 wire \ces_7_3_io_outs_right[13] ;
 wire \ces_7_3_io_outs_right[14] ;
 wire \ces_7_3_io_outs_right[15] ;
 wire \ces_7_3_io_outs_right[16] ;
 wire \ces_7_3_io_outs_right[17] ;
 wire \ces_7_3_io_outs_right[18] ;
 wire \ces_7_3_io_outs_right[19] ;
 wire \ces_7_3_io_outs_right[1] ;
 wire \ces_7_3_io_outs_right[20] ;
 wire \ces_7_3_io_outs_right[21] ;
 wire \ces_7_3_io_outs_right[22] ;
 wire \ces_7_3_io_outs_right[23] ;
 wire \ces_7_3_io_outs_right[24] ;
 wire \ces_7_3_io_outs_right[25] ;
 wire \ces_7_3_io_outs_right[26] ;
 wire \ces_7_3_io_outs_right[27] ;
 wire \ces_7_3_io_outs_right[28] ;
 wire \ces_7_3_io_outs_right[29] ;
 wire \ces_7_3_io_outs_right[2] ;
 wire \ces_7_3_io_outs_right[30] ;
 wire \ces_7_3_io_outs_right[31] ;
 wire \ces_7_3_io_outs_right[32] ;
 wire \ces_7_3_io_outs_right[33] ;
 wire \ces_7_3_io_outs_right[34] ;
 wire \ces_7_3_io_outs_right[35] ;
 wire \ces_7_3_io_outs_right[36] ;
 wire \ces_7_3_io_outs_right[37] ;
 wire \ces_7_3_io_outs_right[38] ;
 wire \ces_7_3_io_outs_right[39] ;
 wire \ces_7_3_io_outs_right[3] ;
 wire \ces_7_3_io_outs_right[40] ;
 wire \ces_7_3_io_outs_right[41] ;
 wire \ces_7_3_io_outs_right[42] ;
 wire \ces_7_3_io_outs_right[43] ;
 wire \ces_7_3_io_outs_right[44] ;
 wire \ces_7_3_io_outs_right[45] ;
 wire \ces_7_3_io_outs_right[46] ;
 wire \ces_7_3_io_outs_right[47] ;
 wire \ces_7_3_io_outs_right[48] ;
 wire \ces_7_3_io_outs_right[49] ;
 wire \ces_7_3_io_outs_right[4] ;
 wire \ces_7_3_io_outs_right[50] ;
 wire \ces_7_3_io_outs_right[51] ;
 wire \ces_7_3_io_outs_right[52] ;
 wire \ces_7_3_io_outs_right[53] ;
 wire \ces_7_3_io_outs_right[54] ;
 wire \ces_7_3_io_outs_right[55] ;
 wire \ces_7_3_io_outs_right[56] ;
 wire \ces_7_3_io_outs_right[57] ;
 wire \ces_7_3_io_outs_right[58] ;
 wire \ces_7_3_io_outs_right[59] ;
 wire \ces_7_3_io_outs_right[5] ;
 wire \ces_7_3_io_outs_right[60] ;
 wire \ces_7_3_io_outs_right[61] ;
 wire \ces_7_3_io_outs_right[62] ;
 wire \ces_7_3_io_outs_right[63] ;
 wire \ces_7_3_io_outs_right[6] ;
 wire \ces_7_3_io_outs_right[7] ;
 wire \ces_7_3_io_outs_right[8] ;
 wire \ces_7_3_io_outs_right[9] ;
 wire \ces_7_4_io_ins_left[0] ;
 wire \ces_7_4_io_ins_left[10] ;
 wire \ces_7_4_io_ins_left[11] ;
 wire \ces_7_4_io_ins_left[12] ;
 wire \ces_7_4_io_ins_left[13] ;
 wire \ces_7_4_io_ins_left[14] ;
 wire \ces_7_4_io_ins_left[15] ;
 wire \ces_7_4_io_ins_left[16] ;
 wire \ces_7_4_io_ins_left[17] ;
 wire \ces_7_4_io_ins_left[18] ;
 wire \ces_7_4_io_ins_left[19] ;
 wire \ces_7_4_io_ins_left[1] ;
 wire \ces_7_4_io_ins_left[20] ;
 wire \ces_7_4_io_ins_left[21] ;
 wire \ces_7_4_io_ins_left[22] ;
 wire \ces_7_4_io_ins_left[23] ;
 wire \ces_7_4_io_ins_left[24] ;
 wire \ces_7_4_io_ins_left[25] ;
 wire \ces_7_4_io_ins_left[26] ;
 wire \ces_7_4_io_ins_left[27] ;
 wire \ces_7_4_io_ins_left[28] ;
 wire \ces_7_4_io_ins_left[29] ;
 wire \ces_7_4_io_ins_left[2] ;
 wire \ces_7_4_io_ins_left[30] ;
 wire \ces_7_4_io_ins_left[31] ;
 wire \ces_7_4_io_ins_left[32] ;
 wire \ces_7_4_io_ins_left[33] ;
 wire \ces_7_4_io_ins_left[34] ;
 wire \ces_7_4_io_ins_left[35] ;
 wire \ces_7_4_io_ins_left[36] ;
 wire \ces_7_4_io_ins_left[37] ;
 wire \ces_7_4_io_ins_left[38] ;
 wire \ces_7_4_io_ins_left[39] ;
 wire \ces_7_4_io_ins_left[3] ;
 wire \ces_7_4_io_ins_left[40] ;
 wire \ces_7_4_io_ins_left[41] ;
 wire \ces_7_4_io_ins_left[42] ;
 wire \ces_7_4_io_ins_left[43] ;
 wire \ces_7_4_io_ins_left[44] ;
 wire \ces_7_4_io_ins_left[45] ;
 wire \ces_7_4_io_ins_left[46] ;
 wire \ces_7_4_io_ins_left[47] ;
 wire \ces_7_4_io_ins_left[48] ;
 wire \ces_7_4_io_ins_left[49] ;
 wire \ces_7_4_io_ins_left[4] ;
 wire \ces_7_4_io_ins_left[50] ;
 wire \ces_7_4_io_ins_left[51] ;
 wire \ces_7_4_io_ins_left[52] ;
 wire \ces_7_4_io_ins_left[53] ;
 wire \ces_7_4_io_ins_left[54] ;
 wire \ces_7_4_io_ins_left[55] ;
 wire \ces_7_4_io_ins_left[56] ;
 wire \ces_7_4_io_ins_left[57] ;
 wire \ces_7_4_io_ins_left[58] ;
 wire \ces_7_4_io_ins_left[59] ;
 wire \ces_7_4_io_ins_left[5] ;
 wire \ces_7_4_io_ins_left[60] ;
 wire \ces_7_4_io_ins_left[61] ;
 wire \ces_7_4_io_ins_left[62] ;
 wire \ces_7_4_io_ins_left[63] ;
 wire \ces_7_4_io_ins_left[6] ;
 wire \ces_7_4_io_ins_left[7] ;
 wire \ces_7_4_io_ins_left[8] ;
 wire \ces_7_4_io_ins_left[9] ;
 wire ces_7_4_io_lsbOuts_0;
 wire ces_7_4_io_lsbOuts_1;
 wire ces_7_4_io_lsbOuts_2;
 wire ces_7_4_io_lsbOuts_3;
 wire ces_7_4_io_lsbOuts_4;
 wire ces_7_4_io_lsbOuts_5;
 wire ces_7_4_io_lsbOuts_6;
 wire ces_7_4_io_lsbOuts_7;
 wire \ces_7_4_io_outs_right[0] ;
 wire \ces_7_4_io_outs_right[10] ;
 wire \ces_7_4_io_outs_right[11] ;
 wire \ces_7_4_io_outs_right[12] ;
 wire \ces_7_4_io_outs_right[13] ;
 wire \ces_7_4_io_outs_right[14] ;
 wire \ces_7_4_io_outs_right[15] ;
 wire \ces_7_4_io_outs_right[16] ;
 wire \ces_7_4_io_outs_right[17] ;
 wire \ces_7_4_io_outs_right[18] ;
 wire \ces_7_4_io_outs_right[19] ;
 wire \ces_7_4_io_outs_right[1] ;
 wire \ces_7_4_io_outs_right[20] ;
 wire \ces_7_4_io_outs_right[21] ;
 wire \ces_7_4_io_outs_right[22] ;
 wire \ces_7_4_io_outs_right[23] ;
 wire \ces_7_4_io_outs_right[24] ;
 wire \ces_7_4_io_outs_right[25] ;
 wire \ces_7_4_io_outs_right[26] ;
 wire \ces_7_4_io_outs_right[27] ;
 wire \ces_7_4_io_outs_right[28] ;
 wire \ces_7_4_io_outs_right[29] ;
 wire \ces_7_4_io_outs_right[2] ;
 wire \ces_7_4_io_outs_right[30] ;
 wire \ces_7_4_io_outs_right[31] ;
 wire \ces_7_4_io_outs_right[32] ;
 wire \ces_7_4_io_outs_right[33] ;
 wire \ces_7_4_io_outs_right[34] ;
 wire \ces_7_4_io_outs_right[35] ;
 wire \ces_7_4_io_outs_right[36] ;
 wire \ces_7_4_io_outs_right[37] ;
 wire \ces_7_4_io_outs_right[38] ;
 wire \ces_7_4_io_outs_right[39] ;
 wire \ces_7_4_io_outs_right[3] ;
 wire \ces_7_4_io_outs_right[40] ;
 wire \ces_7_4_io_outs_right[41] ;
 wire \ces_7_4_io_outs_right[42] ;
 wire \ces_7_4_io_outs_right[43] ;
 wire \ces_7_4_io_outs_right[44] ;
 wire \ces_7_4_io_outs_right[45] ;
 wire \ces_7_4_io_outs_right[46] ;
 wire \ces_7_4_io_outs_right[47] ;
 wire \ces_7_4_io_outs_right[48] ;
 wire \ces_7_4_io_outs_right[49] ;
 wire \ces_7_4_io_outs_right[4] ;
 wire \ces_7_4_io_outs_right[50] ;
 wire \ces_7_4_io_outs_right[51] ;
 wire \ces_7_4_io_outs_right[52] ;
 wire \ces_7_4_io_outs_right[53] ;
 wire \ces_7_4_io_outs_right[54] ;
 wire \ces_7_4_io_outs_right[55] ;
 wire \ces_7_4_io_outs_right[56] ;
 wire \ces_7_4_io_outs_right[57] ;
 wire \ces_7_4_io_outs_right[58] ;
 wire \ces_7_4_io_outs_right[59] ;
 wire \ces_7_4_io_outs_right[5] ;
 wire \ces_7_4_io_outs_right[60] ;
 wire \ces_7_4_io_outs_right[61] ;
 wire \ces_7_4_io_outs_right[62] ;
 wire \ces_7_4_io_outs_right[63] ;
 wire \ces_7_4_io_outs_right[6] ;
 wire \ces_7_4_io_outs_right[7] ;
 wire \ces_7_4_io_outs_right[8] ;
 wire \ces_7_4_io_outs_right[9] ;
 wire \ces_7_5_io_ins_left[0] ;
 wire \ces_7_5_io_ins_left[10] ;
 wire \ces_7_5_io_ins_left[11] ;
 wire \ces_7_5_io_ins_left[12] ;
 wire \ces_7_5_io_ins_left[13] ;
 wire \ces_7_5_io_ins_left[14] ;
 wire \ces_7_5_io_ins_left[15] ;
 wire \ces_7_5_io_ins_left[16] ;
 wire \ces_7_5_io_ins_left[17] ;
 wire \ces_7_5_io_ins_left[18] ;
 wire \ces_7_5_io_ins_left[19] ;
 wire \ces_7_5_io_ins_left[1] ;
 wire \ces_7_5_io_ins_left[20] ;
 wire \ces_7_5_io_ins_left[21] ;
 wire \ces_7_5_io_ins_left[22] ;
 wire \ces_7_5_io_ins_left[23] ;
 wire \ces_7_5_io_ins_left[24] ;
 wire \ces_7_5_io_ins_left[25] ;
 wire \ces_7_5_io_ins_left[26] ;
 wire \ces_7_5_io_ins_left[27] ;
 wire \ces_7_5_io_ins_left[28] ;
 wire \ces_7_5_io_ins_left[29] ;
 wire \ces_7_5_io_ins_left[2] ;
 wire \ces_7_5_io_ins_left[30] ;
 wire \ces_7_5_io_ins_left[31] ;
 wire \ces_7_5_io_ins_left[32] ;
 wire \ces_7_5_io_ins_left[33] ;
 wire \ces_7_5_io_ins_left[34] ;
 wire \ces_7_5_io_ins_left[35] ;
 wire \ces_7_5_io_ins_left[36] ;
 wire \ces_7_5_io_ins_left[37] ;
 wire \ces_7_5_io_ins_left[38] ;
 wire \ces_7_5_io_ins_left[39] ;
 wire \ces_7_5_io_ins_left[3] ;
 wire \ces_7_5_io_ins_left[40] ;
 wire \ces_7_5_io_ins_left[41] ;
 wire \ces_7_5_io_ins_left[42] ;
 wire \ces_7_5_io_ins_left[43] ;
 wire \ces_7_5_io_ins_left[44] ;
 wire \ces_7_5_io_ins_left[45] ;
 wire \ces_7_5_io_ins_left[46] ;
 wire \ces_7_5_io_ins_left[47] ;
 wire \ces_7_5_io_ins_left[48] ;
 wire \ces_7_5_io_ins_left[49] ;
 wire \ces_7_5_io_ins_left[4] ;
 wire \ces_7_5_io_ins_left[50] ;
 wire \ces_7_5_io_ins_left[51] ;
 wire \ces_7_5_io_ins_left[52] ;
 wire \ces_7_5_io_ins_left[53] ;
 wire \ces_7_5_io_ins_left[54] ;
 wire \ces_7_5_io_ins_left[55] ;
 wire \ces_7_5_io_ins_left[56] ;
 wire \ces_7_5_io_ins_left[57] ;
 wire \ces_7_5_io_ins_left[58] ;
 wire \ces_7_5_io_ins_left[59] ;
 wire \ces_7_5_io_ins_left[5] ;
 wire \ces_7_5_io_ins_left[60] ;
 wire \ces_7_5_io_ins_left[61] ;
 wire \ces_7_5_io_ins_left[62] ;
 wire \ces_7_5_io_ins_left[63] ;
 wire \ces_7_5_io_ins_left[6] ;
 wire \ces_7_5_io_ins_left[7] ;
 wire \ces_7_5_io_ins_left[8] ;
 wire \ces_7_5_io_ins_left[9] ;
 wire ces_7_5_io_lsbOuts_0;
 wire ces_7_5_io_lsbOuts_1;
 wire ces_7_5_io_lsbOuts_2;
 wire ces_7_5_io_lsbOuts_3;
 wire ces_7_5_io_lsbOuts_4;
 wire ces_7_5_io_lsbOuts_5;
 wire ces_7_5_io_lsbOuts_6;
 wire ces_7_5_io_lsbOuts_7;
 wire \ces_7_5_io_outs_right[0] ;
 wire \ces_7_5_io_outs_right[10] ;
 wire \ces_7_5_io_outs_right[11] ;
 wire \ces_7_5_io_outs_right[12] ;
 wire \ces_7_5_io_outs_right[13] ;
 wire \ces_7_5_io_outs_right[14] ;
 wire \ces_7_5_io_outs_right[15] ;
 wire \ces_7_5_io_outs_right[16] ;
 wire \ces_7_5_io_outs_right[17] ;
 wire \ces_7_5_io_outs_right[18] ;
 wire \ces_7_5_io_outs_right[19] ;
 wire \ces_7_5_io_outs_right[1] ;
 wire \ces_7_5_io_outs_right[20] ;
 wire \ces_7_5_io_outs_right[21] ;
 wire \ces_7_5_io_outs_right[22] ;
 wire \ces_7_5_io_outs_right[23] ;
 wire \ces_7_5_io_outs_right[24] ;
 wire \ces_7_5_io_outs_right[25] ;
 wire \ces_7_5_io_outs_right[26] ;
 wire \ces_7_5_io_outs_right[27] ;
 wire \ces_7_5_io_outs_right[28] ;
 wire \ces_7_5_io_outs_right[29] ;
 wire \ces_7_5_io_outs_right[2] ;
 wire \ces_7_5_io_outs_right[30] ;
 wire \ces_7_5_io_outs_right[31] ;
 wire \ces_7_5_io_outs_right[32] ;
 wire \ces_7_5_io_outs_right[33] ;
 wire \ces_7_5_io_outs_right[34] ;
 wire \ces_7_5_io_outs_right[35] ;
 wire \ces_7_5_io_outs_right[36] ;
 wire \ces_7_5_io_outs_right[37] ;
 wire \ces_7_5_io_outs_right[38] ;
 wire \ces_7_5_io_outs_right[39] ;
 wire \ces_7_5_io_outs_right[3] ;
 wire \ces_7_5_io_outs_right[40] ;
 wire \ces_7_5_io_outs_right[41] ;
 wire \ces_7_5_io_outs_right[42] ;
 wire \ces_7_5_io_outs_right[43] ;
 wire \ces_7_5_io_outs_right[44] ;
 wire \ces_7_5_io_outs_right[45] ;
 wire \ces_7_5_io_outs_right[46] ;
 wire \ces_7_5_io_outs_right[47] ;
 wire \ces_7_5_io_outs_right[48] ;
 wire \ces_7_5_io_outs_right[49] ;
 wire \ces_7_5_io_outs_right[4] ;
 wire \ces_7_5_io_outs_right[50] ;
 wire \ces_7_5_io_outs_right[51] ;
 wire \ces_7_5_io_outs_right[52] ;
 wire \ces_7_5_io_outs_right[53] ;
 wire \ces_7_5_io_outs_right[54] ;
 wire \ces_7_5_io_outs_right[55] ;
 wire \ces_7_5_io_outs_right[56] ;
 wire \ces_7_5_io_outs_right[57] ;
 wire \ces_7_5_io_outs_right[58] ;
 wire \ces_7_5_io_outs_right[59] ;
 wire \ces_7_5_io_outs_right[5] ;
 wire \ces_7_5_io_outs_right[60] ;
 wire \ces_7_5_io_outs_right[61] ;
 wire \ces_7_5_io_outs_right[62] ;
 wire \ces_7_5_io_outs_right[63] ;
 wire \ces_7_5_io_outs_right[6] ;
 wire \ces_7_5_io_outs_right[7] ;
 wire \ces_7_5_io_outs_right[8] ;
 wire \ces_7_5_io_outs_right[9] ;
 wire \ces_7_6_io_ins_left[0] ;
 wire \ces_7_6_io_ins_left[10] ;
 wire \ces_7_6_io_ins_left[11] ;
 wire \ces_7_6_io_ins_left[12] ;
 wire \ces_7_6_io_ins_left[13] ;
 wire \ces_7_6_io_ins_left[14] ;
 wire \ces_7_6_io_ins_left[15] ;
 wire \ces_7_6_io_ins_left[16] ;
 wire \ces_7_6_io_ins_left[17] ;
 wire \ces_7_6_io_ins_left[18] ;
 wire \ces_7_6_io_ins_left[19] ;
 wire \ces_7_6_io_ins_left[1] ;
 wire \ces_7_6_io_ins_left[20] ;
 wire \ces_7_6_io_ins_left[21] ;
 wire \ces_7_6_io_ins_left[22] ;
 wire \ces_7_6_io_ins_left[23] ;
 wire \ces_7_6_io_ins_left[24] ;
 wire \ces_7_6_io_ins_left[25] ;
 wire \ces_7_6_io_ins_left[26] ;
 wire \ces_7_6_io_ins_left[27] ;
 wire \ces_7_6_io_ins_left[28] ;
 wire \ces_7_6_io_ins_left[29] ;
 wire \ces_7_6_io_ins_left[2] ;
 wire \ces_7_6_io_ins_left[30] ;
 wire \ces_7_6_io_ins_left[31] ;
 wire \ces_7_6_io_ins_left[32] ;
 wire \ces_7_6_io_ins_left[33] ;
 wire \ces_7_6_io_ins_left[34] ;
 wire \ces_7_6_io_ins_left[35] ;
 wire \ces_7_6_io_ins_left[36] ;
 wire \ces_7_6_io_ins_left[37] ;
 wire \ces_7_6_io_ins_left[38] ;
 wire \ces_7_6_io_ins_left[39] ;
 wire \ces_7_6_io_ins_left[3] ;
 wire \ces_7_6_io_ins_left[40] ;
 wire \ces_7_6_io_ins_left[41] ;
 wire \ces_7_6_io_ins_left[42] ;
 wire \ces_7_6_io_ins_left[43] ;
 wire \ces_7_6_io_ins_left[44] ;
 wire \ces_7_6_io_ins_left[45] ;
 wire \ces_7_6_io_ins_left[46] ;
 wire \ces_7_6_io_ins_left[47] ;
 wire \ces_7_6_io_ins_left[48] ;
 wire \ces_7_6_io_ins_left[49] ;
 wire \ces_7_6_io_ins_left[4] ;
 wire \ces_7_6_io_ins_left[50] ;
 wire \ces_7_6_io_ins_left[51] ;
 wire \ces_7_6_io_ins_left[52] ;
 wire \ces_7_6_io_ins_left[53] ;
 wire \ces_7_6_io_ins_left[54] ;
 wire \ces_7_6_io_ins_left[55] ;
 wire \ces_7_6_io_ins_left[56] ;
 wire \ces_7_6_io_ins_left[57] ;
 wire \ces_7_6_io_ins_left[58] ;
 wire \ces_7_6_io_ins_left[59] ;
 wire \ces_7_6_io_ins_left[5] ;
 wire \ces_7_6_io_ins_left[60] ;
 wire \ces_7_6_io_ins_left[61] ;
 wire \ces_7_6_io_ins_left[62] ;
 wire \ces_7_6_io_ins_left[63] ;
 wire \ces_7_6_io_ins_left[6] ;
 wire \ces_7_6_io_ins_left[7] ;
 wire \ces_7_6_io_ins_left[8] ;
 wire \ces_7_6_io_ins_left[9] ;
 wire ces_7_6_io_lsbOuts_0;
 wire ces_7_6_io_lsbOuts_1;
 wire ces_7_6_io_lsbOuts_2;
 wire ces_7_6_io_lsbOuts_3;
 wire ces_7_6_io_lsbOuts_4;
 wire ces_7_6_io_lsbOuts_5;
 wire ces_7_6_io_lsbOuts_6;
 wire ces_7_6_io_lsbOuts_7;
 wire \ces_7_6_io_outs_right[0] ;
 wire \ces_7_6_io_outs_right[10] ;
 wire \ces_7_6_io_outs_right[11] ;
 wire \ces_7_6_io_outs_right[12] ;
 wire \ces_7_6_io_outs_right[13] ;
 wire \ces_7_6_io_outs_right[14] ;
 wire \ces_7_6_io_outs_right[15] ;
 wire \ces_7_6_io_outs_right[16] ;
 wire \ces_7_6_io_outs_right[17] ;
 wire \ces_7_6_io_outs_right[18] ;
 wire \ces_7_6_io_outs_right[19] ;
 wire \ces_7_6_io_outs_right[1] ;
 wire \ces_7_6_io_outs_right[20] ;
 wire \ces_7_6_io_outs_right[21] ;
 wire \ces_7_6_io_outs_right[22] ;
 wire \ces_7_6_io_outs_right[23] ;
 wire \ces_7_6_io_outs_right[24] ;
 wire \ces_7_6_io_outs_right[25] ;
 wire \ces_7_6_io_outs_right[26] ;
 wire \ces_7_6_io_outs_right[27] ;
 wire \ces_7_6_io_outs_right[28] ;
 wire \ces_7_6_io_outs_right[29] ;
 wire \ces_7_6_io_outs_right[2] ;
 wire \ces_7_6_io_outs_right[30] ;
 wire \ces_7_6_io_outs_right[31] ;
 wire \ces_7_6_io_outs_right[32] ;
 wire \ces_7_6_io_outs_right[33] ;
 wire \ces_7_6_io_outs_right[34] ;
 wire \ces_7_6_io_outs_right[35] ;
 wire \ces_7_6_io_outs_right[36] ;
 wire \ces_7_6_io_outs_right[37] ;
 wire \ces_7_6_io_outs_right[38] ;
 wire \ces_7_6_io_outs_right[39] ;
 wire \ces_7_6_io_outs_right[3] ;
 wire \ces_7_6_io_outs_right[40] ;
 wire \ces_7_6_io_outs_right[41] ;
 wire \ces_7_6_io_outs_right[42] ;
 wire \ces_7_6_io_outs_right[43] ;
 wire \ces_7_6_io_outs_right[44] ;
 wire \ces_7_6_io_outs_right[45] ;
 wire \ces_7_6_io_outs_right[46] ;
 wire \ces_7_6_io_outs_right[47] ;
 wire \ces_7_6_io_outs_right[48] ;
 wire \ces_7_6_io_outs_right[49] ;
 wire \ces_7_6_io_outs_right[4] ;
 wire \ces_7_6_io_outs_right[50] ;
 wire \ces_7_6_io_outs_right[51] ;
 wire \ces_7_6_io_outs_right[52] ;
 wire \ces_7_6_io_outs_right[53] ;
 wire \ces_7_6_io_outs_right[54] ;
 wire \ces_7_6_io_outs_right[55] ;
 wire \ces_7_6_io_outs_right[56] ;
 wire \ces_7_6_io_outs_right[57] ;
 wire \ces_7_6_io_outs_right[58] ;
 wire \ces_7_6_io_outs_right[59] ;
 wire \ces_7_6_io_outs_right[5] ;
 wire \ces_7_6_io_outs_right[60] ;
 wire \ces_7_6_io_outs_right[61] ;
 wire \ces_7_6_io_outs_right[62] ;
 wire \ces_7_6_io_outs_right[63] ;
 wire \ces_7_6_io_outs_right[6] ;
 wire \ces_7_6_io_outs_right[7] ;
 wire \ces_7_6_io_outs_right[8] ;
 wire \ces_7_6_io_outs_right[9] ;
 wire ces_7_7_io_lsbOuts_0;
 wire ces_7_7_io_lsbOuts_1;
 wire ces_7_7_io_lsbOuts_2;
 wire ces_7_7_io_lsbOuts_3;
 wire ces_7_7_io_lsbOuts_4;
 wire ces_7_7_io_lsbOuts_5;
 wire ces_7_7_io_lsbOuts_6;
 wire ces_7_7_io_lsbOuts_7;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire clknet_0_clock;
 wire clknet_1_0_0_clock;
 wire clknet_1_1_0_clock;
 wire clknet_2_0_0_clock;
 wire clknet_2_1_0_clock;
 wire clknet_2_2_0_clock;
 wire clknet_2_3_0_clock;
 wire clknet_3_0_0_clock;
 wire clknet_3_1_0_clock;
 wire clknet_3_2_0_clock;
 wire clknet_3_3_0_clock;
 wire clknet_3_4_0_clock;
 wire clknet_3_5_0_clock;
 wire clknet_3_6_0_clock;
 wire clknet_3_7_0_clock;
 wire clknet_0_clock_regs;
 wire clknet_3_0_0_clock_regs;
 wire clknet_3_1_0_clock_regs;
 wire clknet_3_2_0_clock_regs;
 wire clknet_3_3_0_clock_regs;
 wire clknet_3_4_0_clock_regs;
 wire clknet_3_5_0_clock_regs;
 wire clknet_3_6_0_clock_regs;
 wire clknet_3_7_0_clock_regs;
 wire delaynet_0_clock;
 wire delaynet_1_clock;
 wire delaynet_2_clock;
 wire delaynet_3_clock;
 wire delaynet_4_clock;
 wire delaynet_5_clock;
 wire net4217;
 wire net4218;

 INVx4_ASAP7_75t_R _065_ (.A(_000_),
    .Y(net2050));
 INVx4_ASAP7_75t_R _066_ (.A(_001_),
    .Y(net2049));
 INVx4_ASAP7_75t_R _067_ (.A(_002_),
    .Y(net2061));
 INVx3_ASAP7_75t_R _068_ (.A(_003_),
    .Y(net2072));
 INVx3_ASAP7_75t_R _069_ (.A(_004_),
    .Y(net2083));
 INVx4_ASAP7_75t_R _070_ (.A(_005_),
    .Y(net2094));
 INVx4_ASAP7_75t_R _071_ (.A(_006_),
    .Y(net2105));
 INVx4_ASAP7_75t_R _072_ (.A(_007_),
    .Y(net2110));
 INVx3_ASAP7_75t_R _073_ (.A(_008_),
    .Y(net2111));
 INVx3_ASAP7_75t_R _074_ (.A(_009_),
    .Y(net2112));
 INVx3_ASAP7_75t_R _075_ (.A(_010_),
    .Y(net2051));
 INVx3_ASAP7_75t_R _076_ (.A(_011_),
    .Y(net2052));
 INVx3_ASAP7_75t_R _077_ (.A(_012_),
    .Y(net2053));
 INVx3_ASAP7_75t_R _078_ (.A(_013_),
    .Y(net2054));
 INVx3_ASAP7_75t_R _079_ (.A(_014_),
    .Y(net2055));
 INVx3_ASAP7_75t_R _080_ (.A(_015_),
    .Y(net2056));
 INVx3_ASAP7_75t_R _081_ (.A(_016_),
    .Y(net2057));
 INVx3_ASAP7_75t_R _082_ (.A(_017_),
    .Y(net2058));
 INVx3_ASAP7_75t_R _083_ (.A(_018_),
    .Y(net2059));
 INVx3_ASAP7_75t_R _084_ (.A(_019_),
    .Y(net2060));
 INVx3_ASAP7_75t_R _085_ (.A(_020_),
    .Y(net2062));
 INVx3_ASAP7_75t_R _086_ (.A(_021_),
    .Y(net2063));
 INVx3_ASAP7_75t_R _087_ (.A(_022_),
    .Y(net2064));
 INVx3_ASAP7_75t_R _088_ (.A(_023_),
    .Y(net2065));
 INVx3_ASAP7_75t_R _089_ (.A(_024_),
    .Y(net2066));
 INVx3_ASAP7_75t_R _090_ (.A(_025_),
    .Y(net2067));
 INVx3_ASAP7_75t_R _091_ (.A(_026_),
    .Y(net2068));
 INVx3_ASAP7_75t_R _092_ (.A(_027_),
    .Y(net2069));
 INVx3_ASAP7_75t_R _093_ (.A(_028_),
    .Y(net2070));
 INVx3_ASAP7_75t_R _094_ (.A(_029_),
    .Y(net2071));
 INVx3_ASAP7_75t_R _095_ (.A(_030_),
    .Y(net2073));
 INVx3_ASAP7_75t_R _096_ (.A(_031_),
    .Y(net2074));
 INVx3_ASAP7_75t_R _097_ (.A(_032_),
    .Y(net2075));
 INVx3_ASAP7_75t_R _098_ (.A(_033_),
    .Y(net2076));
 INVx3_ASAP7_75t_R _099_ (.A(_034_),
    .Y(net2077));
 INVx3_ASAP7_75t_R _100_ (.A(_035_),
    .Y(net2078));
 INVx3_ASAP7_75t_R _101_ (.A(_036_),
    .Y(net2079));
 INVx3_ASAP7_75t_R _102_ (.A(_037_),
    .Y(net2080));
 INVx3_ASAP7_75t_R _103_ (.A(_038_),
    .Y(net2081));
 INVx3_ASAP7_75t_R _104_ (.A(_039_),
    .Y(net2082));
 INVx3_ASAP7_75t_R _105_ (.A(_040_),
    .Y(net2084));
 INVx3_ASAP7_75t_R _106_ (.A(_041_),
    .Y(net2085));
 INVx3_ASAP7_75t_R _107_ (.A(_042_),
    .Y(net2086));
 INVx3_ASAP7_75t_R _108_ (.A(_043_),
    .Y(net2087));
 INVx3_ASAP7_75t_R _109_ (.A(_044_),
    .Y(net2088));
 INVx3_ASAP7_75t_R _110_ (.A(_045_),
    .Y(net2089));
 INVx3_ASAP7_75t_R _111_ (.A(_046_),
    .Y(net2090));
 INVx3_ASAP7_75t_R _112_ (.A(_047_),
    .Y(net2091));
 INVx3_ASAP7_75t_R _113_ (.A(_048_),
    .Y(net2092));
 INVx3_ASAP7_75t_R _114_ (.A(_049_),
    .Y(net2093));
 INVx3_ASAP7_75t_R _115_ (.A(_050_),
    .Y(net2095));
 INVx3_ASAP7_75t_R _116_ (.A(_051_),
    .Y(net2096));
 INVx3_ASAP7_75t_R _117_ (.A(_052_),
    .Y(net2097));
 INVx3_ASAP7_75t_R _118_ (.A(_053_),
    .Y(net2098));
 INVx3_ASAP7_75t_R _119_ (.A(_054_),
    .Y(net2099));
 INVx3_ASAP7_75t_R _120_ (.A(_055_),
    .Y(net2100));
 INVx4_ASAP7_75t_R _121_ (.A(_056_),
    .Y(net2101));
 INVx4_ASAP7_75t_R _122_ (.A(_057_),
    .Y(net2102));
 INVx4_ASAP7_75t_R _123_ (.A(_058_),
    .Y(net2103));
 INVx4_ASAP7_75t_R _124_ (.A(_059_),
    .Y(net2104));
 INVx4_ASAP7_75t_R _125_ (.A(_060_),
    .Y(net2106));
 INVx4_ASAP7_75t_R _126_ (.A(_061_),
    .Y(net2107));
 INVx4_ASAP7_75t_R _127_ (.A(_062_),
    .Y(net2108));
 INVx4_ASAP7_75t_R _128_ (.A(_063_),
    .Y(net2109));
 BUFx24_ASAP7_75t_R clkbuf_regs_0_clock (.A(net4217),
    .Y(delaynet_0_clock));
 Element ces_0_0 (.clock(clknet_3_0_0_clock),
    .io_lsbIns_1(net4161),
    .io_lsbIns_2(net4162),
    .io_lsbIns_3(net4163),
    .io_lsbIns_4(net4164),
    .io_lsbIns_5(net4165),
    .io_lsbIns_6(net4166),
    .io_lsbIns_7(net4167),
    .io_lsbOuts_0(ces_0_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_0_io_lsbOuts_7),
    .io_ins_down({\ces_0_0_io_ins_down[63] ,
    \ces_0_0_io_ins_down[62] ,
    \ces_0_0_io_ins_down[61] ,
    \ces_0_0_io_ins_down[60] ,
    \ces_0_0_io_ins_down[59] ,
    \ces_0_0_io_ins_down[58] ,
    \ces_0_0_io_ins_down[57] ,
    \ces_0_0_io_ins_down[56] ,
    \ces_0_0_io_ins_down[55] ,
    \ces_0_0_io_ins_down[54] ,
    \ces_0_0_io_ins_down[53] ,
    \ces_0_0_io_ins_down[52] ,
    \ces_0_0_io_ins_down[51] ,
    \ces_0_0_io_ins_down[50] ,
    \ces_0_0_io_ins_down[49] ,
    \ces_0_0_io_ins_down[48] ,
    \ces_0_0_io_ins_down[47] ,
    \ces_0_0_io_ins_down[46] ,
    \ces_0_0_io_ins_down[45] ,
    \ces_0_0_io_ins_down[44] ,
    \ces_0_0_io_ins_down[43] ,
    \ces_0_0_io_ins_down[42] ,
    \ces_0_0_io_ins_down[41] ,
    \ces_0_0_io_ins_down[40] ,
    \ces_0_0_io_ins_down[39] ,
    \ces_0_0_io_ins_down[38] ,
    \ces_0_0_io_ins_down[37] ,
    \ces_0_0_io_ins_down[36] ,
    \ces_0_0_io_ins_down[35] ,
    \ces_0_0_io_ins_down[34] ,
    \ces_0_0_io_ins_down[33] ,
    \ces_0_0_io_ins_down[32] ,
    \ces_0_0_io_ins_down[31] ,
    \ces_0_0_io_ins_down[30] ,
    \ces_0_0_io_ins_down[29] ,
    \ces_0_0_io_ins_down[28] ,
    \ces_0_0_io_ins_down[27] ,
    \ces_0_0_io_ins_down[26] ,
    \ces_0_0_io_ins_down[25] ,
    \ces_0_0_io_ins_down[24] ,
    \ces_0_0_io_ins_down[23] ,
    \ces_0_0_io_ins_down[22] ,
    \ces_0_0_io_ins_down[21] ,
    \ces_0_0_io_ins_down[20] ,
    \ces_0_0_io_ins_down[19] ,
    \ces_0_0_io_ins_down[18] ,
    \ces_0_0_io_ins_down[17] ,
    \ces_0_0_io_ins_down[16] ,
    \ces_0_0_io_ins_down[15] ,
    \ces_0_0_io_ins_down[14] ,
    \ces_0_0_io_ins_down[13] ,
    \ces_0_0_io_ins_down[12] ,
    \ces_0_0_io_ins_down[11] ,
    \ces_0_0_io_ins_down[10] ,
    \ces_0_0_io_ins_down[9] ,
    \ces_0_0_io_ins_down[8] ,
    \ces_0_0_io_ins_down[7] ,
    \ces_0_0_io_ins_down[6] ,
    \ces_0_0_io_ins_down[5] ,
    \ces_0_0_io_ins_down[4] ,
    \ces_0_0_io_ins_down[3] ,
    \ces_0_0_io_ins_down[2] ,
    \ces_0_0_io_ins_down[1] ,
    \ces_0_0_io_ins_down[0] }),
    .io_ins_left({\ces_0_0_io_ins_left[63] ,
    \ces_0_0_io_ins_left[62] ,
    \ces_0_0_io_ins_left[61] ,
    \ces_0_0_io_ins_left[60] ,
    \ces_0_0_io_ins_left[59] ,
    \ces_0_0_io_ins_left[58] ,
    \ces_0_0_io_ins_left[57] ,
    \ces_0_0_io_ins_left[56] ,
    \ces_0_0_io_ins_left[55] ,
    \ces_0_0_io_ins_left[54] ,
    \ces_0_0_io_ins_left[53] ,
    \ces_0_0_io_ins_left[52] ,
    \ces_0_0_io_ins_left[51] ,
    \ces_0_0_io_ins_left[50] ,
    \ces_0_0_io_ins_left[49] ,
    \ces_0_0_io_ins_left[48] ,
    \ces_0_0_io_ins_left[47] ,
    \ces_0_0_io_ins_left[46] ,
    \ces_0_0_io_ins_left[45] ,
    \ces_0_0_io_ins_left[44] ,
    \ces_0_0_io_ins_left[43] ,
    \ces_0_0_io_ins_left[42] ,
    \ces_0_0_io_ins_left[41] ,
    \ces_0_0_io_ins_left[40] ,
    \ces_0_0_io_ins_left[39] ,
    \ces_0_0_io_ins_left[38] ,
    \ces_0_0_io_ins_left[37] ,
    \ces_0_0_io_ins_left[36] ,
    \ces_0_0_io_ins_left[35] ,
    \ces_0_0_io_ins_left[34] ,
    \ces_0_0_io_ins_left[33] ,
    \ces_0_0_io_ins_left[32] ,
    \ces_0_0_io_ins_left[31] ,
    \ces_0_0_io_ins_left[30] ,
    \ces_0_0_io_ins_left[29] ,
    \ces_0_0_io_ins_left[28] ,
    \ces_0_0_io_ins_left[27] ,
    \ces_0_0_io_ins_left[26] ,
    \ces_0_0_io_ins_left[25] ,
    \ces_0_0_io_ins_left[24] ,
    \ces_0_0_io_ins_left[23] ,
    \ces_0_0_io_ins_left[22] ,
    \ces_0_0_io_ins_left[21] ,
    \ces_0_0_io_ins_left[20] ,
    \ces_0_0_io_ins_left[19] ,
    \ces_0_0_io_ins_left[18] ,
    \ces_0_0_io_ins_left[17] ,
    \ces_0_0_io_ins_left[16] ,
    \ces_0_0_io_ins_left[15] ,
    \ces_0_0_io_ins_left[14] ,
    \ces_0_0_io_ins_left[13] ,
    \ces_0_0_io_ins_left[12] ,
    \ces_0_0_io_ins_left[11] ,
    \ces_0_0_io_ins_left[10] ,
    \ces_0_0_io_ins_left[9] ,
    \ces_0_0_io_ins_left[8] ,
    \ces_0_0_io_ins_left[7] ,
    \ces_0_0_io_ins_left[6] ,
    \ces_0_0_io_ins_left[5] ,
    \ces_0_0_io_ins_left[4] ,
    \ces_0_0_io_ins_left[3] ,
    \ces_0_0_io_ins_left[2] ,
    \ces_0_0_io_ins_left[1] ,
    \ces_0_0_io_ins_left[0] }),
    .io_ins_right({net1084,
    net1083,
    net1082,
    net1081,
    net1079,
    net1078,
    net1077,
    net1076,
    net1075,
    net1074,
    net1073,
    net1072,
    net1071,
    net1070,
    net1068,
    net1067,
    net1066,
    net1065,
    net1064,
    net1063,
    net1062,
    net1061,
    net1060,
    net1059,
    net1057,
    net1056,
    net1055,
    net1054,
    net1053,
    net1052,
    net1051,
    net1050,
    net1049,
    net1048,
    net1046,
    net1045,
    net1044,
    net1043,
    net1042,
    net1041,
    net1040,
    net1039,
    net1038,
    net1037,
    net1035,
    net1034,
    net1033,
    net1032,
    net1031,
    net1030,
    net1029,
    net1028,
    net1027,
    net1026,
    net1088,
    net1087,
    net1086,
    net1085,
    net1080,
    net1069,
    net1058,
    net1047,
    net1036,
    net1025}),
    .io_ins_up({net1596,
    net1595,
    net1594,
    net1593,
    net1591,
    net1590,
    net1589,
    net1588,
    net1587,
    net1586,
    net1585,
    net1584,
    net1583,
    net1582,
    net1580,
    net1579,
    net1578,
    net1577,
    net1576,
    net1575,
    net1574,
    net1573,
    net1572,
    net1571,
    net1569,
    net1568,
    net1567,
    net1566,
    net1565,
    net1564,
    net1563,
    net1562,
    net1561,
    net1560,
    net1558,
    net1557,
    net1556,
    net1555,
    net1554,
    net1553,
    net1552,
    net1551,
    net1550,
    net1549,
    net1547,
    net1546,
    net1545,
    net1544,
    net1543,
    net1542,
    net1541,
    net1540,
    net1539,
    net1538,
    net1600,
    net1599,
    net1598,
    net1597,
    net1592,
    net1581,
    net1570,
    net1559,
    net1548,
    net1537}),
    .io_outs_down({net2172,
    net2171,
    net2170,
    net2169,
    net2167,
    net2166,
    net2165,
    net2164,
    net2163,
    net2162,
    net2161,
    net2160,
    net2159,
    net2158,
    net2156,
    net2155,
    net2154,
    net2153,
    net2152,
    net2151,
    net2150,
    net2149,
    net2148,
    net2147,
    net2145,
    net2144,
    net2143,
    net2142,
    net2141,
    net2140,
    net2139,
    net2138,
    net2137,
    net2136,
    net2134,
    net2133,
    net2132,
    net2131,
    net2130,
    net2129,
    net2128,
    net2127,
    net2126,
    net2125,
    net2123,
    net2122,
    net2121,
    net2120,
    net2119,
    net2118,
    net2117,
    net2116,
    net2115,
    net2114,
    net2176,
    net2175,
    net2174,
    net2173,
    net2168,
    net2157,
    net2146,
    net2135,
    net2124,
    net2113}),
    .io_outs_left({net2684,
    net2683,
    net2682,
    net2681,
    net2679,
    net2678,
    net2677,
    net2676,
    net2675,
    net2674,
    net2673,
    net2672,
    net2671,
    net2670,
    net2668,
    net2667,
    net2666,
    net2665,
    net2664,
    net2663,
    net2662,
    net2661,
    net2660,
    net2659,
    net2657,
    net2656,
    net2655,
    net2654,
    net2653,
    net2652,
    net2651,
    net2650,
    net2649,
    net2648,
    net2646,
    net2645,
    net2644,
    net2643,
    net2642,
    net2641,
    net2640,
    net2639,
    net2638,
    net2637,
    net2635,
    net2634,
    net2633,
    net2632,
    net2631,
    net2630,
    net2629,
    net2628,
    net2627,
    net2626,
    net2688,
    net2687,
    net2686,
    net2685,
    net2680,
    net2669,
    net2658,
    net2647,
    net2636,
    net2625}),
    .io_outs_right({\ces_0_0_io_outs_right[63] ,
    \ces_0_0_io_outs_right[62] ,
    \ces_0_0_io_outs_right[61] ,
    \ces_0_0_io_outs_right[60] ,
    \ces_0_0_io_outs_right[59] ,
    \ces_0_0_io_outs_right[58] ,
    \ces_0_0_io_outs_right[57] ,
    \ces_0_0_io_outs_right[56] ,
    \ces_0_0_io_outs_right[55] ,
    \ces_0_0_io_outs_right[54] ,
    \ces_0_0_io_outs_right[53] ,
    \ces_0_0_io_outs_right[52] ,
    \ces_0_0_io_outs_right[51] ,
    \ces_0_0_io_outs_right[50] ,
    \ces_0_0_io_outs_right[49] ,
    \ces_0_0_io_outs_right[48] ,
    \ces_0_0_io_outs_right[47] ,
    \ces_0_0_io_outs_right[46] ,
    \ces_0_0_io_outs_right[45] ,
    \ces_0_0_io_outs_right[44] ,
    \ces_0_0_io_outs_right[43] ,
    \ces_0_0_io_outs_right[42] ,
    \ces_0_0_io_outs_right[41] ,
    \ces_0_0_io_outs_right[40] ,
    \ces_0_0_io_outs_right[39] ,
    \ces_0_0_io_outs_right[38] ,
    \ces_0_0_io_outs_right[37] ,
    \ces_0_0_io_outs_right[36] ,
    \ces_0_0_io_outs_right[35] ,
    \ces_0_0_io_outs_right[34] ,
    \ces_0_0_io_outs_right[33] ,
    \ces_0_0_io_outs_right[32] ,
    \ces_0_0_io_outs_right[31] ,
    \ces_0_0_io_outs_right[30] ,
    \ces_0_0_io_outs_right[29] ,
    \ces_0_0_io_outs_right[28] ,
    \ces_0_0_io_outs_right[27] ,
    \ces_0_0_io_outs_right[26] ,
    \ces_0_0_io_outs_right[25] ,
    \ces_0_0_io_outs_right[24] ,
    \ces_0_0_io_outs_right[23] ,
    \ces_0_0_io_outs_right[22] ,
    \ces_0_0_io_outs_right[21] ,
    \ces_0_0_io_outs_right[20] ,
    \ces_0_0_io_outs_right[19] ,
    \ces_0_0_io_outs_right[18] ,
    \ces_0_0_io_outs_right[17] ,
    \ces_0_0_io_outs_right[16] ,
    \ces_0_0_io_outs_right[15] ,
    \ces_0_0_io_outs_right[14] ,
    \ces_0_0_io_outs_right[13] ,
    \ces_0_0_io_outs_right[12] ,
    \ces_0_0_io_outs_right[11] ,
    \ces_0_0_io_outs_right[10] ,
    \ces_0_0_io_outs_right[9] ,
    \ces_0_0_io_outs_right[8] ,
    \ces_0_0_io_outs_right[7] ,
    \ces_0_0_io_outs_right[6] ,
    \ces_0_0_io_outs_right[5] ,
    \ces_0_0_io_outs_right[4] ,
    \ces_0_0_io_outs_right[3] ,
    \ces_0_0_io_outs_right[2] ,
    \ces_0_0_io_outs_right[1] ,
    \ces_0_0_io_outs_right[0] }),
    .io_outs_up({\ces_0_0_io_outs_up[63] ,
    \ces_0_0_io_outs_up[62] ,
    \ces_0_0_io_outs_up[61] ,
    \ces_0_0_io_outs_up[60] ,
    \ces_0_0_io_outs_up[59] ,
    \ces_0_0_io_outs_up[58] ,
    \ces_0_0_io_outs_up[57] ,
    \ces_0_0_io_outs_up[56] ,
    \ces_0_0_io_outs_up[55] ,
    \ces_0_0_io_outs_up[54] ,
    \ces_0_0_io_outs_up[53] ,
    \ces_0_0_io_outs_up[52] ,
    \ces_0_0_io_outs_up[51] ,
    \ces_0_0_io_outs_up[50] ,
    \ces_0_0_io_outs_up[49] ,
    \ces_0_0_io_outs_up[48] ,
    \ces_0_0_io_outs_up[47] ,
    \ces_0_0_io_outs_up[46] ,
    \ces_0_0_io_outs_up[45] ,
    \ces_0_0_io_outs_up[44] ,
    \ces_0_0_io_outs_up[43] ,
    \ces_0_0_io_outs_up[42] ,
    \ces_0_0_io_outs_up[41] ,
    \ces_0_0_io_outs_up[40] ,
    \ces_0_0_io_outs_up[39] ,
    \ces_0_0_io_outs_up[38] ,
    \ces_0_0_io_outs_up[37] ,
    \ces_0_0_io_outs_up[36] ,
    \ces_0_0_io_outs_up[35] ,
    \ces_0_0_io_outs_up[34] ,
    \ces_0_0_io_outs_up[33] ,
    \ces_0_0_io_outs_up[32] ,
    \ces_0_0_io_outs_up[31] ,
    \ces_0_0_io_outs_up[30] ,
    \ces_0_0_io_outs_up[29] ,
    \ces_0_0_io_outs_up[28] ,
    \ces_0_0_io_outs_up[27] ,
    \ces_0_0_io_outs_up[26] ,
    \ces_0_0_io_outs_up[25] ,
    \ces_0_0_io_outs_up[24] ,
    \ces_0_0_io_outs_up[23] ,
    \ces_0_0_io_outs_up[22] ,
    \ces_0_0_io_outs_up[21] ,
    \ces_0_0_io_outs_up[20] ,
    \ces_0_0_io_outs_up[19] ,
    \ces_0_0_io_outs_up[18] ,
    \ces_0_0_io_outs_up[17] ,
    \ces_0_0_io_outs_up[16] ,
    \ces_0_0_io_outs_up[15] ,
    \ces_0_0_io_outs_up[14] ,
    \ces_0_0_io_outs_up[13] ,
    \ces_0_0_io_outs_up[12] ,
    \ces_0_0_io_outs_up[11] ,
    \ces_0_0_io_outs_up[10] ,
    \ces_0_0_io_outs_up[9] ,
    \ces_0_0_io_outs_up[8] ,
    \ces_0_0_io_outs_up[7] ,
    \ces_0_0_io_outs_up[6] ,
    \ces_0_0_io_outs_up[5] ,
    \ces_0_0_io_outs_up[4] ,
    \ces_0_0_io_outs_up[3] ,
    \ces_0_0_io_outs_up[2] ,
    \ces_0_0_io_outs_up[1] ,
    \ces_0_0_io_outs_up[0] }));
 Element ces_0_1 (.clock(clknet_3_0_0_clock),
    .io_lsbIns_1(ces_0_0_io_lsbOuts_1),
    .io_lsbIns_2(ces_0_0_io_lsbOuts_2),
    .io_lsbIns_3(ces_0_0_io_lsbOuts_3),
    .io_lsbIns_4(ces_0_0_io_lsbOuts_4),
    .io_lsbIns_5(ces_0_0_io_lsbOuts_5),
    .io_lsbIns_6(ces_0_0_io_lsbOuts_6),
    .io_lsbIns_7(ces_0_0_io_lsbOuts_7),
    .io_lsbOuts_0(ces_0_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_1_io_lsbOuts_7),
    .io_ins_down({\ces_0_1_io_ins_down[63] ,
    \ces_0_1_io_ins_down[62] ,
    \ces_0_1_io_ins_down[61] ,
    \ces_0_1_io_ins_down[60] ,
    \ces_0_1_io_ins_down[59] ,
    \ces_0_1_io_ins_down[58] ,
    \ces_0_1_io_ins_down[57] ,
    \ces_0_1_io_ins_down[56] ,
    \ces_0_1_io_ins_down[55] ,
    \ces_0_1_io_ins_down[54] ,
    \ces_0_1_io_ins_down[53] ,
    \ces_0_1_io_ins_down[52] ,
    \ces_0_1_io_ins_down[51] ,
    \ces_0_1_io_ins_down[50] ,
    \ces_0_1_io_ins_down[49] ,
    \ces_0_1_io_ins_down[48] ,
    \ces_0_1_io_ins_down[47] ,
    \ces_0_1_io_ins_down[46] ,
    \ces_0_1_io_ins_down[45] ,
    \ces_0_1_io_ins_down[44] ,
    \ces_0_1_io_ins_down[43] ,
    \ces_0_1_io_ins_down[42] ,
    \ces_0_1_io_ins_down[41] ,
    \ces_0_1_io_ins_down[40] ,
    \ces_0_1_io_ins_down[39] ,
    \ces_0_1_io_ins_down[38] ,
    \ces_0_1_io_ins_down[37] ,
    \ces_0_1_io_ins_down[36] ,
    \ces_0_1_io_ins_down[35] ,
    \ces_0_1_io_ins_down[34] ,
    \ces_0_1_io_ins_down[33] ,
    \ces_0_1_io_ins_down[32] ,
    \ces_0_1_io_ins_down[31] ,
    \ces_0_1_io_ins_down[30] ,
    \ces_0_1_io_ins_down[29] ,
    \ces_0_1_io_ins_down[28] ,
    \ces_0_1_io_ins_down[27] ,
    \ces_0_1_io_ins_down[26] ,
    \ces_0_1_io_ins_down[25] ,
    \ces_0_1_io_ins_down[24] ,
    \ces_0_1_io_ins_down[23] ,
    \ces_0_1_io_ins_down[22] ,
    \ces_0_1_io_ins_down[21] ,
    \ces_0_1_io_ins_down[20] ,
    \ces_0_1_io_ins_down[19] ,
    \ces_0_1_io_ins_down[18] ,
    \ces_0_1_io_ins_down[17] ,
    \ces_0_1_io_ins_down[16] ,
    \ces_0_1_io_ins_down[15] ,
    \ces_0_1_io_ins_down[14] ,
    \ces_0_1_io_ins_down[13] ,
    \ces_0_1_io_ins_down[12] ,
    \ces_0_1_io_ins_down[11] ,
    \ces_0_1_io_ins_down[10] ,
    \ces_0_1_io_ins_down[9] ,
    \ces_0_1_io_ins_down[8] ,
    \ces_0_1_io_ins_down[7] ,
    \ces_0_1_io_ins_down[6] ,
    \ces_0_1_io_ins_down[5] ,
    \ces_0_1_io_ins_down[4] ,
    \ces_0_1_io_ins_down[3] ,
    \ces_0_1_io_ins_down[2] ,
    \ces_0_1_io_ins_down[1] ,
    \ces_0_1_io_ins_down[0] }),
    .io_ins_left({\ces_0_1_io_ins_left[63] ,
    \ces_0_1_io_ins_left[62] ,
    \ces_0_1_io_ins_left[61] ,
    \ces_0_1_io_ins_left[60] ,
    \ces_0_1_io_ins_left[59] ,
    \ces_0_1_io_ins_left[58] ,
    \ces_0_1_io_ins_left[57] ,
    \ces_0_1_io_ins_left[56] ,
    \ces_0_1_io_ins_left[55] ,
    \ces_0_1_io_ins_left[54] ,
    \ces_0_1_io_ins_left[53] ,
    \ces_0_1_io_ins_left[52] ,
    \ces_0_1_io_ins_left[51] ,
    \ces_0_1_io_ins_left[50] ,
    \ces_0_1_io_ins_left[49] ,
    \ces_0_1_io_ins_left[48] ,
    \ces_0_1_io_ins_left[47] ,
    \ces_0_1_io_ins_left[46] ,
    \ces_0_1_io_ins_left[45] ,
    \ces_0_1_io_ins_left[44] ,
    \ces_0_1_io_ins_left[43] ,
    \ces_0_1_io_ins_left[42] ,
    \ces_0_1_io_ins_left[41] ,
    \ces_0_1_io_ins_left[40] ,
    \ces_0_1_io_ins_left[39] ,
    \ces_0_1_io_ins_left[38] ,
    \ces_0_1_io_ins_left[37] ,
    \ces_0_1_io_ins_left[36] ,
    \ces_0_1_io_ins_left[35] ,
    \ces_0_1_io_ins_left[34] ,
    \ces_0_1_io_ins_left[33] ,
    \ces_0_1_io_ins_left[32] ,
    \ces_0_1_io_ins_left[31] ,
    \ces_0_1_io_ins_left[30] ,
    \ces_0_1_io_ins_left[29] ,
    \ces_0_1_io_ins_left[28] ,
    \ces_0_1_io_ins_left[27] ,
    \ces_0_1_io_ins_left[26] ,
    \ces_0_1_io_ins_left[25] ,
    \ces_0_1_io_ins_left[24] ,
    \ces_0_1_io_ins_left[23] ,
    \ces_0_1_io_ins_left[22] ,
    \ces_0_1_io_ins_left[21] ,
    \ces_0_1_io_ins_left[20] ,
    \ces_0_1_io_ins_left[19] ,
    \ces_0_1_io_ins_left[18] ,
    \ces_0_1_io_ins_left[17] ,
    \ces_0_1_io_ins_left[16] ,
    \ces_0_1_io_ins_left[15] ,
    \ces_0_1_io_ins_left[14] ,
    \ces_0_1_io_ins_left[13] ,
    \ces_0_1_io_ins_left[12] ,
    \ces_0_1_io_ins_left[11] ,
    \ces_0_1_io_ins_left[10] ,
    \ces_0_1_io_ins_left[9] ,
    \ces_0_1_io_ins_left[8] ,
    \ces_0_1_io_ins_left[7] ,
    \ces_0_1_io_ins_left[6] ,
    \ces_0_1_io_ins_left[5] ,
    \ces_0_1_io_ins_left[4] ,
    \ces_0_1_io_ins_left[3] ,
    \ces_0_1_io_ins_left[2] ,
    \ces_0_1_io_ins_left[1] ,
    \ces_0_1_io_ins_left[0] }),
    .io_ins_right({\ces_0_0_io_outs_right[63] ,
    \ces_0_0_io_outs_right[62] ,
    \ces_0_0_io_outs_right[61] ,
    \ces_0_0_io_outs_right[60] ,
    \ces_0_0_io_outs_right[59] ,
    \ces_0_0_io_outs_right[58] ,
    \ces_0_0_io_outs_right[57] ,
    \ces_0_0_io_outs_right[56] ,
    \ces_0_0_io_outs_right[55] ,
    \ces_0_0_io_outs_right[54] ,
    \ces_0_0_io_outs_right[53] ,
    \ces_0_0_io_outs_right[52] ,
    \ces_0_0_io_outs_right[51] ,
    \ces_0_0_io_outs_right[50] ,
    \ces_0_0_io_outs_right[49] ,
    \ces_0_0_io_outs_right[48] ,
    \ces_0_0_io_outs_right[47] ,
    \ces_0_0_io_outs_right[46] ,
    \ces_0_0_io_outs_right[45] ,
    \ces_0_0_io_outs_right[44] ,
    \ces_0_0_io_outs_right[43] ,
    \ces_0_0_io_outs_right[42] ,
    \ces_0_0_io_outs_right[41] ,
    \ces_0_0_io_outs_right[40] ,
    \ces_0_0_io_outs_right[39] ,
    \ces_0_0_io_outs_right[38] ,
    \ces_0_0_io_outs_right[37] ,
    \ces_0_0_io_outs_right[36] ,
    \ces_0_0_io_outs_right[35] ,
    \ces_0_0_io_outs_right[34] ,
    \ces_0_0_io_outs_right[33] ,
    \ces_0_0_io_outs_right[32] ,
    \ces_0_0_io_outs_right[31] ,
    \ces_0_0_io_outs_right[30] ,
    \ces_0_0_io_outs_right[29] ,
    \ces_0_0_io_outs_right[28] ,
    \ces_0_0_io_outs_right[27] ,
    \ces_0_0_io_outs_right[26] ,
    \ces_0_0_io_outs_right[25] ,
    \ces_0_0_io_outs_right[24] ,
    \ces_0_0_io_outs_right[23] ,
    \ces_0_0_io_outs_right[22] ,
    \ces_0_0_io_outs_right[21] ,
    \ces_0_0_io_outs_right[20] ,
    \ces_0_0_io_outs_right[19] ,
    \ces_0_0_io_outs_right[18] ,
    \ces_0_0_io_outs_right[17] ,
    \ces_0_0_io_outs_right[16] ,
    \ces_0_0_io_outs_right[15] ,
    \ces_0_0_io_outs_right[14] ,
    \ces_0_0_io_outs_right[13] ,
    \ces_0_0_io_outs_right[12] ,
    \ces_0_0_io_outs_right[11] ,
    \ces_0_0_io_outs_right[10] ,
    \ces_0_0_io_outs_right[9] ,
    \ces_0_0_io_outs_right[8] ,
    \ces_0_0_io_outs_right[7] ,
    \ces_0_0_io_outs_right[6] ,
    \ces_0_0_io_outs_right[5] ,
    \ces_0_0_io_outs_right[4] ,
    \ces_0_0_io_outs_right[3] ,
    \ces_0_0_io_outs_right[2] ,
    \ces_0_0_io_outs_right[1] ,
    \ces_0_0_io_outs_right[0] }),
    .io_ins_up({net1660,
    net1659,
    net1658,
    net1657,
    net1655,
    net1654,
    net1653,
    net1652,
    net1651,
    net1650,
    net1649,
    net1648,
    net1647,
    net1646,
    net1644,
    net1643,
    net1642,
    net1641,
    net1640,
    net1639,
    net1638,
    net1637,
    net1636,
    net1635,
    net1633,
    net1632,
    net1631,
    net1630,
    net1629,
    net1628,
    net1627,
    net1626,
    net1625,
    net1624,
    net1622,
    net1621,
    net1620,
    net1619,
    net1618,
    net1617,
    net1616,
    net1615,
    net1614,
    net1613,
    net1611,
    net1610,
    net1609,
    net1608,
    net1607,
    net1606,
    net1605,
    net1604,
    net1603,
    net1602,
    net1664,
    net1663,
    net1662,
    net1661,
    net1656,
    net1645,
    net1634,
    net1623,
    net1612,
    net1601}),
    .io_outs_down({net2236,
    net2235,
    net2234,
    net2233,
    net2231,
    net2230,
    net2229,
    net2228,
    net2227,
    net2226,
    net2225,
    net2224,
    net2223,
    net2222,
    net2220,
    net2219,
    net2218,
    net2217,
    net2216,
    net2215,
    net2214,
    net2213,
    net2212,
    net2211,
    net2209,
    net2208,
    net2207,
    net2206,
    net2205,
    net2204,
    net2203,
    net2202,
    net2201,
    net2200,
    net2198,
    net2197,
    net2196,
    net2195,
    net2194,
    net2193,
    net2192,
    net2191,
    net2190,
    net2189,
    net2187,
    net2186,
    net2185,
    net2184,
    net2183,
    net2182,
    net2181,
    net2180,
    net2179,
    net2178,
    net2240,
    net2239,
    net2238,
    net2237,
    net2232,
    net2221,
    net2210,
    net2199,
    net2188,
    net2177}),
    .io_outs_left({\ces_0_0_io_ins_left[63] ,
    \ces_0_0_io_ins_left[62] ,
    \ces_0_0_io_ins_left[61] ,
    \ces_0_0_io_ins_left[60] ,
    \ces_0_0_io_ins_left[59] ,
    \ces_0_0_io_ins_left[58] ,
    \ces_0_0_io_ins_left[57] ,
    \ces_0_0_io_ins_left[56] ,
    \ces_0_0_io_ins_left[55] ,
    \ces_0_0_io_ins_left[54] ,
    \ces_0_0_io_ins_left[53] ,
    \ces_0_0_io_ins_left[52] ,
    \ces_0_0_io_ins_left[51] ,
    \ces_0_0_io_ins_left[50] ,
    \ces_0_0_io_ins_left[49] ,
    \ces_0_0_io_ins_left[48] ,
    \ces_0_0_io_ins_left[47] ,
    \ces_0_0_io_ins_left[46] ,
    \ces_0_0_io_ins_left[45] ,
    \ces_0_0_io_ins_left[44] ,
    \ces_0_0_io_ins_left[43] ,
    \ces_0_0_io_ins_left[42] ,
    \ces_0_0_io_ins_left[41] ,
    \ces_0_0_io_ins_left[40] ,
    \ces_0_0_io_ins_left[39] ,
    \ces_0_0_io_ins_left[38] ,
    \ces_0_0_io_ins_left[37] ,
    \ces_0_0_io_ins_left[36] ,
    \ces_0_0_io_ins_left[35] ,
    \ces_0_0_io_ins_left[34] ,
    \ces_0_0_io_ins_left[33] ,
    \ces_0_0_io_ins_left[32] ,
    \ces_0_0_io_ins_left[31] ,
    \ces_0_0_io_ins_left[30] ,
    \ces_0_0_io_ins_left[29] ,
    \ces_0_0_io_ins_left[28] ,
    \ces_0_0_io_ins_left[27] ,
    \ces_0_0_io_ins_left[26] ,
    \ces_0_0_io_ins_left[25] ,
    \ces_0_0_io_ins_left[24] ,
    \ces_0_0_io_ins_left[23] ,
    \ces_0_0_io_ins_left[22] ,
    \ces_0_0_io_ins_left[21] ,
    \ces_0_0_io_ins_left[20] ,
    \ces_0_0_io_ins_left[19] ,
    \ces_0_0_io_ins_left[18] ,
    \ces_0_0_io_ins_left[17] ,
    \ces_0_0_io_ins_left[16] ,
    \ces_0_0_io_ins_left[15] ,
    \ces_0_0_io_ins_left[14] ,
    \ces_0_0_io_ins_left[13] ,
    \ces_0_0_io_ins_left[12] ,
    \ces_0_0_io_ins_left[11] ,
    \ces_0_0_io_ins_left[10] ,
    \ces_0_0_io_ins_left[9] ,
    \ces_0_0_io_ins_left[8] ,
    \ces_0_0_io_ins_left[7] ,
    \ces_0_0_io_ins_left[6] ,
    \ces_0_0_io_ins_left[5] ,
    \ces_0_0_io_ins_left[4] ,
    \ces_0_0_io_ins_left[3] ,
    \ces_0_0_io_ins_left[2] ,
    \ces_0_0_io_ins_left[1] ,
    \ces_0_0_io_ins_left[0] }),
    .io_outs_right({\ces_0_1_io_outs_right[63] ,
    \ces_0_1_io_outs_right[62] ,
    \ces_0_1_io_outs_right[61] ,
    \ces_0_1_io_outs_right[60] ,
    \ces_0_1_io_outs_right[59] ,
    \ces_0_1_io_outs_right[58] ,
    \ces_0_1_io_outs_right[57] ,
    \ces_0_1_io_outs_right[56] ,
    \ces_0_1_io_outs_right[55] ,
    \ces_0_1_io_outs_right[54] ,
    \ces_0_1_io_outs_right[53] ,
    \ces_0_1_io_outs_right[52] ,
    \ces_0_1_io_outs_right[51] ,
    \ces_0_1_io_outs_right[50] ,
    \ces_0_1_io_outs_right[49] ,
    \ces_0_1_io_outs_right[48] ,
    \ces_0_1_io_outs_right[47] ,
    \ces_0_1_io_outs_right[46] ,
    \ces_0_1_io_outs_right[45] ,
    \ces_0_1_io_outs_right[44] ,
    \ces_0_1_io_outs_right[43] ,
    \ces_0_1_io_outs_right[42] ,
    \ces_0_1_io_outs_right[41] ,
    \ces_0_1_io_outs_right[40] ,
    \ces_0_1_io_outs_right[39] ,
    \ces_0_1_io_outs_right[38] ,
    \ces_0_1_io_outs_right[37] ,
    \ces_0_1_io_outs_right[36] ,
    \ces_0_1_io_outs_right[35] ,
    \ces_0_1_io_outs_right[34] ,
    \ces_0_1_io_outs_right[33] ,
    \ces_0_1_io_outs_right[32] ,
    \ces_0_1_io_outs_right[31] ,
    \ces_0_1_io_outs_right[30] ,
    \ces_0_1_io_outs_right[29] ,
    \ces_0_1_io_outs_right[28] ,
    \ces_0_1_io_outs_right[27] ,
    \ces_0_1_io_outs_right[26] ,
    \ces_0_1_io_outs_right[25] ,
    \ces_0_1_io_outs_right[24] ,
    \ces_0_1_io_outs_right[23] ,
    \ces_0_1_io_outs_right[22] ,
    \ces_0_1_io_outs_right[21] ,
    \ces_0_1_io_outs_right[20] ,
    \ces_0_1_io_outs_right[19] ,
    \ces_0_1_io_outs_right[18] ,
    \ces_0_1_io_outs_right[17] ,
    \ces_0_1_io_outs_right[16] ,
    \ces_0_1_io_outs_right[15] ,
    \ces_0_1_io_outs_right[14] ,
    \ces_0_1_io_outs_right[13] ,
    \ces_0_1_io_outs_right[12] ,
    \ces_0_1_io_outs_right[11] ,
    \ces_0_1_io_outs_right[10] ,
    \ces_0_1_io_outs_right[9] ,
    \ces_0_1_io_outs_right[8] ,
    \ces_0_1_io_outs_right[7] ,
    \ces_0_1_io_outs_right[6] ,
    \ces_0_1_io_outs_right[5] ,
    \ces_0_1_io_outs_right[4] ,
    \ces_0_1_io_outs_right[3] ,
    \ces_0_1_io_outs_right[2] ,
    \ces_0_1_io_outs_right[1] ,
    \ces_0_1_io_outs_right[0] }),
    .io_outs_up({\ces_0_1_io_outs_up[63] ,
    \ces_0_1_io_outs_up[62] ,
    \ces_0_1_io_outs_up[61] ,
    \ces_0_1_io_outs_up[60] ,
    \ces_0_1_io_outs_up[59] ,
    \ces_0_1_io_outs_up[58] ,
    \ces_0_1_io_outs_up[57] ,
    \ces_0_1_io_outs_up[56] ,
    \ces_0_1_io_outs_up[55] ,
    \ces_0_1_io_outs_up[54] ,
    \ces_0_1_io_outs_up[53] ,
    \ces_0_1_io_outs_up[52] ,
    \ces_0_1_io_outs_up[51] ,
    \ces_0_1_io_outs_up[50] ,
    \ces_0_1_io_outs_up[49] ,
    \ces_0_1_io_outs_up[48] ,
    \ces_0_1_io_outs_up[47] ,
    \ces_0_1_io_outs_up[46] ,
    \ces_0_1_io_outs_up[45] ,
    \ces_0_1_io_outs_up[44] ,
    \ces_0_1_io_outs_up[43] ,
    \ces_0_1_io_outs_up[42] ,
    \ces_0_1_io_outs_up[41] ,
    \ces_0_1_io_outs_up[40] ,
    \ces_0_1_io_outs_up[39] ,
    \ces_0_1_io_outs_up[38] ,
    \ces_0_1_io_outs_up[37] ,
    \ces_0_1_io_outs_up[36] ,
    \ces_0_1_io_outs_up[35] ,
    \ces_0_1_io_outs_up[34] ,
    \ces_0_1_io_outs_up[33] ,
    \ces_0_1_io_outs_up[32] ,
    \ces_0_1_io_outs_up[31] ,
    \ces_0_1_io_outs_up[30] ,
    \ces_0_1_io_outs_up[29] ,
    \ces_0_1_io_outs_up[28] ,
    \ces_0_1_io_outs_up[27] ,
    \ces_0_1_io_outs_up[26] ,
    \ces_0_1_io_outs_up[25] ,
    \ces_0_1_io_outs_up[24] ,
    \ces_0_1_io_outs_up[23] ,
    \ces_0_1_io_outs_up[22] ,
    \ces_0_1_io_outs_up[21] ,
    \ces_0_1_io_outs_up[20] ,
    \ces_0_1_io_outs_up[19] ,
    \ces_0_1_io_outs_up[18] ,
    \ces_0_1_io_outs_up[17] ,
    \ces_0_1_io_outs_up[16] ,
    \ces_0_1_io_outs_up[15] ,
    \ces_0_1_io_outs_up[14] ,
    \ces_0_1_io_outs_up[13] ,
    \ces_0_1_io_outs_up[12] ,
    \ces_0_1_io_outs_up[11] ,
    \ces_0_1_io_outs_up[10] ,
    \ces_0_1_io_outs_up[9] ,
    \ces_0_1_io_outs_up[8] ,
    \ces_0_1_io_outs_up[7] ,
    \ces_0_1_io_outs_up[6] ,
    \ces_0_1_io_outs_up[5] ,
    \ces_0_1_io_outs_up[4] ,
    \ces_0_1_io_outs_up[3] ,
    \ces_0_1_io_outs_up[2] ,
    \ces_0_1_io_outs_up[1] ,
    \ces_0_1_io_outs_up[0] }));
 Element ces_0_2 (.clock(clknet_3_0_0_clock),
    .io_lsbIns_1(ces_0_1_io_lsbOuts_1),
    .io_lsbIns_2(ces_0_1_io_lsbOuts_2),
    .io_lsbIns_3(ces_0_1_io_lsbOuts_3),
    .io_lsbIns_4(ces_0_1_io_lsbOuts_4),
    .io_lsbIns_5(ces_0_1_io_lsbOuts_5),
    .io_lsbIns_6(ces_0_1_io_lsbOuts_6),
    .io_lsbIns_7(ces_0_1_io_lsbOuts_7),
    .io_lsbOuts_0(ces_0_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_2_io_lsbOuts_7),
    .io_ins_down({\ces_0_2_io_ins_down[63] ,
    \ces_0_2_io_ins_down[62] ,
    \ces_0_2_io_ins_down[61] ,
    \ces_0_2_io_ins_down[60] ,
    \ces_0_2_io_ins_down[59] ,
    \ces_0_2_io_ins_down[58] ,
    \ces_0_2_io_ins_down[57] ,
    \ces_0_2_io_ins_down[56] ,
    \ces_0_2_io_ins_down[55] ,
    \ces_0_2_io_ins_down[54] ,
    \ces_0_2_io_ins_down[53] ,
    \ces_0_2_io_ins_down[52] ,
    \ces_0_2_io_ins_down[51] ,
    \ces_0_2_io_ins_down[50] ,
    \ces_0_2_io_ins_down[49] ,
    \ces_0_2_io_ins_down[48] ,
    \ces_0_2_io_ins_down[47] ,
    \ces_0_2_io_ins_down[46] ,
    \ces_0_2_io_ins_down[45] ,
    \ces_0_2_io_ins_down[44] ,
    \ces_0_2_io_ins_down[43] ,
    \ces_0_2_io_ins_down[42] ,
    \ces_0_2_io_ins_down[41] ,
    \ces_0_2_io_ins_down[40] ,
    \ces_0_2_io_ins_down[39] ,
    \ces_0_2_io_ins_down[38] ,
    \ces_0_2_io_ins_down[37] ,
    \ces_0_2_io_ins_down[36] ,
    \ces_0_2_io_ins_down[35] ,
    \ces_0_2_io_ins_down[34] ,
    \ces_0_2_io_ins_down[33] ,
    \ces_0_2_io_ins_down[32] ,
    \ces_0_2_io_ins_down[31] ,
    \ces_0_2_io_ins_down[30] ,
    \ces_0_2_io_ins_down[29] ,
    \ces_0_2_io_ins_down[28] ,
    \ces_0_2_io_ins_down[27] ,
    \ces_0_2_io_ins_down[26] ,
    \ces_0_2_io_ins_down[25] ,
    \ces_0_2_io_ins_down[24] ,
    \ces_0_2_io_ins_down[23] ,
    \ces_0_2_io_ins_down[22] ,
    \ces_0_2_io_ins_down[21] ,
    \ces_0_2_io_ins_down[20] ,
    \ces_0_2_io_ins_down[19] ,
    \ces_0_2_io_ins_down[18] ,
    \ces_0_2_io_ins_down[17] ,
    \ces_0_2_io_ins_down[16] ,
    \ces_0_2_io_ins_down[15] ,
    \ces_0_2_io_ins_down[14] ,
    \ces_0_2_io_ins_down[13] ,
    \ces_0_2_io_ins_down[12] ,
    \ces_0_2_io_ins_down[11] ,
    \ces_0_2_io_ins_down[10] ,
    \ces_0_2_io_ins_down[9] ,
    \ces_0_2_io_ins_down[8] ,
    \ces_0_2_io_ins_down[7] ,
    \ces_0_2_io_ins_down[6] ,
    \ces_0_2_io_ins_down[5] ,
    \ces_0_2_io_ins_down[4] ,
    \ces_0_2_io_ins_down[3] ,
    \ces_0_2_io_ins_down[2] ,
    \ces_0_2_io_ins_down[1] ,
    \ces_0_2_io_ins_down[0] }),
    .io_ins_left({\ces_0_2_io_ins_left[63] ,
    \ces_0_2_io_ins_left[62] ,
    \ces_0_2_io_ins_left[61] ,
    \ces_0_2_io_ins_left[60] ,
    \ces_0_2_io_ins_left[59] ,
    \ces_0_2_io_ins_left[58] ,
    \ces_0_2_io_ins_left[57] ,
    \ces_0_2_io_ins_left[56] ,
    \ces_0_2_io_ins_left[55] ,
    \ces_0_2_io_ins_left[54] ,
    \ces_0_2_io_ins_left[53] ,
    \ces_0_2_io_ins_left[52] ,
    \ces_0_2_io_ins_left[51] ,
    \ces_0_2_io_ins_left[50] ,
    \ces_0_2_io_ins_left[49] ,
    \ces_0_2_io_ins_left[48] ,
    \ces_0_2_io_ins_left[47] ,
    \ces_0_2_io_ins_left[46] ,
    \ces_0_2_io_ins_left[45] ,
    \ces_0_2_io_ins_left[44] ,
    \ces_0_2_io_ins_left[43] ,
    \ces_0_2_io_ins_left[42] ,
    \ces_0_2_io_ins_left[41] ,
    \ces_0_2_io_ins_left[40] ,
    \ces_0_2_io_ins_left[39] ,
    \ces_0_2_io_ins_left[38] ,
    \ces_0_2_io_ins_left[37] ,
    \ces_0_2_io_ins_left[36] ,
    \ces_0_2_io_ins_left[35] ,
    \ces_0_2_io_ins_left[34] ,
    \ces_0_2_io_ins_left[33] ,
    \ces_0_2_io_ins_left[32] ,
    \ces_0_2_io_ins_left[31] ,
    \ces_0_2_io_ins_left[30] ,
    \ces_0_2_io_ins_left[29] ,
    \ces_0_2_io_ins_left[28] ,
    \ces_0_2_io_ins_left[27] ,
    \ces_0_2_io_ins_left[26] ,
    \ces_0_2_io_ins_left[25] ,
    \ces_0_2_io_ins_left[24] ,
    \ces_0_2_io_ins_left[23] ,
    \ces_0_2_io_ins_left[22] ,
    \ces_0_2_io_ins_left[21] ,
    \ces_0_2_io_ins_left[20] ,
    \ces_0_2_io_ins_left[19] ,
    \ces_0_2_io_ins_left[18] ,
    \ces_0_2_io_ins_left[17] ,
    \ces_0_2_io_ins_left[16] ,
    \ces_0_2_io_ins_left[15] ,
    \ces_0_2_io_ins_left[14] ,
    \ces_0_2_io_ins_left[13] ,
    \ces_0_2_io_ins_left[12] ,
    \ces_0_2_io_ins_left[11] ,
    \ces_0_2_io_ins_left[10] ,
    \ces_0_2_io_ins_left[9] ,
    \ces_0_2_io_ins_left[8] ,
    \ces_0_2_io_ins_left[7] ,
    \ces_0_2_io_ins_left[6] ,
    \ces_0_2_io_ins_left[5] ,
    \ces_0_2_io_ins_left[4] ,
    \ces_0_2_io_ins_left[3] ,
    \ces_0_2_io_ins_left[2] ,
    \ces_0_2_io_ins_left[1] ,
    \ces_0_2_io_ins_left[0] }),
    .io_ins_right({\ces_0_1_io_outs_right[63] ,
    \ces_0_1_io_outs_right[62] ,
    \ces_0_1_io_outs_right[61] ,
    \ces_0_1_io_outs_right[60] ,
    \ces_0_1_io_outs_right[59] ,
    \ces_0_1_io_outs_right[58] ,
    \ces_0_1_io_outs_right[57] ,
    \ces_0_1_io_outs_right[56] ,
    \ces_0_1_io_outs_right[55] ,
    \ces_0_1_io_outs_right[54] ,
    \ces_0_1_io_outs_right[53] ,
    \ces_0_1_io_outs_right[52] ,
    \ces_0_1_io_outs_right[51] ,
    \ces_0_1_io_outs_right[50] ,
    \ces_0_1_io_outs_right[49] ,
    \ces_0_1_io_outs_right[48] ,
    \ces_0_1_io_outs_right[47] ,
    \ces_0_1_io_outs_right[46] ,
    \ces_0_1_io_outs_right[45] ,
    \ces_0_1_io_outs_right[44] ,
    \ces_0_1_io_outs_right[43] ,
    \ces_0_1_io_outs_right[42] ,
    \ces_0_1_io_outs_right[41] ,
    \ces_0_1_io_outs_right[40] ,
    \ces_0_1_io_outs_right[39] ,
    \ces_0_1_io_outs_right[38] ,
    \ces_0_1_io_outs_right[37] ,
    \ces_0_1_io_outs_right[36] ,
    \ces_0_1_io_outs_right[35] ,
    \ces_0_1_io_outs_right[34] ,
    \ces_0_1_io_outs_right[33] ,
    \ces_0_1_io_outs_right[32] ,
    \ces_0_1_io_outs_right[31] ,
    \ces_0_1_io_outs_right[30] ,
    \ces_0_1_io_outs_right[29] ,
    \ces_0_1_io_outs_right[28] ,
    \ces_0_1_io_outs_right[27] ,
    \ces_0_1_io_outs_right[26] ,
    \ces_0_1_io_outs_right[25] ,
    \ces_0_1_io_outs_right[24] ,
    \ces_0_1_io_outs_right[23] ,
    \ces_0_1_io_outs_right[22] ,
    \ces_0_1_io_outs_right[21] ,
    \ces_0_1_io_outs_right[20] ,
    \ces_0_1_io_outs_right[19] ,
    \ces_0_1_io_outs_right[18] ,
    \ces_0_1_io_outs_right[17] ,
    \ces_0_1_io_outs_right[16] ,
    \ces_0_1_io_outs_right[15] ,
    \ces_0_1_io_outs_right[14] ,
    \ces_0_1_io_outs_right[13] ,
    \ces_0_1_io_outs_right[12] ,
    \ces_0_1_io_outs_right[11] ,
    \ces_0_1_io_outs_right[10] ,
    \ces_0_1_io_outs_right[9] ,
    \ces_0_1_io_outs_right[8] ,
    \ces_0_1_io_outs_right[7] ,
    \ces_0_1_io_outs_right[6] ,
    \ces_0_1_io_outs_right[5] ,
    \ces_0_1_io_outs_right[4] ,
    \ces_0_1_io_outs_right[3] ,
    \ces_0_1_io_outs_right[2] ,
    \ces_0_1_io_outs_right[1] ,
    \ces_0_1_io_outs_right[0] }),
    .io_ins_up({net1724,
    net1723,
    net1722,
    net1721,
    net1719,
    net1718,
    net1717,
    net1716,
    net1715,
    net1714,
    net1713,
    net1712,
    net1711,
    net1710,
    net1708,
    net1707,
    net1706,
    net1705,
    net1704,
    net1703,
    net1702,
    net1701,
    net1700,
    net1699,
    net1697,
    net1696,
    net1695,
    net1694,
    net1693,
    net1692,
    net1691,
    net1690,
    net1689,
    net1688,
    net1686,
    net1685,
    net1684,
    net1683,
    net1682,
    net1681,
    net1680,
    net1679,
    net1678,
    net1677,
    net1675,
    net1674,
    net1673,
    net1672,
    net1671,
    net1670,
    net1669,
    net1668,
    net1667,
    net1666,
    net1728,
    net1727,
    net1726,
    net1725,
    net1720,
    net1709,
    net1698,
    net1687,
    net1676,
    net1665}),
    .io_outs_down({net2300,
    net2299,
    net2298,
    net2297,
    net2295,
    net2294,
    net2293,
    net2292,
    net2291,
    net2290,
    net2289,
    net2288,
    net2287,
    net2286,
    net2284,
    net2283,
    net2282,
    net2281,
    net2280,
    net2279,
    net2278,
    net2277,
    net2276,
    net2275,
    net2273,
    net2272,
    net2271,
    net2270,
    net2269,
    net2268,
    net2267,
    net2266,
    net2265,
    net2264,
    net2262,
    net2261,
    net2260,
    net2259,
    net2258,
    net2257,
    net2256,
    net2255,
    net2254,
    net2253,
    net2251,
    net2250,
    net2249,
    net2248,
    net2247,
    net2246,
    net2245,
    net2244,
    net2243,
    net2242,
    net2304,
    net2303,
    net2302,
    net2301,
    net2296,
    net2285,
    net2274,
    net2263,
    net2252,
    net2241}),
    .io_outs_left({\ces_0_1_io_ins_left[63] ,
    \ces_0_1_io_ins_left[62] ,
    \ces_0_1_io_ins_left[61] ,
    \ces_0_1_io_ins_left[60] ,
    \ces_0_1_io_ins_left[59] ,
    \ces_0_1_io_ins_left[58] ,
    \ces_0_1_io_ins_left[57] ,
    \ces_0_1_io_ins_left[56] ,
    \ces_0_1_io_ins_left[55] ,
    \ces_0_1_io_ins_left[54] ,
    \ces_0_1_io_ins_left[53] ,
    \ces_0_1_io_ins_left[52] ,
    \ces_0_1_io_ins_left[51] ,
    \ces_0_1_io_ins_left[50] ,
    \ces_0_1_io_ins_left[49] ,
    \ces_0_1_io_ins_left[48] ,
    \ces_0_1_io_ins_left[47] ,
    \ces_0_1_io_ins_left[46] ,
    \ces_0_1_io_ins_left[45] ,
    \ces_0_1_io_ins_left[44] ,
    \ces_0_1_io_ins_left[43] ,
    \ces_0_1_io_ins_left[42] ,
    \ces_0_1_io_ins_left[41] ,
    \ces_0_1_io_ins_left[40] ,
    \ces_0_1_io_ins_left[39] ,
    \ces_0_1_io_ins_left[38] ,
    \ces_0_1_io_ins_left[37] ,
    \ces_0_1_io_ins_left[36] ,
    \ces_0_1_io_ins_left[35] ,
    \ces_0_1_io_ins_left[34] ,
    \ces_0_1_io_ins_left[33] ,
    \ces_0_1_io_ins_left[32] ,
    \ces_0_1_io_ins_left[31] ,
    \ces_0_1_io_ins_left[30] ,
    \ces_0_1_io_ins_left[29] ,
    \ces_0_1_io_ins_left[28] ,
    \ces_0_1_io_ins_left[27] ,
    \ces_0_1_io_ins_left[26] ,
    \ces_0_1_io_ins_left[25] ,
    \ces_0_1_io_ins_left[24] ,
    \ces_0_1_io_ins_left[23] ,
    \ces_0_1_io_ins_left[22] ,
    \ces_0_1_io_ins_left[21] ,
    \ces_0_1_io_ins_left[20] ,
    \ces_0_1_io_ins_left[19] ,
    \ces_0_1_io_ins_left[18] ,
    \ces_0_1_io_ins_left[17] ,
    \ces_0_1_io_ins_left[16] ,
    \ces_0_1_io_ins_left[15] ,
    \ces_0_1_io_ins_left[14] ,
    \ces_0_1_io_ins_left[13] ,
    \ces_0_1_io_ins_left[12] ,
    \ces_0_1_io_ins_left[11] ,
    \ces_0_1_io_ins_left[10] ,
    \ces_0_1_io_ins_left[9] ,
    \ces_0_1_io_ins_left[8] ,
    \ces_0_1_io_ins_left[7] ,
    \ces_0_1_io_ins_left[6] ,
    \ces_0_1_io_ins_left[5] ,
    \ces_0_1_io_ins_left[4] ,
    \ces_0_1_io_ins_left[3] ,
    \ces_0_1_io_ins_left[2] ,
    \ces_0_1_io_ins_left[1] ,
    \ces_0_1_io_ins_left[0] }),
    .io_outs_right({\ces_0_2_io_outs_right[63] ,
    \ces_0_2_io_outs_right[62] ,
    \ces_0_2_io_outs_right[61] ,
    \ces_0_2_io_outs_right[60] ,
    \ces_0_2_io_outs_right[59] ,
    \ces_0_2_io_outs_right[58] ,
    \ces_0_2_io_outs_right[57] ,
    \ces_0_2_io_outs_right[56] ,
    \ces_0_2_io_outs_right[55] ,
    \ces_0_2_io_outs_right[54] ,
    \ces_0_2_io_outs_right[53] ,
    \ces_0_2_io_outs_right[52] ,
    \ces_0_2_io_outs_right[51] ,
    \ces_0_2_io_outs_right[50] ,
    \ces_0_2_io_outs_right[49] ,
    \ces_0_2_io_outs_right[48] ,
    \ces_0_2_io_outs_right[47] ,
    \ces_0_2_io_outs_right[46] ,
    \ces_0_2_io_outs_right[45] ,
    \ces_0_2_io_outs_right[44] ,
    \ces_0_2_io_outs_right[43] ,
    \ces_0_2_io_outs_right[42] ,
    \ces_0_2_io_outs_right[41] ,
    \ces_0_2_io_outs_right[40] ,
    \ces_0_2_io_outs_right[39] ,
    \ces_0_2_io_outs_right[38] ,
    \ces_0_2_io_outs_right[37] ,
    \ces_0_2_io_outs_right[36] ,
    \ces_0_2_io_outs_right[35] ,
    \ces_0_2_io_outs_right[34] ,
    \ces_0_2_io_outs_right[33] ,
    \ces_0_2_io_outs_right[32] ,
    \ces_0_2_io_outs_right[31] ,
    \ces_0_2_io_outs_right[30] ,
    \ces_0_2_io_outs_right[29] ,
    \ces_0_2_io_outs_right[28] ,
    \ces_0_2_io_outs_right[27] ,
    \ces_0_2_io_outs_right[26] ,
    \ces_0_2_io_outs_right[25] ,
    \ces_0_2_io_outs_right[24] ,
    \ces_0_2_io_outs_right[23] ,
    \ces_0_2_io_outs_right[22] ,
    \ces_0_2_io_outs_right[21] ,
    \ces_0_2_io_outs_right[20] ,
    \ces_0_2_io_outs_right[19] ,
    \ces_0_2_io_outs_right[18] ,
    \ces_0_2_io_outs_right[17] ,
    \ces_0_2_io_outs_right[16] ,
    \ces_0_2_io_outs_right[15] ,
    \ces_0_2_io_outs_right[14] ,
    \ces_0_2_io_outs_right[13] ,
    \ces_0_2_io_outs_right[12] ,
    \ces_0_2_io_outs_right[11] ,
    \ces_0_2_io_outs_right[10] ,
    \ces_0_2_io_outs_right[9] ,
    \ces_0_2_io_outs_right[8] ,
    \ces_0_2_io_outs_right[7] ,
    \ces_0_2_io_outs_right[6] ,
    \ces_0_2_io_outs_right[5] ,
    \ces_0_2_io_outs_right[4] ,
    \ces_0_2_io_outs_right[3] ,
    \ces_0_2_io_outs_right[2] ,
    \ces_0_2_io_outs_right[1] ,
    \ces_0_2_io_outs_right[0] }),
    .io_outs_up({\ces_0_2_io_outs_up[63] ,
    \ces_0_2_io_outs_up[62] ,
    \ces_0_2_io_outs_up[61] ,
    \ces_0_2_io_outs_up[60] ,
    \ces_0_2_io_outs_up[59] ,
    \ces_0_2_io_outs_up[58] ,
    \ces_0_2_io_outs_up[57] ,
    \ces_0_2_io_outs_up[56] ,
    \ces_0_2_io_outs_up[55] ,
    \ces_0_2_io_outs_up[54] ,
    \ces_0_2_io_outs_up[53] ,
    \ces_0_2_io_outs_up[52] ,
    \ces_0_2_io_outs_up[51] ,
    \ces_0_2_io_outs_up[50] ,
    \ces_0_2_io_outs_up[49] ,
    \ces_0_2_io_outs_up[48] ,
    \ces_0_2_io_outs_up[47] ,
    \ces_0_2_io_outs_up[46] ,
    \ces_0_2_io_outs_up[45] ,
    \ces_0_2_io_outs_up[44] ,
    \ces_0_2_io_outs_up[43] ,
    \ces_0_2_io_outs_up[42] ,
    \ces_0_2_io_outs_up[41] ,
    \ces_0_2_io_outs_up[40] ,
    \ces_0_2_io_outs_up[39] ,
    \ces_0_2_io_outs_up[38] ,
    \ces_0_2_io_outs_up[37] ,
    \ces_0_2_io_outs_up[36] ,
    \ces_0_2_io_outs_up[35] ,
    \ces_0_2_io_outs_up[34] ,
    \ces_0_2_io_outs_up[33] ,
    \ces_0_2_io_outs_up[32] ,
    \ces_0_2_io_outs_up[31] ,
    \ces_0_2_io_outs_up[30] ,
    \ces_0_2_io_outs_up[29] ,
    \ces_0_2_io_outs_up[28] ,
    \ces_0_2_io_outs_up[27] ,
    \ces_0_2_io_outs_up[26] ,
    \ces_0_2_io_outs_up[25] ,
    \ces_0_2_io_outs_up[24] ,
    \ces_0_2_io_outs_up[23] ,
    \ces_0_2_io_outs_up[22] ,
    \ces_0_2_io_outs_up[21] ,
    \ces_0_2_io_outs_up[20] ,
    \ces_0_2_io_outs_up[19] ,
    \ces_0_2_io_outs_up[18] ,
    \ces_0_2_io_outs_up[17] ,
    \ces_0_2_io_outs_up[16] ,
    \ces_0_2_io_outs_up[15] ,
    \ces_0_2_io_outs_up[14] ,
    \ces_0_2_io_outs_up[13] ,
    \ces_0_2_io_outs_up[12] ,
    \ces_0_2_io_outs_up[11] ,
    \ces_0_2_io_outs_up[10] ,
    \ces_0_2_io_outs_up[9] ,
    \ces_0_2_io_outs_up[8] ,
    \ces_0_2_io_outs_up[7] ,
    \ces_0_2_io_outs_up[6] ,
    \ces_0_2_io_outs_up[5] ,
    \ces_0_2_io_outs_up[4] ,
    \ces_0_2_io_outs_up[3] ,
    \ces_0_2_io_outs_up[2] ,
    \ces_0_2_io_outs_up[1] ,
    \ces_0_2_io_outs_up[0] }));
 Element ces_0_3 (.clock(clknet_3_0_0_clock),
    .io_lsbIns_1(ces_0_2_io_lsbOuts_1),
    .io_lsbIns_2(ces_0_2_io_lsbOuts_2),
    .io_lsbIns_3(ces_0_2_io_lsbOuts_3),
    .io_lsbIns_4(ces_0_2_io_lsbOuts_4),
    .io_lsbIns_5(ces_0_2_io_lsbOuts_5),
    .io_lsbIns_6(ces_0_2_io_lsbOuts_6),
    .io_lsbIns_7(ces_0_2_io_lsbOuts_7),
    .io_lsbOuts_0(ces_0_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_3_io_lsbOuts_7),
    .io_ins_down({\ces_0_3_io_ins_down[63] ,
    \ces_0_3_io_ins_down[62] ,
    \ces_0_3_io_ins_down[61] ,
    \ces_0_3_io_ins_down[60] ,
    \ces_0_3_io_ins_down[59] ,
    \ces_0_3_io_ins_down[58] ,
    \ces_0_3_io_ins_down[57] ,
    \ces_0_3_io_ins_down[56] ,
    \ces_0_3_io_ins_down[55] ,
    \ces_0_3_io_ins_down[54] ,
    \ces_0_3_io_ins_down[53] ,
    \ces_0_3_io_ins_down[52] ,
    \ces_0_3_io_ins_down[51] ,
    \ces_0_3_io_ins_down[50] ,
    \ces_0_3_io_ins_down[49] ,
    \ces_0_3_io_ins_down[48] ,
    \ces_0_3_io_ins_down[47] ,
    \ces_0_3_io_ins_down[46] ,
    \ces_0_3_io_ins_down[45] ,
    \ces_0_3_io_ins_down[44] ,
    \ces_0_3_io_ins_down[43] ,
    \ces_0_3_io_ins_down[42] ,
    \ces_0_3_io_ins_down[41] ,
    \ces_0_3_io_ins_down[40] ,
    \ces_0_3_io_ins_down[39] ,
    \ces_0_3_io_ins_down[38] ,
    \ces_0_3_io_ins_down[37] ,
    \ces_0_3_io_ins_down[36] ,
    \ces_0_3_io_ins_down[35] ,
    \ces_0_3_io_ins_down[34] ,
    \ces_0_3_io_ins_down[33] ,
    \ces_0_3_io_ins_down[32] ,
    \ces_0_3_io_ins_down[31] ,
    \ces_0_3_io_ins_down[30] ,
    \ces_0_3_io_ins_down[29] ,
    \ces_0_3_io_ins_down[28] ,
    \ces_0_3_io_ins_down[27] ,
    \ces_0_3_io_ins_down[26] ,
    \ces_0_3_io_ins_down[25] ,
    \ces_0_3_io_ins_down[24] ,
    \ces_0_3_io_ins_down[23] ,
    \ces_0_3_io_ins_down[22] ,
    \ces_0_3_io_ins_down[21] ,
    \ces_0_3_io_ins_down[20] ,
    \ces_0_3_io_ins_down[19] ,
    \ces_0_3_io_ins_down[18] ,
    \ces_0_3_io_ins_down[17] ,
    \ces_0_3_io_ins_down[16] ,
    \ces_0_3_io_ins_down[15] ,
    \ces_0_3_io_ins_down[14] ,
    \ces_0_3_io_ins_down[13] ,
    \ces_0_3_io_ins_down[12] ,
    \ces_0_3_io_ins_down[11] ,
    \ces_0_3_io_ins_down[10] ,
    \ces_0_3_io_ins_down[9] ,
    \ces_0_3_io_ins_down[8] ,
    \ces_0_3_io_ins_down[7] ,
    \ces_0_3_io_ins_down[6] ,
    \ces_0_3_io_ins_down[5] ,
    \ces_0_3_io_ins_down[4] ,
    \ces_0_3_io_ins_down[3] ,
    \ces_0_3_io_ins_down[2] ,
    \ces_0_3_io_ins_down[1] ,
    \ces_0_3_io_ins_down[0] }),
    .io_ins_left({\ces_0_3_io_ins_left[63] ,
    \ces_0_3_io_ins_left[62] ,
    \ces_0_3_io_ins_left[61] ,
    \ces_0_3_io_ins_left[60] ,
    \ces_0_3_io_ins_left[59] ,
    \ces_0_3_io_ins_left[58] ,
    \ces_0_3_io_ins_left[57] ,
    \ces_0_3_io_ins_left[56] ,
    \ces_0_3_io_ins_left[55] ,
    \ces_0_3_io_ins_left[54] ,
    \ces_0_3_io_ins_left[53] ,
    \ces_0_3_io_ins_left[52] ,
    \ces_0_3_io_ins_left[51] ,
    \ces_0_3_io_ins_left[50] ,
    \ces_0_3_io_ins_left[49] ,
    \ces_0_3_io_ins_left[48] ,
    \ces_0_3_io_ins_left[47] ,
    \ces_0_3_io_ins_left[46] ,
    \ces_0_3_io_ins_left[45] ,
    \ces_0_3_io_ins_left[44] ,
    \ces_0_3_io_ins_left[43] ,
    \ces_0_3_io_ins_left[42] ,
    \ces_0_3_io_ins_left[41] ,
    \ces_0_3_io_ins_left[40] ,
    \ces_0_3_io_ins_left[39] ,
    \ces_0_3_io_ins_left[38] ,
    \ces_0_3_io_ins_left[37] ,
    \ces_0_3_io_ins_left[36] ,
    \ces_0_3_io_ins_left[35] ,
    \ces_0_3_io_ins_left[34] ,
    \ces_0_3_io_ins_left[33] ,
    \ces_0_3_io_ins_left[32] ,
    \ces_0_3_io_ins_left[31] ,
    \ces_0_3_io_ins_left[30] ,
    \ces_0_3_io_ins_left[29] ,
    \ces_0_3_io_ins_left[28] ,
    \ces_0_3_io_ins_left[27] ,
    \ces_0_3_io_ins_left[26] ,
    \ces_0_3_io_ins_left[25] ,
    \ces_0_3_io_ins_left[24] ,
    \ces_0_3_io_ins_left[23] ,
    \ces_0_3_io_ins_left[22] ,
    \ces_0_3_io_ins_left[21] ,
    \ces_0_3_io_ins_left[20] ,
    \ces_0_3_io_ins_left[19] ,
    \ces_0_3_io_ins_left[18] ,
    \ces_0_3_io_ins_left[17] ,
    \ces_0_3_io_ins_left[16] ,
    \ces_0_3_io_ins_left[15] ,
    \ces_0_3_io_ins_left[14] ,
    \ces_0_3_io_ins_left[13] ,
    \ces_0_3_io_ins_left[12] ,
    \ces_0_3_io_ins_left[11] ,
    \ces_0_3_io_ins_left[10] ,
    \ces_0_3_io_ins_left[9] ,
    \ces_0_3_io_ins_left[8] ,
    \ces_0_3_io_ins_left[7] ,
    \ces_0_3_io_ins_left[6] ,
    \ces_0_3_io_ins_left[5] ,
    \ces_0_3_io_ins_left[4] ,
    \ces_0_3_io_ins_left[3] ,
    \ces_0_3_io_ins_left[2] ,
    \ces_0_3_io_ins_left[1] ,
    \ces_0_3_io_ins_left[0] }),
    .io_ins_right({\ces_0_2_io_outs_right[63] ,
    \ces_0_2_io_outs_right[62] ,
    \ces_0_2_io_outs_right[61] ,
    \ces_0_2_io_outs_right[60] ,
    \ces_0_2_io_outs_right[59] ,
    \ces_0_2_io_outs_right[58] ,
    \ces_0_2_io_outs_right[57] ,
    \ces_0_2_io_outs_right[56] ,
    \ces_0_2_io_outs_right[55] ,
    \ces_0_2_io_outs_right[54] ,
    \ces_0_2_io_outs_right[53] ,
    \ces_0_2_io_outs_right[52] ,
    \ces_0_2_io_outs_right[51] ,
    \ces_0_2_io_outs_right[50] ,
    \ces_0_2_io_outs_right[49] ,
    \ces_0_2_io_outs_right[48] ,
    \ces_0_2_io_outs_right[47] ,
    \ces_0_2_io_outs_right[46] ,
    \ces_0_2_io_outs_right[45] ,
    \ces_0_2_io_outs_right[44] ,
    \ces_0_2_io_outs_right[43] ,
    \ces_0_2_io_outs_right[42] ,
    \ces_0_2_io_outs_right[41] ,
    \ces_0_2_io_outs_right[40] ,
    \ces_0_2_io_outs_right[39] ,
    \ces_0_2_io_outs_right[38] ,
    \ces_0_2_io_outs_right[37] ,
    \ces_0_2_io_outs_right[36] ,
    \ces_0_2_io_outs_right[35] ,
    \ces_0_2_io_outs_right[34] ,
    \ces_0_2_io_outs_right[33] ,
    \ces_0_2_io_outs_right[32] ,
    \ces_0_2_io_outs_right[31] ,
    \ces_0_2_io_outs_right[30] ,
    \ces_0_2_io_outs_right[29] ,
    \ces_0_2_io_outs_right[28] ,
    \ces_0_2_io_outs_right[27] ,
    \ces_0_2_io_outs_right[26] ,
    \ces_0_2_io_outs_right[25] ,
    \ces_0_2_io_outs_right[24] ,
    \ces_0_2_io_outs_right[23] ,
    \ces_0_2_io_outs_right[22] ,
    \ces_0_2_io_outs_right[21] ,
    \ces_0_2_io_outs_right[20] ,
    \ces_0_2_io_outs_right[19] ,
    \ces_0_2_io_outs_right[18] ,
    \ces_0_2_io_outs_right[17] ,
    \ces_0_2_io_outs_right[16] ,
    \ces_0_2_io_outs_right[15] ,
    \ces_0_2_io_outs_right[14] ,
    \ces_0_2_io_outs_right[13] ,
    \ces_0_2_io_outs_right[12] ,
    \ces_0_2_io_outs_right[11] ,
    \ces_0_2_io_outs_right[10] ,
    \ces_0_2_io_outs_right[9] ,
    \ces_0_2_io_outs_right[8] ,
    \ces_0_2_io_outs_right[7] ,
    \ces_0_2_io_outs_right[6] ,
    \ces_0_2_io_outs_right[5] ,
    \ces_0_2_io_outs_right[4] ,
    \ces_0_2_io_outs_right[3] ,
    \ces_0_2_io_outs_right[2] ,
    \ces_0_2_io_outs_right[1] ,
    \ces_0_2_io_outs_right[0] }),
    .io_ins_up({net1788,
    net1787,
    net1786,
    net1785,
    net1783,
    net1782,
    net1781,
    net1780,
    net1779,
    net1778,
    net1777,
    net1776,
    net1775,
    net1774,
    net1772,
    net1771,
    net1770,
    net1769,
    net1768,
    net1767,
    net1766,
    net1765,
    net1764,
    net1763,
    net1761,
    net1760,
    net1759,
    net1758,
    net1757,
    net1756,
    net1755,
    net1754,
    net1753,
    net1752,
    net1750,
    net1749,
    net1748,
    net1747,
    net1746,
    net1745,
    net1744,
    net1743,
    net1742,
    net1741,
    net1739,
    net1738,
    net1737,
    net1736,
    net1735,
    net1734,
    net1733,
    net1732,
    net1731,
    net1730,
    net1792,
    net1791,
    net1790,
    net1789,
    net1784,
    net1773,
    net1762,
    net1751,
    net1740,
    net1729}),
    .io_outs_down({net2364,
    net2363,
    net2362,
    net2361,
    net2359,
    net2358,
    net2357,
    net2356,
    net2355,
    net2354,
    net2353,
    net2352,
    net2351,
    net2350,
    net2348,
    net2347,
    net2346,
    net2345,
    net2344,
    net2343,
    net2342,
    net2341,
    net2340,
    net2339,
    net2337,
    net2336,
    net2335,
    net2334,
    net2333,
    net2332,
    net2331,
    net2330,
    net2329,
    net2328,
    net2326,
    net2325,
    net2324,
    net2323,
    net2322,
    net2321,
    net2320,
    net2319,
    net2318,
    net2317,
    net2315,
    net2314,
    net2313,
    net2312,
    net2311,
    net2310,
    net2309,
    net2308,
    net2307,
    net2306,
    net2368,
    net2367,
    net2366,
    net2365,
    net2360,
    net2349,
    net2338,
    net2327,
    net2316,
    net2305}),
    .io_outs_left({\ces_0_2_io_ins_left[63] ,
    \ces_0_2_io_ins_left[62] ,
    \ces_0_2_io_ins_left[61] ,
    \ces_0_2_io_ins_left[60] ,
    \ces_0_2_io_ins_left[59] ,
    \ces_0_2_io_ins_left[58] ,
    \ces_0_2_io_ins_left[57] ,
    \ces_0_2_io_ins_left[56] ,
    \ces_0_2_io_ins_left[55] ,
    \ces_0_2_io_ins_left[54] ,
    \ces_0_2_io_ins_left[53] ,
    \ces_0_2_io_ins_left[52] ,
    \ces_0_2_io_ins_left[51] ,
    \ces_0_2_io_ins_left[50] ,
    \ces_0_2_io_ins_left[49] ,
    \ces_0_2_io_ins_left[48] ,
    \ces_0_2_io_ins_left[47] ,
    \ces_0_2_io_ins_left[46] ,
    \ces_0_2_io_ins_left[45] ,
    \ces_0_2_io_ins_left[44] ,
    \ces_0_2_io_ins_left[43] ,
    \ces_0_2_io_ins_left[42] ,
    \ces_0_2_io_ins_left[41] ,
    \ces_0_2_io_ins_left[40] ,
    \ces_0_2_io_ins_left[39] ,
    \ces_0_2_io_ins_left[38] ,
    \ces_0_2_io_ins_left[37] ,
    \ces_0_2_io_ins_left[36] ,
    \ces_0_2_io_ins_left[35] ,
    \ces_0_2_io_ins_left[34] ,
    \ces_0_2_io_ins_left[33] ,
    \ces_0_2_io_ins_left[32] ,
    \ces_0_2_io_ins_left[31] ,
    \ces_0_2_io_ins_left[30] ,
    \ces_0_2_io_ins_left[29] ,
    \ces_0_2_io_ins_left[28] ,
    \ces_0_2_io_ins_left[27] ,
    \ces_0_2_io_ins_left[26] ,
    \ces_0_2_io_ins_left[25] ,
    \ces_0_2_io_ins_left[24] ,
    \ces_0_2_io_ins_left[23] ,
    \ces_0_2_io_ins_left[22] ,
    \ces_0_2_io_ins_left[21] ,
    \ces_0_2_io_ins_left[20] ,
    \ces_0_2_io_ins_left[19] ,
    \ces_0_2_io_ins_left[18] ,
    \ces_0_2_io_ins_left[17] ,
    \ces_0_2_io_ins_left[16] ,
    \ces_0_2_io_ins_left[15] ,
    \ces_0_2_io_ins_left[14] ,
    \ces_0_2_io_ins_left[13] ,
    \ces_0_2_io_ins_left[12] ,
    \ces_0_2_io_ins_left[11] ,
    \ces_0_2_io_ins_left[10] ,
    \ces_0_2_io_ins_left[9] ,
    \ces_0_2_io_ins_left[8] ,
    \ces_0_2_io_ins_left[7] ,
    \ces_0_2_io_ins_left[6] ,
    \ces_0_2_io_ins_left[5] ,
    \ces_0_2_io_ins_left[4] ,
    \ces_0_2_io_ins_left[3] ,
    \ces_0_2_io_ins_left[2] ,
    \ces_0_2_io_ins_left[1] ,
    \ces_0_2_io_ins_left[0] }),
    .io_outs_right({\ces_0_3_io_outs_right[63] ,
    \ces_0_3_io_outs_right[62] ,
    \ces_0_3_io_outs_right[61] ,
    \ces_0_3_io_outs_right[60] ,
    \ces_0_3_io_outs_right[59] ,
    \ces_0_3_io_outs_right[58] ,
    \ces_0_3_io_outs_right[57] ,
    \ces_0_3_io_outs_right[56] ,
    \ces_0_3_io_outs_right[55] ,
    \ces_0_3_io_outs_right[54] ,
    \ces_0_3_io_outs_right[53] ,
    \ces_0_3_io_outs_right[52] ,
    \ces_0_3_io_outs_right[51] ,
    \ces_0_3_io_outs_right[50] ,
    \ces_0_3_io_outs_right[49] ,
    \ces_0_3_io_outs_right[48] ,
    \ces_0_3_io_outs_right[47] ,
    \ces_0_3_io_outs_right[46] ,
    \ces_0_3_io_outs_right[45] ,
    \ces_0_3_io_outs_right[44] ,
    \ces_0_3_io_outs_right[43] ,
    \ces_0_3_io_outs_right[42] ,
    \ces_0_3_io_outs_right[41] ,
    \ces_0_3_io_outs_right[40] ,
    \ces_0_3_io_outs_right[39] ,
    \ces_0_3_io_outs_right[38] ,
    \ces_0_3_io_outs_right[37] ,
    \ces_0_3_io_outs_right[36] ,
    \ces_0_3_io_outs_right[35] ,
    \ces_0_3_io_outs_right[34] ,
    \ces_0_3_io_outs_right[33] ,
    \ces_0_3_io_outs_right[32] ,
    \ces_0_3_io_outs_right[31] ,
    \ces_0_3_io_outs_right[30] ,
    \ces_0_3_io_outs_right[29] ,
    \ces_0_3_io_outs_right[28] ,
    \ces_0_3_io_outs_right[27] ,
    \ces_0_3_io_outs_right[26] ,
    \ces_0_3_io_outs_right[25] ,
    \ces_0_3_io_outs_right[24] ,
    \ces_0_3_io_outs_right[23] ,
    \ces_0_3_io_outs_right[22] ,
    \ces_0_3_io_outs_right[21] ,
    \ces_0_3_io_outs_right[20] ,
    \ces_0_3_io_outs_right[19] ,
    \ces_0_3_io_outs_right[18] ,
    \ces_0_3_io_outs_right[17] ,
    \ces_0_3_io_outs_right[16] ,
    \ces_0_3_io_outs_right[15] ,
    \ces_0_3_io_outs_right[14] ,
    \ces_0_3_io_outs_right[13] ,
    \ces_0_3_io_outs_right[12] ,
    \ces_0_3_io_outs_right[11] ,
    \ces_0_3_io_outs_right[10] ,
    \ces_0_3_io_outs_right[9] ,
    \ces_0_3_io_outs_right[8] ,
    \ces_0_3_io_outs_right[7] ,
    \ces_0_3_io_outs_right[6] ,
    \ces_0_3_io_outs_right[5] ,
    \ces_0_3_io_outs_right[4] ,
    \ces_0_3_io_outs_right[3] ,
    \ces_0_3_io_outs_right[2] ,
    \ces_0_3_io_outs_right[1] ,
    \ces_0_3_io_outs_right[0] }),
    .io_outs_up({\ces_0_3_io_outs_up[63] ,
    \ces_0_3_io_outs_up[62] ,
    \ces_0_3_io_outs_up[61] ,
    \ces_0_3_io_outs_up[60] ,
    \ces_0_3_io_outs_up[59] ,
    \ces_0_3_io_outs_up[58] ,
    \ces_0_3_io_outs_up[57] ,
    \ces_0_3_io_outs_up[56] ,
    \ces_0_3_io_outs_up[55] ,
    \ces_0_3_io_outs_up[54] ,
    \ces_0_3_io_outs_up[53] ,
    \ces_0_3_io_outs_up[52] ,
    \ces_0_3_io_outs_up[51] ,
    \ces_0_3_io_outs_up[50] ,
    \ces_0_3_io_outs_up[49] ,
    \ces_0_3_io_outs_up[48] ,
    \ces_0_3_io_outs_up[47] ,
    \ces_0_3_io_outs_up[46] ,
    \ces_0_3_io_outs_up[45] ,
    \ces_0_3_io_outs_up[44] ,
    \ces_0_3_io_outs_up[43] ,
    \ces_0_3_io_outs_up[42] ,
    \ces_0_3_io_outs_up[41] ,
    \ces_0_3_io_outs_up[40] ,
    \ces_0_3_io_outs_up[39] ,
    \ces_0_3_io_outs_up[38] ,
    \ces_0_3_io_outs_up[37] ,
    \ces_0_3_io_outs_up[36] ,
    \ces_0_3_io_outs_up[35] ,
    \ces_0_3_io_outs_up[34] ,
    \ces_0_3_io_outs_up[33] ,
    \ces_0_3_io_outs_up[32] ,
    \ces_0_3_io_outs_up[31] ,
    \ces_0_3_io_outs_up[30] ,
    \ces_0_3_io_outs_up[29] ,
    \ces_0_3_io_outs_up[28] ,
    \ces_0_3_io_outs_up[27] ,
    \ces_0_3_io_outs_up[26] ,
    \ces_0_3_io_outs_up[25] ,
    \ces_0_3_io_outs_up[24] ,
    \ces_0_3_io_outs_up[23] ,
    \ces_0_3_io_outs_up[22] ,
    \ces_0_3_io_outs_up[21] ,
    \ces_0_3_io_outs_up[20] ,
    \ces_0_3_io_outs_up[19] ,
    \ces_0_3_io_outs_up[18] ,
    \ces_0_3_io_outs_up[17] ,
    \ces_0_3_io_outs_up[16] ,
    \ces_0_3_io_outs_up[15] ,
    \ces_0_3_io_outs_up[14] ,
    \ces_0_3_io_outs_up[13] ,
    \ces_0_3_io_outs_up[12] ,
    \ces_0_3_io_outs_up[11] ,
    \ces_0_3_io_outs_up[10] ,
    \ces_0_3_io_outs_up[9] ,
    \ces_0_3_io_outs_up[8] ,
    \ces_0_3_io_outs_up[7] ,
    \ces_0_3_io_outs_up[6] ,
    \ces_0_3_io_outs_up[5] ,
    \ces_0_3_io_outs_up[4] ,
    \ces_0_3_io_outs_up[3] ,
    \ces_0_3_io_outs_up[2] ,
    \ces_0_3_io_outs_up[1] ,
    \ces_0_3_io_outs_up[0] }));
 Element ces_0_4 (.clock(clknet_3_2_0_clock),
    .io_lsbIns_1(ces_0_3_io_lsbOuts_1),
    .io_lsbIns_2(ces_0_3_io_lsbOuts_2),
    .io_lsbIns_3(ces_0_3_io_lsbOuts_3),
    .io_lsbIns_4(ces_0_3_io_lsbOuts_4),
    .io_lsbIns_5(ces_0_3_io_lsbOuts_5),
    .io_lsbIns_6(ces_0_3_io_lsbOuts_6),
    .io_lsbIns_7(ces_0_3_io_lsbOuts_7),
    .io_lsbOuts_0(ces_0_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_4_io_lsbOuts_7),
    .io_ins_down({\ces_0_4_io_ins_down[63] ,
    \ces_0_4_io_ins_down[62] ,
    \ces_0_4_io_ins_down[61] ,
    \ces_0_4_io_ins_down[60] ,
    \ces_0_4_io_ins_down[59] ,
    \ces_0_4_io_ins_down[58] ,
    \ces_0_4_io_ins_down[57] ,
    \ces_0_4_io_ins_down[56] ,
    \ces_0_4_io_ins_down[55] ,
    \ces_0_4_io_ins_down[54] ,
    \ces_0_4_io_ins_down[53] ,
    \ces_0_4_io_ins_down[52] ,
    \ces_0_4_io_ins_down[51] ,
    \ces_0_4_io_ins_down[50] ,
    \ces_0_4_io_ins_down[49] ,
    \ces_0_4_io_ins_down[48] ,
    \ces_0_4_io_ins_down[47] ,
    \ces_0_4_io_ins_down[46] ,
    \ces_0_4_io_ins_down[45] ,
    \ces_0_4_io_ins_down[44] ,
    \ces_0_4_io_ins_down[43] ,
    \ces_0_4_io_ins_down[42] ,
    \ces_0_4_io_ins_down[41] ,
    \ces_0_4_io_ins_down[40] ,
    \ces_0_4_io_ins_down[39] ,
    \ces_0_4_io_ins_down[38] ,
    \ces_0_4_io_ins_down[37] ,
    \ces_0_4_io_ins_down[36] ,
    \ces_0_4_io_ins_down[35] ,
    \ces_0_4_io_ins_down[34] ,
    \ces_0_4_io_ins_down[33] ,
    \ces_0_4_io_ins_down[32] ,
    \ces_0_4_io_ins_down[31] ,
    \ces_0_4_io_ins_down[30] ,
    \ces_0_4_io_ins_down[29] ,
    \ces_0_4_io_ins_down[28] ,
    \ces_0_4_io_ins_down[27] ,
    \ces_0_4_io_ins_down[26] ,
    \ces_0_4_io_ins_down[25] ,
    \ces_0_4_io_ins_down[24] ,
    \ces_0_4_io_ins_down[23] ,
    \ces_0_4_io_ins_down[22] ,
    \ces_0_4_io_ins_down[21] ,
    \ces_0_4_io_ins_down[20] ,
    \ces_0_4_io_ins_down[19] ,
    \ces_0_4_io_ins_down[18] ,
    \ces_0_4_io_ins_down[17] ,
    \ces_0_4_io_ins_down[16] ,
    \ces_0_4_io_ins_down[15] ,
    \ces_0_4_io_ins_down[14] ,
    \ces_0_4_io_ins_down[13] ,
    \ces_0_4_io_ins_down[12] ,
    \ces_0_4_io_ins_down[11] ,
    \ces_0_4_io_ins_down[10] ,
    \ces_0_4_io_ins_down[9] ,
    \ces_0_4_io_ins_down[8] ,
    \ces_0_4_io_ins_down[7] ,
    \ces_0_4_io_ins_down[6] ,
    \ces_0_4_io_ins_down[5] ,
    \ces_0_4_io_ins_down[4] ,
    \ces_0_4_io_ins_down[3] ,
    \ces_0_4_io_ins_down[2] ,
    \ces_0_4_io_ins_down[1] ,
    \ces_0_4_io_ins_down[0] }),
    .io_ins_left({\ces_0_4_io_ins_left[63] ,
    \ces_0_4_io_ins_left[62] ,
    \ces_0_4_io_ins_left[61] ,
    \ces_0_4_io_ins_left[60] ,
    \ces_0_4_io_ins_left[59] ,
    \ces_0_4_io_ins_left[58] ,
    \ces_0_4_io_ins_left[57] ,
    \ces_0_4_io_ins_left[56] ,
    \ces_0_4_io_ins_left[55] ,
    \ces_0_4_io_ins_left[54] ,
    \ces_0_4_io_ins_left[53] ,
    \ces_0_4_io_ins_left[52] ,
    \ces_0_4_io_ins_left[51] ,
    \ces_0_4_io_ins_left[50] ,
    \ces_0_4_io_ins_left[49] ,
    \ces_0_4_io_ins_left[48] ,
    \ces_0_4_io_ins_left[47] ,
    \ces_0_4_io_ins_left[46] ,
    \ces_0_4_io_ins_left[45] ,
    \ces_0_4_io_ins_left[44] ,
    \ces_0_4_io_ins_left[43] ,
    \ces_0_4_io_ins_left[42] ,
    \ces_0_4_io_ins_left[41] ,
    \ces_0_4_io_ins_left[40] ,
    \ces_0_4_io_ins_left[39] ,
    \ces_0_4_io_ins_left[38] ,
    \ces_0_4_io_ins_left[37] ,
    \ces_0_4_io_ins_left[36] ,
    \ces_0_4_io_ins_left[35] ,
    \ces_0_4_io_ins_left[34] ,
    \ces_0_4_io_ins_left[33] ,
    \ces_0_4_io_ins_left[32] ,
    \ces_0_4_io_ins_left[31] ,
    \ces_0_4_io_ins_left[30] ,
    \ces_0_4_io_ins_left[29] ,
    \ces_0_4_io_ins_left[28] ,
    \ces_0_4_io_ins_left[27] ,
    \ces_0_4_io_ins_left[26] ,
    \ces_0_4_io_ins_left[25] ,
    \ces_0_4_io_ins_left[24] ,
    \ces_0_4_io_ins_left[23] ,
    \ces_0_4_io_ins_left[22] ,
    \ces_0_4_io_ins_left[21] ,
    \ces_0_4_io_ins_left[20] ,
    \ces_0_4_io_ins_left[19] ,
    \ces_0_4_io_ins_left[18] ,
    \ces_0_4_io_ins_left[17] ,
    \ces_0_4_io_ins_left[16] ,
    \ces_0_4_io_ins_left[15] ,
    \ces_0_4_io_ins_left[14] ,
    \ces_0_4_io_ins_left[13] ,
    \ces_0_4_io_ins_left[12] ,
    \ces_0_4_io_ins_left[11] ,
    \ces_0_4_io_ins_left[10] ,
    \ces_0_4_io_ins_left[9] ,
    \ces_0_4_io_ins_left[8] ,
    \ces_0_4_io_ins_left[7] ,
    \ces_0_4_io_ins_left[6] ,
    \ces_0_4_io_ins_left[5] ,
    \ces_0_4_io_ins_left[4] ,
    \ces_0_4_io_ins_left[3] ,
    \ces_0_4_io_ins_left[2] ,
    \ces_0_4_io_ins_left[1] ,
    \ces_0_4_io_ins_left[0] }),
    .io_ins_right({\ces_0_3_io_outs_right[63] ,
    \ces_0_3_io_outs_right[62] ,
    \ces_0_3_io_outs_right[61] ,
    \ces_0_3_io_outs_right[60] ,
    \ces_0_3_io_outs_right[59] ,
    \ces_0_3_io_outs_right[58] ,
    \ces_0_3_io_outs_right[57] ,
    \ces_0_3_io_outs_right[56] ,
    \ces_0_3_io_outs_right[55] ,
    \ces_0_3_io_outs_right[54] ,
    \ces_0_3_io_outs_right[53] ,
    \ces_0_3_io_outs_right[52] ,
    \ces_0_3_io_outs_right[51] ,
    \ces_0_3_io_outs_right[50] ,
    \ces_0_3_io_outs_right[49] ,
    \ces_0_3_io_outs_right[48] ,
    \ces_0_3_io_outs_right[47] ,
    \ces_0_3_io_outs_right[46] ,
    \ces_0_3_io_outs_right[45] ,
    \ces_0_3_io_outs_right[44] ,
    \ces_0_3_io_outs_right[43] ,
    \ces_0_3_io_outs_right[42] ,
    \ces_0_3_io_outs_right[41] ,
    \ces_0_3_io_outs_right[40] ,
    \ces_0_3_io_outs_right[39] ,
    \ces_0_3_io_outs_right[38] ,
    \ces_0_3_io_outs_right[37] ,
    \ces_0_3_io_outs_right[36] ,
    \ces_0_3_io_outs_right[35] ,
    \ces_0_3_io_outs_right[34] ,
    \ces_0_3_io_outs_right[33] ,
    \ces_0_3_io_outs_right[32] ,
    \ces_0_3_io_outs_right[31] ,
    \ces_0_3_io_outs_right[30] ,
    \ces_0_3_io_outs_right[29] ,
    \ces_0_3_io_outs_right[28] ,
    \ces_0_3_io_outs_right[27] ,
    \ces_0_3_io_outs_right[26] ,
    \ces_0_3_io_outs_right[25] ,
    \ces_0_3_io_outs_right[24] ,
    \ces_0_3_io_outs_right[23] ,
    \ces_0_3_io_outs_right[22] ,
    \ces_0_3_io_outs_right[21] ,
    \ces_0_3_io_outs_right[20] ,
    \ces_0_3_io_outs_right[19] ,
    \ces_0_3_io_outs_right[18] ,
    \ces_0_3_io_outs_right[17] ,
    \ces_0_3_io_outs_right[16] ,
    \ces_0_3_io_outs_right[15] ,
    \ces_0_3_io_outs_right[14] ,
    \ces_0_3_io_outs_right[13] ,
    \ces_0_3_io_outs_right[12] ,
    \ces_0_3_io_outs_right[11] ,
    \ces_0_3_io_outs_right[10] ,
    \ces_0_3_io_outs_right[9] ,
    \ces_0_3_io_outs_right[8] ,
    \ces_0_3_io_outs_right[7] ,
    \ces_0_3_io_outs_right[6] ,
    \ces_0_3_io_outs_right[5] ,
    \ces_0_3_io_outs_right[4] ,
    \ces_0_3_io_outs_right[3] ,
    \ces_0_3_io_outs_right[2] ,
    \ces_0_3_io_outs_right[1] ,
    \ces_0_3_io_outs_right[0] }),
    .io_ins_up({net1852,
    net1851,
    net1850,
    net1849,
    net1847,
    net1846,
    net1845,
    net1844,
    net1843,
    net1842,
    net1841,
    net1840,
    net1839,
    net1838,
    net1836,
    net1835,
    net1834,
    net1833,
    net1832,
    net1831,
    net1830,
    net1829,
    net1828,
    net1827,
    net1825,
    net1824,
    net1823,
    net1822,
    net1821,
    net1820,
    net1819,
    net1818,
    net1817,
    net1816,
    net1814,
    net1813,
    net1812,
    net1811,
    net1810,
    net1809,
    net1808,
    net1807,
    net1806,
    net1805,
    net1803,
    net1802,
    net1801,
    net1800,
    net1799,
    net1798,
    net1797,
    net1796,
    net1795,
    net1794,
    net1856,
    net1855,
    net1854,
    net1853,
    net1848,
    net1837,
    net1826,
    net1815,
    net1804,
    net1793}),
    .io_outs_down({net2428,
    net2427,
    net2426,
    net2425,
    net2423,
    net2422,
    net2421,
    net2420,
    net2419,
    net2418,
    net2417,
    net2416,
    net2415,
    net2414,
    net2412,
    net2411,
    net2410,
    net2409,
    net2408,
    net2407,
    net2406,
    net2405,
    net2404,
    net2403,
    net2401,
    net2400,
    net2399,
    net2398,
    net2397,
    net2396,
    net2395,
    net2394,
    net2393,
    net2392,
    net2390,
    net2389,
    net2388,
    net2387,
    net2386,
    net2385,
    net2384,
    net2383,
    net2382,
    net2381,
    net2379,
    net2378,
    net2377,
    net2376,
    net2375,
    net2374,
    net2373,
    net2372,
    net2371,
    net2370,
    net2432,
    net2431,
    net2430,
    net2429,
    net2424,
    net2413,
    net2402,
    net2391,
    net2380,
    net2369}),
    .io_outs_left({\ces_0_3_io_ins_left[63] ,
    \ces_0_3_io_ins_left[62] ,
    \ces_0_3_io_ins_left[61] ,
    \ces_0_3_io_ins_left[60] ,
    \ces_0_3_io_ins_left[59] ,
    \ces_0_3_io_ins_left[58] ,
    \ces_0_3_io_ins_left[57] ,
    \ces_0_3_io_ins_left[56] ,
    \ces_0_3_io_ins_left[55] ,
    \ces_0_3_io_ins_left[54] ,
    \ces_0_3_io_ins_left[53] ,
    \ces_0_3_io_ins_left[52] ,
    \ces_0_3_io_ins_left[51] ,
    \ces_0_3_io_ins_left[50] ,
    \ces_0_3_io_ins_left[49] ,
    \ces_0_3_io_ins_left[48] ,
    \ces_0_3_io_ins_left[47] ,
    \ces_0_3_io_ins_left[46] ,
    \ces_0_3_io_ins_left[45] ,
    \ces_0_3_io_ins_left[44] ,
    \ces_0_3_io_ins_left[43] ,
    \ces_0_3_io_ins_left[42] ,
    \ces_0_3_io_ins_left[41] ,
    \ces_0_3_io_ins_left[40] ,
    \ces_0_3_io_ins_left[39] ,
    \ces_0_3_io_ins_left[38] ,
    \ces_0_3_io_ins_left[37] ,
    \ces_0_3_io_ins_left[36] ,
    \ces_0_3_io_ins_left[35] ,
    \ces_0_3_io_ins_left[34] ,
    \ces_0_3_io_ins_left[33] ,
    \ces_0_3_io_ins_left[32] ,
    \ces_0_3_io_ins_left[31] ,
    \ces_0_3_io_ins_left[30] ,
    \ces_0_3_io_ins_left[29] ,
    \ces_0_3_io_ins_left[28] ,
    \ces_0_3_io_ins_left[27] ,
    \ces_0_3_io_ins_left[26] ,
    \ces_0_3_io_ins_left[25] ,
    \ces_0_3_io_ins_left[24] ,
    \ces_0_3_io_ins_left[23] ,
    \ces_0_3_io_ins_left[22] ,
    \ces_0_3_io_ins_left[21] ,
    \ces_0_3_io_ins_left[20] ,
    \ces_0_3_io_ins_left[19] ,
    \ces_0_3_io_ins_left[18] ,
    \ces_0_3_io_ins_left[17] ,
    \ces_0_3_io_ins_left[16] ,
    \ces_0_3_io_ins_left[15] ,
    \ces_0_3_io_ins_left[14] ,
    \ces_0_3_io_ins_left[13] ,
    \ces_0_3_io_ins_left[12] ,
    \ces_0_3_io_ins_left[11] ,
    \ces_0_3_io_ins_left[10] ,
    \ces_0_3_io_ins_left[9] ,
    \ces_0_3_io_ins_left[8] ,
    \ces_0_3_io_ins_left[7] ,
    \ces_0_3_io_ins_left[6] ,
    \ces_0_3_io_ins_left[5] ,
    \ces_0_3_io_ins_left[4] ,
    \ces_0_3_io_ins_left[3] ,
    \ces_0_3_io_ins_left[2] ,
    \ces_0_3_io_ins_left[1] ,
    \ces_0_3_io_ins_left[0] }),
    .io_outs_right({\ces_0_4_io_outs_right[63] ,
    \ces_0_4_io_outs_right[62] ,
    \ces_0_4_io_outs_right[61] ,
    \ces_0_4_io_outs_right[60] ,
    \ces_0_4_io_outs_right[59] ,
    \ces_0_4_io_outs_right[58] ,
    \ces_0_4_io_outs_right[57] ,
    \ces_0_4_io_outs_right[56] ,
    \ces_0_4_io_outs_right[55] ,
    \ces_0_4_io_outs_right[54] ,
    \ces_0_4_io_outs_right[53] ,
    \ces_0_4_io_outs_right[52] ,
    \ces_0_4_io_outs_right[51] ,
    \ces_0_4_io_outs_right[50] ,
    \ces_0_4_io_outs_right[49] ,
    \ces_0_4_io_outs_right[48] ,
    \ces_0_4_io_outs_right[47] ,
    \ces_0_4_io_outs_right[46] ,
    \ces_0_4_io_outs_right[45] ,
    \ces_0_4_io_outs_right[44] ,
    \ces_0_4_io_outs_right[43] ,
    \ces_0_4_io_outs_right[42] ,
    \ces_0_4_io_outs_right[41] ,
    \ces_0_4_io_outs_right[40] ,
    \ces_0_4_io_outs_right[39] ,
    \ces_0_4_io_outs_right[38] ,
    \ces_0_4_io_outs_right[37] ,
    \ces_0_4_io_outs_right[36] ,
    \ces_0_4_io_outs_right[35] ,
    \ces_0_4_io_outs_right[34] ,
    \ces_0_4_io_outs_right[33] ,
    \ces_0_4_io_outs_right[32] ,
    \ces_0_4_io_outs_right[31] ,
    \ces_0_4_io_outs_right[30] ,
    \ces_0_4_io_outs_right[29] ,
    \ces_0_4_io_outs_right[28] ,
    \ces_0_4_io_outs_right[27] ,
    \ces_0_4_io_outs_right[26] ,
    \ces_0_4_io_outs_right[25] ,
    \ces_0_4_io_outs_right[24] ,
    \ces_0_4_io_outs_right[23] ,
    \ces_0_4_io_outs_right[22] ,
    \ces_0_4_io_outs_right[21] ,
    \ces_0_4_io_outs_right[20] ,
    \ces_0_4_io_outs_right[19] ,
    \ces_0_4_io_outs_right[18] ,
    \ces_0_4_io_outs_right[17] ,
    \ces_0_4_io_outs_right[16] ,
    \ces_0_4_io_outs_right[15] ,
    \ces_0_4_io_outs_right[14] ,
    \ces_0_4_io_outs_right[13] ,
    \ces_0_4_io_outs_right[12] ,
    \ces_0_4_io_outs_right[11] ,
    \ces_0_4_io_outs_right[10] ,
    \ces_0_4_io_outs_right[9] ,
    \ces_0_4_io_outs_right[8] ,
    \ces_0_4_io_outs_right[7] ,
    \ces_0_4_io_outs_right[6] ,
    \ces_0_4_io_outs_right[5] ,
    \ces_0_4_io_outs_right[4] ,
    \ces_0_4_io_outs_right[3] ,
    \ces_0_4_io_outs_right[2] ,
    \ces_0_4_io_outs_right[1] ,
    \ces_0_4_io_outs_right[0] }),
    .io_outs_up({\ces_0_4_io_outs_up[63] ,
    \ces_0_4_io_outs_up[62] ,
    \ces_0_4_io_outs_up[61] ,
    \ces_0_4_io_outs_up[60] ,
    \ces_0_4_io_outs_up[59] ,
    \ces_0_4_io_outs_up[58] ,
    \ces_0_4_io_outs_up[57] ,
    \ces_0_4_io_outs_up[56] ,
    \ces_0_4_io_outs_up[55] ,
    \ces_0_4_io_outs_up[54] ,
    \ces_0_4_io_outs_up[53] ,
    \ces_0_4_io_outs_up[52] ,
    \ces_0_4_io_outs_up[51] ,
    \ces_0_4_io_outs_up[50] ,
    \ces_0_4_io_outs_up[49] ,
    \ces_0_4_io_outs_up[48] ,
    \ces_0_4_io_outs_up[47] ,
    \ces_0_4_io_outs_up[46] ,
    \ces_0_4_io_outs_up[45] ,
    \ces_0_4_io_outs_up[44] ,
    \ces_0_4_io_outs_up[43] ,
    \ces_0_4_io_outs_up[42] ,
    \ces_0_4_io_outs_up[41] ,
    \ces_0_4_io_outs_up[40] ,
    \ces_0_4_io_outs_up[39] ,
    \ces_0_4_io_outs_up[38] ,
    \ces_0_4_io_outs_up[37] ,
    \ces_0_4_io_outs_up[36] ,
    \ces_0_4_io_outs_up[35] ,
    \ces_0_4_io_outs_up[34] ,
    \ces_0_4_io_outs_up[33] ,
    \ces_0_4_io_outs_up[32] ,
    \ces_0_4_io_outs_up[31] ,
    \ces_0_4_io_outs_up[30] ,
    \ces_0_4_io_outs_up[29] ,
    \ces_0_4_io_outs_up[28] ,
    \ces_0_4_io_outs_up[27] ,
    \ces_0_4_io_outs_up[26] ,
    \ces_0_4_io_outs_up[25] ,
    \ces_0_4_io_outs_up[24] ,
    \ces_0_4_io_outs_up[23] ,
    \ces_0_4_io_outs_up[22] ,
    \ces_0_4_io_outs_up[21] ,
    \ces_0_4_io_outs_up[20] ,
    \ces_0_4_io_outs_up[19] ,
    \ces_0_4_io_outs_up[18] ,
    \ces_0_4_io_outs_up[17] ,
    \ces_0_4_io_outs_up[16] ,
    \ces_0_4_io_outs_up[15] ,
    \ces_0_4_io_outs_up[14] ,
    \ces_0_4_io_outs_up[13] ,
    \ces_0_4_io_outs_up[12] ,
    \ces_0_4_io_outs_up[11] ,
    \ces_0_4_io_outs_up[10] ,
    \ces_0_4_io_outs_up[9] ,
    \ces_0_4_io_outs_up[8] ,
    \ces_0_4_io_outs_up[7] ,
    \ces_0_4_io_outs_up[6] ,
    \ces_0_4_io_outs_up[5] ,
    \ces_0_4_io_outs_up[4] ,
    \ces_0_4_io_outs_up[3] ,
    \ces_0_4_io_outs_up[2] ,
    \ces_0_4_io_outs_up[1] ,
    \ces_0_4_io_outs_up[0] }));
 Element ces_0_5 (.clock(clknet_3_2_0_clock),
    .io_lsbIns_1(ces_0_4_io_lsbOuts_1),
    .io_lsbIns_2(ces_0_4_io_lsbOuts_2),
    .io_lsbIns_3(ces_0_4_io_lsbOuts_3),
    .io_lsbIns_4(ces_0_4_io_lsbOuts_4),
    .io_lsbIns_5(ces_0_4_io_lsbOuts_5),
    .io_lsbIns_6(ces_0_4_io_lsbOuts_6),
    .io_lsbIns_7(ces_0_4_io_lsbOuts_7),
    .io_lsbOuts_0(ces_0_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_5_io_lsbOuts_7),
    .io_ins_down({\ces_0_5_io_ins_down[63] ,
    \ces_0_5_io_ins_down[62] ,
    \ces_0_5_io_ins_down[61] ,
    \ces_0_5_io_ins_down[60] ,
    \ces_0_5_io_ins_down[59] ,
    \ces_0_5_io_ins_down[58] ,
    \ces_0_5_io_ins_down[57] ,
    \ces_0_5_io_ins_down[56] ,
    \ces_0_5_io_ins_down[55] ,
    \ces_0_5_io_ins_down[54] ,
    \ces_0_5_io_ins_down[53] ,
    \ces_0_5_io_ins_down[52] ,
    \ces_0_5_io_ins_down[51] ,
    \ces_0_5_io_ins_down[50] ,
    \ces_0_5_io_ins_down[49] ,
    \ces_0_5_io_ins_down[48] ,
    \ces_0_5_io_ins_down[47] ,
    \ces_0_5_io_ins_down[46] ,
    \ces_0_5_io_ins_down[45] ,
    \ces_0_5_io_ins_down[44] ,
    \ces_0_5_io_ins_down[43] ,
    \ces_0_5_io_ins_down[42] ,
    \ces_0_5_io_ins_down[41] ,
    \ces_0_5_io_ins_down[40] ,
    \ces_0_5_io_ins_down[39] ,
    \ces_0_5_io_ins_down[38] ,
    \ces_0_5_io_ins_down[37] ,
    \ces_0_5_io_ins_down[36] ,
    \ces_0_5_io_ins_down[35] ,
    \ces_0_5_io_ins_down[34] ,
    \ces_0_5_io_ins_down[33] ,
    \ces_0_5_io_ins_down[32] ,
    \ces_0_5_io_ins_down[31] ,
    \ces_0_5_io_ins_down[30] ,
    \ces_0_5_io_ins_down[29] ,
    \ces_0_5_io_ins_down[28] ,
    \ces_0_5_io_ins_down[27] ,
    \ces_0_5_io_ins_down[26] ,
    \ces_0_5_io_ins_down[25] ,
    \ces_0_5_io_ins_down[24] ,
    \ces_0_5_io_ins_down[23] ,
    \ces_0_5_io_ins_down[22] ,
    \ces_0_5_io_ins_down[21] ,
    \ces_0_5_io_ins_down[20] ,
    \ces_0_5_io_ins_down[19] ,
    \ces_0_5_io_ins_down[18] ,
    \ces_0_5_io_ins_down[17] ,
    \ces_0_5_io_ins_down[16] ,
    \ces_0_5_io_ins_down[15] ,
    \ces_0_5_io_ins_down[14] ,
    \ces_0_5_io_ins_down[13] ,
    \ces_0_5_io_ins_down[12] ,
    \ces_0_5_io_ins_down[11] ,
    \ces_0_5_io_ins_down[10] ,
    \ces_0_5_io_ins_down[9] ,
    \ces_0_5_io_ins_down[8] ,
    \ces_0_5_io_ins_down[7] ,
    \ces_0_5_io_ins_down[6] ,
    \ces_0_5_io_ins_down[5] ,
    \ces_0_5_io_ins_down[4] ,
    \ces_0_5_io_ins_down[3] ,
    \ces_0_5_io_ins_down[2] ,
    \ces_0_5_io_ins_down[1] ,
    \ces_0_5_io_ins_down[0] }),
    .io_ins_left({\ces_0_5_io_ins_left[63] ,
    \ces_0_5_io_ins_left[62] ,
    \ces_0_5_io_ins_left[61] ,
    \ces_0_5_io_ins_left[60] ,
    \ces_0_5_io_ins_left[59] ,
    \ces_0_5_io_ins_left[58] ,
    \ces_0_5_io_ins_left[57] ,
    \ces_0_5_io_ins_left[56] ,
    \ces_0_5_io_ins_left[55] ,
    \ces_0_5_io_ins_left[54] ,
    \ces_0_5_io_ins_left[53] ,
    \ces_0_5_io_ins_left[52] ,
    \ces_0_5_io_ins_left[51] ,
    \ces_0_5_io_ins_left[50] ,
    \ces_0_5_io_ins_left[49] ,
    \ces_0_5_io_ins_left[48] ,
    \ces_0_5_io_ins_left[47] ,
    \ces_0_5_io_ins_left[46] ,
    \ces_0_5_io_ins_left[45] ,
    \ces_0_5_io_ins_left[44] ,
    \ces_0_5_io_ins_left[43] ,
    \ces_0_5_io_ins_left[42] ,
    \ces_0_5_io_ins_left[41] ,
    \ces_0_5_io_ins_left[40] ,
    \ces_0_5_io_ins_left[39] ,
    \ces_0_5_io_ins_left[38] ,
    \ces_0_5_io_ins_left[37] ,
    \ces_0_5_io_ins_left[36] ,
    \ces_0_5_io_ins_left[35] ,
    \ces_0_5_io_ins_left[34] ,
    \ces_0_5_io_ins_left[33] ,
    \ces_0_5_io_ins_left[32] ,
    \ces_0_5_io_ins_left[31] ,
    \ces_0_5_io_ins_left[30] ,
    \ces_0_5_io_ins_left[29] ,
    \ces_0_5_io_ins_left[28] ,
    \ces_0_5_io_ins_left[27] ,
    \ces_0_5_io_ins_left[26] ,
    \ces_0_5_io_ins_left[25] ,
    \ces_0_5_io_ins_left[24] ,
    \ces_0_5_io_ins_left[23] ,
    \ces_0_5_io_ins_left[22] ,
    \ces_0_5_io_ins_left[21] ,
    \ces_0_5_io_ins_left[20] ,
    \ces_0_5_io_ins_left[19] ,
    \ces_0_5_io_ins_left[18] ,
    \ces_0_5_io_ins_left[17] ,
    \ces_0_5_io_ins_left[16] ,
    \ces_0_5_io_ins_left[15] ,
    \ces_0_5_io_ins_left[14] ,
    \ces_0_5_io_ins_left[13] ,
    \ces_0_5_io_ins_left[12] ,
    \ces_0_5_io_ins_left[11] ,
    \ces_0_5_io_ins_left[10] ,
    \ces_0_5_io_ins_left[9] ,
    \ces_0_5_io_ins_left[8] ,
    \ces_0_5_io_ins_left[7] ,
    \ces_0_5_io_ins_left[6] ,
    \ces_0_5_io_ins_left[5] ,
    \ces_0_5_io_ins_left[4] ,
    \ces_0_5_io_ins_left[3] ,
    \ces_0_5_io_ins_left[2] ,
    \ces_0_5_io_ins_left[1] ,
    \ces_0_5_io_ins_left[0] }),
    .io_ins_right({\ces_0_4_io_outs_right[63] ,
    \ces_0_4_io_outs_right[62] ,
    \ces_0_4_io_outs_right[61] ,
    \ces_0_4_io_outs_right[60] ,
    \ces_0_4_io_outs_right[59] ,
    \ces_0_4_io_outs_right[58] ,
    \ces_0_4_io_outs_right[57] ,
    \ces_0_4_io_outs_right[56] ,
    \ces_0_4_io_outs_right[55] ,
    \ces_0_4_io_outs_right[54] ,
    \ces_0_4_io_outs_right[53] ,
    \ces_0_4_io_outs_right[52] ,
    \ces_0_4_io_outs_right[51] ,
    \ces_0_4_io_outs_right[50] ,
    \ces_0_4_io_outs_right[49] ,
    \ces_0_4_io_outs_right[48] ,
    \ces_0_4_io_outs_right[47] ,
    \ces_0_4_io_outs_right[46] ,
    \ces_0_4_io_outs_right[45] ,
    \ces_0_4_io_outs_right[44] ,
    \ces_0_4_io_outs_right[43] ,
    \ces_0_4_io_outs_right[42] ,
    \ces_0_4_io_outs_right[41] ,
    \ces_0_4_io_outs_right[40] ,
    \ces_0_4_io_outs_right[39] ,
    \ces_0_4_io_outs_right[38] ,
    \ces_0_4_io_outs_right[37] ,
    \ces_0_4_io_outs_right[36] ,
    \ces_0_4_io_outs_right[35] ,
    \ces_0_4_io_outs_right[34] ,
    \ces_0_4_io_outs_right[33] ,
    \ces_0_4_io_outs_right[32] ,
    \ces_0_4_io_outs_right[31] ,
    \ces_0_4_io_outs_right[30] ,
    \ces_0_4_io_outs_right[29] ,
    \ces_0_4_io_outs_right[28] ,
    \ces_0_4_io_outs_right[27] ,
    \ces_0_4_io_outs_right[26] ,
    \ces_0_4_io_outs_right[25] ,
    \ces_0_4_io_outs_right[24] ,
    \ces_0_4_io_outs_right[23] ,
    \ces_0_4_io_outs_right[22] ,
    \ces_0_4_io_outs_right[21] ,
    \ces_0_4_io_outs_right[20] ,
    \ces_0_4_io_outs_right[19] ,
    \ces_0_4_io_outs_right[18] ,
    \ces_0_4_io_outs_right[17] ,
    \ces_0_4_io_outs_right[16] ,
    \ces_0_4_io_outs_right[15] ,
    \ces_0_4_io_outs_right[14] ,
    \ces_0_4_io_outs_right[13] ,
    \ces_0_4_io_outs_right[12] ,
    \ces_0_4_io_outs_right[11] ,
    \ces_0_4_io_outs_right[10] ,
    \ces_0_4_io_outs_right[9] ,
    \ces_0_4_io_outs_right[8] ,
    \ces_0_4_io_outs_right[7] ,
    \ces_0_4_io_outs_right[6] ,
    \ces_0_4_io_outs_right[5] ,
    \ces_0_4_io_outs_right[4] ,
    \ces_0_4_io_outs_right[3] ,
    \ces_0_4_io_outs_right[2] ,
    \ces_0_4_io_outs_right[1] ,
    \ces_0_4_io_outs_right[0] }),
    .io_ins_up({net1916,
    net1915,
    net1914,
    net1913,
    net1911,
    net1910,
    net1909,
    net1908,
    net1907,
    net1906,
    net1905,
    net1904,
    net1903,
    net1902,
    net1900,
    net1899,
    net1898,
    net1897,
    net1896,
    net1895,
    net1894,
    net1893,
    net1892,
    net1891,
    net1889,
    net1888,
    net1887,
    net1886,
    net1885,
    net1884,
    net1883,
    net1882,
    net1881,
    net1880,
    net1878,
    net1877,
    net1876,
    net1875,
    net1874,
    net1873,
    net1872,
    net1871,
    net1870,
    net1869,
    net1867,
    net1866,
    net1865,
    net1864,
    net1863,
    net1862,
    net1861,
    net1860,
    net1859,
    net1858,
    net1920,
    net1919,
    net1918,
    net1917,
    net1912,
    net1901,
    net1890,
    net1879,
    net1868,
    net1857}),
    .io_outs_down({net2492,
    net2491,
    net2490,
    net2489,
    net2487,
    net2486,
    net2485,
    net2484,
    net2483,
    net2482,
    net2481,
    net2480,
    net2479,
    net2478,
    net2476,
    net2475,
    net2474,
    net2473,
    net2472,
    net2471,
    net2470,
    net2469,
    net2468,
    net2467,
    net2465,
    net2464,
    net2463,
    net2462,
    net2461,
    net2460,
    net2459,
    net2458,
    net2457,
    net2456,
    net2454,
    net2453,
    net2452,
    net2451,
    net2450,
    net2449,
    net2448,
    net2447,
    net2446,
    net2445,
    net2443,
    net2442,
    net2441,
    net2440,
    net2439,
    net2438,
    net2437,
    net2436,
    net2435,
    net2434,
    net2496,
    net2495,
    net2494,
    net2493,
    net2488,
    net2477,
    net2466,
    net2455,
    net2444,
    net2433}),
    .io_outs_left({\ces_0_4_io_ins_left[63] ,
    \ces_0_4_io_ins_left[62] ,
    \ces_0_4_io_ins_left[61] ,
    \ces_0_4_io_ins_left[60] ,
    \ces_0_4_io_ins_left[59] ,
    \ces_0_4_io_ins_left[58] ,
    \ces_0_4_io_ins_left[57] ,
    \ces_0_4_io_ins_left[56] ,
    \ces_0_4_io_ins_left[55] ,
    \ces_0_4_io_ins_left[54] ,
    \ces_0_4_io_ins_left[53] ,
    \ces_0_4_io_ins_left[52] ,
    \ces_0_4_io_ins_left[51] ,
    \ces_0_4_io_ins_left[50] ,
    \ces_0_4_io_ins_left[49] ,
    \ces_0_4_io_ins_left[48] ,
    \ces_0_4_io_ins_left[47] ,
    \ces_0_4_io_ins_left[46] ,
    \ces_0_4_io_ins_left[45] ,
    \ces_0_4_io_ins_left[44] ,
    \ces_0_4_io_ins_left[43] ,
    \ces_0_4_io_ins_left[42] ,
    \ces_0_4_io_ins_left[41] ,
    \ces_0_4_io_ins_left[40] ,
    \ces_0_4_io_ins_left[39] ,
    \ces_0_4_io_ins_left[38] ,
    \ces_0_4_io_ins_left[37] ,
    \ces_0_4_io_ins_left[36] ,
    \ces_0_4_io_ins_left[35] ,
    \ces_0_4_io_ins_left[34] ,
    \ces_0_4_io_ins_left[33] ,
    \ces_0_4_io_ins_left[32] ,
    \ces_0_4_io_ins_left[31] ,
    \ces_0_4_io_ins_left[30] ,
    \ces_0_4_io_ins_left[29] ,
    \ces_0_4_io_ins_left[28] ,
    \ces_0_4_io_ins_left[27] ,
    \ces_0_4_io_ins_left[26] ,
    \ces_0_4_io_ins_left[25] ,
    \ces_0_4_io_ins_left[24] ,
    \ces_0_4_io_ins_left[23] ,
    \ces_0_4_io_ins_left[22] ,
    \ces_0_4_io_ins_left[21] ,
    \ces_0_4_io_ins_left[20] ,
    \ces_0_4_io_ins_left[19] ,
    \ces_0_4_io_ins_left[18] ,
    \ces_0_4_io_ins_left[17] ,
    \ces_0_4_io_ins_left[16] ,
    \ces_0_4_io_ins_left[15] ,
    \ces_0_4_io_ins_left[14] ,
    \ces_0_4_io_ins_left[13] ,
    \ces_0_4_io_ins_left[12] ,
    \ces_0_4_io_ins_left[11] ,
    \ces_0_4_io_ins_left[10] ,
    \ces_0_4_io_ins_left[9] ,
    \ces_0_4_io_ins_left[8] ,
    \ces_0_4_io_ins_left[7] ,
    \ces_0_4_io_ins_left[6] ,
    \ces_0_4_io_ins_left[5] ,
    \ces_0_4_io_ins_left[4] ,
    \ces_0_4_io_ins_left[3] ,
    \ces_0_4_io_ins_left[2] ,
    \ces_0_4_io_ins_left[1] ,
    \ces_0_4_io_ins_left[0] }),
    .io_outs_right({\ces_0_5_io_outs_right[63] ,
    \ces_0_5_io_outs_right[62] ,
    \ces_0_5_io_outs_right[61] ,
    \ces_0_5_io_outs_right[60] ,
    \ces_0_5_io_outs_right[59] ,
    \ces_0_5_io_outs_right[58] ,
    \ces_0_5_io_outs_right[57] ,
    \ces_0_5_io_outs_right[56] ,
    \ces_0_5_io_outs_right[55] ,
    \ces_0_5_io_outs_right[54] ,
    \ces_0_5_io_outs_right[53] ,
    \ces_0_5_io_outs_right[52] ,
    \ces_0_5_io_outs_right[51] ,
    \ces_0_5_io_outs_right[50] ,
    \ces_0_5_io_outs_right[49] ,
    \ces_0_5_io_outs_right[48] ,
    \ces_0_5_io_outs_right[47] ,
    \ces_0_5_io_outs_right[46] ,
    \ces_0_5_io_outs_right[45] ,
    \ces_0_5_io_outs_right[44] ,
    \ces_0_5_io_outs_right[43] ,
    \ces_0_5_io_outs_right[42] ,
    \ces_0_5_io_outs_right[41] ,
    \ces_0_5_io_outs_right[40] ,
    \ces_0_5_io_outs_right[39] ,
    \ces_0_5_io_outs_right[38] ,
    \ces_0_5_io_outs_right[37] ,
    \ces_0_5_io_outs_right[36] ,
    \ces_0_5_io_outs_right[35] ,
    \ces_0_5_io_outs_right[34] ,
    \ces_0_5_io_outs_right[33] ,
    \ces_0_5_io_outs_right[32] ,
    \ces_0_5_io_outs_right[31] ,
    \ces_0_5_io_outs_right[30] ,
    \ces_0_5_io_outs_right[29] ,
    \ces_0_5_io_outs_right[28] ,
    \ces_0_5_io_outs_right[27] ,
    \ces_0_5_io_outs_right[26] ,
    \ces_0_5_io_outs_right[25] ,
    \ces_0_5_io_outs_right[24] ,
    \ces_0_5_io_outs_right[23] ,
    \ces_0_5_io_outs_right[22] ,
    \ces_0_5_io_outs_right[21] ,
    \ces_0_5_io_outs_right[20] ,
    \ces_0_5_io_outs_right[19] ,
    \ces_0_5_io_outs_right[18] ,
    \ces_0_5_io_outs_right[17] ,
    \ces_0_5_io_outs_right[16] ,
    \ces_0_5_io_outs_right[15] ,
    \ces_0_5_io_outs_right[14] ,
    \ces_0_5_io_outs_right[13] ,
    \ces_0_5_io_outs_right[12] ,
    \ces_0_5_io_outs_right[11] ,
    \ces_0_5_io_outs_right[10] ,
    \ces_0_5_io_outs_right[9] ,
    \ces_0_5_io_outs_right[8] ,
    \ces_0_5_io_outs_right[7] ,
    \ces_0_5_io_outs_right[6] ,
    \ces_0_5_io_outs_right[5] ,
    \ces_0_5_io_outs_right[4] ,
    \ces_0_5_io_outs_right[3] ,
    \ces_0_5_io_outs_right[2] ,
    \ces_0_5_io_outs_right[1] ,
    \ces_0_5_io_outs_right[0] }),
    .io_outs_up({\ces_0_5_io_outs_up[63] ,
    \ces_0_5_io_outs_up[62] ,
    \ces_0_5_io_outs_up[61] ,
    \ces_0_5_io_outs_up[60] ,
    \ces_0_5_io_outs_up[59] ,
    \ces_0_5_io_outs_up[58] ,
    \ces_0_5_io_outs_up[57] ,
    \ces_0_5_io_outs_up[56] ,
    \ces_0_5_io_outs_up[55] ,
    \ces_0_5_io_outs_up[54] ,
    \ces_0_5_io_outs_up[53] ,
    \ces_0_5_io_outs_up[52] ,
    \ces_0_5_io_outs_up[51] ,
    \ces_0_5_io_outs_up[50] ,
    \ces_0_5_io_outs_up[49] ,
    \ces_0_5_io_outs_up[48] ,
    \ces_0_5_io_outs_up[47] ,
    \ces_0_5_io_outs_up[46] ,
    \ces_0_5_io_outs_up[45] ,
    \ces_0_5_io_outs_up[44] ,
    \ces_0_5_io_outs_up[43] ,
    \ces_0_5_io_outs_up[42] ,
    \ces_0_5_io_outs_up[41] ,
    \ces_0_5_io_outs_up[40] ,
    \ces_0_5_io_outs_up[39] ,
    \ces_0_5_io_outs_up[38] ,
    \ces_0_5_io_outs_up[37] ,
    \ces_0_5_io_outs_up[36] ,
    \ces_0_5_io_outs_up[35] ,
    \ces_0_5_io_outs_up[34] ,
    \ces_0_5_io_outs_up[33] ,
    \ces_0_5_io_outs_up[32] ,
    \ces_0_5_io_outs_up[31] ,
    \ces_0_5_io_outs_up[30] ,
    \ces_0_5_io_outs_up[29] ,
    \ces_0_5_io_outs_up[28] ,
    \ces_0_5_io_outs_up[27] ,
    \ces_0_5_io_outs_up[26] ,
    \ces_0_5_io_outs_up[25] ,
    \ces_0_5_io_outs_up[24] ,
    \ces_0_5_io_outs_up[23] ,
    \ces_0_5_io_outs_up[22] ,
    \ces_0_5_io_outs_up[21] ,
    \ces_0_5_io_outs_up[20] ,
    \ces_0_5_io_outs_up[19] ,
    \ces_0_5_io_outs_up[18] ,
    \ces_0_5_io_outs_up[17] ,
    \ces_0_5_io_outs_up[16] ,
    \ces_0_5_io_outs_up[15] ,
    \ces_0_5_io_outs_up[14] ,
    \ces_0_5_io_outs_up[13] ,
    \ces_0_5_io_outs_up[12] ,
    \ces_0_5_io_outs_up[11] ,
    \ces_0_5_io_outs_up[10] ,
    \ces_0_5_io_outs_up[9] ,
    \ces_0_5_io_outs_up[8] ,
    \ces_0_5_io_outs_up[7] ,
    \ces_0_5_io_outs_up[6] ,
    \ces_0_5_io_outs_up[5] ,
    \ces_0_5_io_outs_up[4] ,
    \ces_0_5_io_outs_up[3] ,
    \ces_0_5_io_outs_up[2] ,
    \ces_0_5_io_outs_up[1] ,
    \ces_0_5_io_outs_up[0] }));
 Element ces_0_6 (.clock(clknet_3_2_0_clock),
    .io_lsbIns_1(ces_0_5_io_lsbOuts_1),
    .io_lsbIns_2(ces_0_5_io_lsbOuts_2),
    .io_lsbIns_3(ces_0_5_io_lsbOuts_3),
    .io_lsbIns_4(ces_0_5_io_lsbOuts_4),
    .io_lsbIns_5(ces_0_5_io_lsbOuts_5),
    .io_lsbIns_6(ces_0_5_io_lsbOuts_6),
    .io_lsbIns_7(ces_0_5_io_lsbOuts_7),
    .io_lsbOuts_0(ces_0_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_6_io_lsbOuts_7),
    .io_ins_down({\ces_0_6_io_ins_down[63] ,
    \ces_0_6_io_ins_down[62] ,
    \ces_0_6_io_ins_down[61] ,
    \ces_0_6_io_ins_down[60] ,
    \ces_0_6_io_ins_down[59] ,
    \ces_0_6_io_ins_down[58] ,
    \ces_0_6_io_ins_down[57] ,
    \ces_0_6_io_ins_down[56] ,
    \ces_0_6_io_ins_down[55] ,
    \ces_0_6_io_ins_down[54] ,
    \ces_0_6_io_ins_down[53] ,
    \ces_0_6_io_ins_down[52] ,
    \ces_0_6_io_ins_down[51] ,
    \ces_0_6_io_ins_down[50] ,
    \ces_0_6_io_ins_down[49] ,
    \ces_0_6_io_ins_down[48] ,
    \ces_0_6_io_ins_down[47] ,
    \ces_0_6_io_ins_down[46] ,
    \ces_0_6_io_ins_down[45] ,
    \ces_0_6_io_ins_down[44] ,
    \ces_0_6_io_ins_down[43] ,
    \ces_0_6_io_ins_down[42] ,
    \ces_0_6_io_ins_down[41] ,
    \ces_0_6_io_ins_down[40] ,
    \ces_0_6_io_ins_down[39] ,
    \ces_0_6_io_ins_down[38] ,
    \ces_0_6_io_ins_down[37] ,
    \ces_0_6_io_ins_down[36] ,
    \ces_0_6_io_ins_down[35] ,
    \ces_0_6_io_ins_down[34] ,
    \ces_0_6_io_ins_down[33] ,
    \ces_0_6_io_ins_down[32] ,
    \ces_0_6_io_ins_down[31] ,
    \ces_0_6_io_ins_down[30] ,
    \ces_0_6_io_ins_down[29] ,
    \ces_0_6_io_ins_down[28] ,
    \ces_0_6_io_ins_down[27] ,
    \ces_0_6_io_ins_down[26] ,
    \ces_0_6_io_ins_down[25] ,
    \ces_0_6_io_ins_down[24] ,
    \ces_0_6_io_ins_down[23] ,
    \ces_0_6_io_ins_down[22] ,
    \ces_0_6_io_ins_down[21] ,
    \ces_0_6_io_ins_down[20] ,
    \ces_0_6_io_ins_down[19] ,
    \ces_0_6_io_ins_down[18] ,
    \ces_0_6_io_ins_down[17] ,
    \ces_0_6_io_ins_down[16] ,
    \ces_0_6_io_ins_down[15] ,
    \ces_0_6_io_ins_down[14] ,
    \ces_0_6_io_ins_down[13] ,
    \ces_0_6_io_ins_down[12] ,
    \ces_0_6_io_ins_down[11] ,
    \ces_0_6_io_ins_down[10] ,
    \ces_0_6_io_ins_down[9] ,
    \ces_0_6_io_ins_down[8] ,
    \ces_0_6_io_ins_down[7] ,
    \ces_0_6_io_ins_down[6] ,
    \ces_0_6_io_ins_down[5] ,
    \ces_0_6_io_ins_down[4] ,
    \ces_0_6_io_ins_down[3] ,
    \ces_0_6_io_ins_down[2] ,
    \ces_0_6_io_ins_down[1] ,
    \ces_0_6_io_ins_down[0] }),
    .io_ins_left({\ces_0_6_io_ins_left[63] ,
    \ces_0_6_io_ins_left[62] ,
    \ces_0_6_io_ins_left[61] ,
    \ces_0_6_io_ins_left[60] ,
    \ces_0_6_io_ins_left[59] ,
    \ces_0_6_io_ins_left[58] ,
    \ces_0_6_io_ins_left[57] ,
    \ces_0_6_io_ins_left[56] ,
    \ces_0_6_io_ins_left[55] ,
    \ces_0_6_io_ins_left[54] ,
    \ces_0_6_io_ins_left[53] ,
    \ces_0_6_io_ins_left[52] ,
    \ces_0_6_io_ins_left[51] ,
    \ces_0_6_io_ins_left[50] ,
    \ces_0_6_io_ins_left[49] ,
    \ces_0_6_io_ins_left[48] ,
    \ces_0_6_io_ins_left[47] ,
    \ces_0_6_io_ins_left[46] ,
    \ces_0_6_io_ins_left[45] ,
    \ces_0_6_io_ins_left[44] ,
    \ces_0_6_io_ins_left[43] ,
    \ces_0_6_io_ins_left[42] ,
    \ces_0_6_io_ins_left[41] ,
    \ces_0_6_io_ins_left[40] ,
    \ces_0_6_io_ins_left[39] ,
    \ces_0_6_io_ins_left[38] ,
    \ces_0_6_io_ins_left[37] ,
    \ces_0_6_io_ins_left[36] ,
    \ces_0_6_io_ins_left[35] ,
    \ces_0_6_io_ins_left[34] ,
    \ces_0_6_io_ins_left[33] ,
    \ces_0_6_io_ins_left[32] ,
    \ces_0_6_io_ins_left[31] ,
    \ces_0_6_io_ins_left[30] ,
    \ces_0_6_io_ins_left[29] ,
    \ces_0_6_io_ins_left[28] ,
    \ces_0_6_io_ins_left[27] ,
    \ces_0_6_io_ins_left[26] ,
    \ces_0_6_io_ins_left[25] ,
    \ces_0_6_io_ins_left[24] ,
    \ces_0_6_io_ins_left[23] ,
    \ces_0_6_io_ins_left[22] ,
    \ces_0_6_io_ins_left[21] ,
    \ces_0_6_io_ins_left[20] ,
    \ces_0_6_io_ins_left[19] ,
    \ces_0_6_io_ins_left[18] ,
    \ces_0_6_io_ins_left[17] ,
    \ces_0_6_io_ins_left[16] ,
    \ces_0_6_io_ins_left[15] ,
    \ces_0_6_io_ins_left[14] ,
    \ces_0_6_io_ins_left[13] ,
    \ces_0_6_io_ins_left[12] ,
    \ces_0_6_io_ins_left[11] ,
    \ces_0_6_io_ins_left[10] ,
    \ces_0_6_io_ins_left[9] ,
    \ces_0_6_io_ins_left[8] ,
    \ces_0_6_io_ins_left[7] ,
    \ces_0_6_io_ins_left[6] ,
    \ces_0_6_io_ins_left[5] ,
    \ces_0_6_io_ins_left[4] ,
    \ces_0_6_io_ins_left[3] ,
    \ces_0_6_io_ins_left[2] ,
    \ces_0_6_io_ins_left[1] ,
    \ces_0_6_io_ins_left[0] }),
    .io_ins_right({\ces_0_5_io_outs_right[63] ,
    \ces_0_5_io_outs_right[62] ,
    \ces_0_5_io_outs_right[61] ,
    \ces_0_5_io_outs_right[60] ,
    \ces_0_5_io_outs_right[59] ,
    \ces_0_5_io_outs_right[58] ,
    \ces_0_5_io_outs_right[57] ,
    \ces_0_5_io_outs_right[56] ,
    \ces_0_5_io_outs_right[55] ,
    \ces_0_5_io_outs_right[54] ,
    \ces_0_5_io_outs_right[53] ,
    \ces_0_5_io_outs_right[52] ,
    \ces_0_5_io_outs_right[51] ,
    \ces_0_5_io_outs_right[50] ,
    \ces_0_5_io_outs_right[49] ,
    \ces_0_5_io_outs_right[48] ,
    \ces_0_5_io_outs_right[47] ,
    \ces_0_5_io_outs_right[46] ,
    \ces_0_5_io_outs_right[45] ,
    \ces_0_5_io_outs_right[44] ,
    \ces_0_5_io_outs_right[43] ,
    \ces_0_5_io_outs_right[42] ,
    \ces_0_5_io_outs_right[41] ,
    \ces_0_5_io_outs_right[40] ,
    \ces_0_5_io_outs_right[39] ,
    \ces_0_5_io_outs_right[38] ,
    \ces_0_5_io_outs_right[37] ,
    \ces_0_5_io_outs_right[36] ,
    \ces_0_5_io_outs_right[35] ,
    \ces_0_5_io_outs_right[34] ,
    \ces_0_5_io_outs_right[33] ,
    \ces_0_5_io_outs_right[32] ,
    \ces_0_5_io_outs_right[31] ,
    \ces_0_5_io_outs_right[30] ,
    \ces_0_5_io_outs_right[29] ,
    \ces_0_5_io_outs_right[28] ,
    \ces_0_5_io_outs_right[27] ,
    \ces_0_5_io_outs_right[26] ,
    \ces_0_5_io_outs_right[25] ,
    \ces_0_5_io_outs_right[24] ,
    \ces_0_5_io_outs_right[23] ,
    \ces_0_5_io_outs_right[22] ,
    \ces_0_5_io_outs_right[21] ,
    \ces_0_5_io_outs_right[20] ,
    \ces_0_5_io_outs_right[19] ,
    \ces_0_5_io_outs_right[18] ,
    \ces_0_5_io_outs_right[17] ,
    \ces_0_5_io_outs_right[16] ,
    \ces_0_5_io_outs_right[15] ,
    \ces_0_5_io_outs_right[14] ,
    \ces_0_5_io_outs_right[13] ,
    \ces_0_5_io_outs_right[12] ,
    \ces_0_5_io_outs_right[11] ,
    \ces_0_5_io_outs_right[10] ,
    \ces_0_5_io_outs_right[9] ,
    \ces_0_5_io_outs_right[8] ,
    \ces_0_5_io_outs_right[7] ,
    \ces_0_5_io_outs_right[6] ,
    \ces_0_5_io_outs_right[5] ,
    \ces_0_5_io_outs_right[4] ,
    \ces_0_5_io_outs_right[3] ,
    \ces_0_5_io_outs_right[2] ,
    \ces_0_5_io_outs_right[1] ,
    \ces_0_5_io_outs_right[0] }),
    .io_ins_up({net1980,
    net1979,
    net1978,
    net1977,
    net1975,
    net1974,
    net1973,
    net1972,
    net1971,
    net1970,
    net1969,
    net1968,
    net1967,
    net1966,
    net1964,
    net1963,
    net1962,
    net1961,
    net1960,
    net1959,
    net1958,
    net1957,
    net1956,
    net1955,
    net1953,
    net1952,
    net1951,
    net1950,
    net1949,
    net1948,
    net1947,
    net1946,
    net1945,
    net1944,
    net1942,
    net1941,
    net1940,
    net1939,
    net1938,
    net1937,
    net1936,
    net1935,
    net1934,
    net1933,
    net1931,
    net1930,
    net1929,
    net1928,
    net1927,
    net1926,
    net1925,
    net1924,
    net1923,
    net1922,
    net1984,
    net1983,
    net1982,
    net1981,
    net1976,
    net1965,
    net1954,
    net1943,
    net1932,
    net1921}),
    .io_outs_down({net2556,
    net2555,
    net2554,
    net2553,
    net2551,
    net2550,
    net2549,
    net2548,
    net2547,
    net2546,
    net2545,
    net2544,
    net2543,
    net2542,
    net2540,
    net2539,
    net2538,
    net2537,
    net2536,
    net2535,
    net2534,
    net2533,
    net2532,
    net2531,
    net2529,
    net2528,
    net2527,
    net2526,
    net2525,
    net2524,
    net2523,
    net2522,
    net2521,
    net2520,
    net2518,
    net2517,
    net2516,
    net2515,
    net2514,
    net2513,
    net2512,
    net2511,
    net2510,
    net2509,
    net2507,
    net2506,
    net2505,
    net2504,
    net2503,
    net2502,
    net2501,
    net2500,
    net2499,
    net2498,
    net2560,
    net2559,
    net2558,
    net2557,
    net2552,
    net2541,
    net2530,
    net2519,
    net2508,
    net2497}),
    .io_outs_left({\ces_0_5_io_ins_left[63] ,
    \ces_0_5_io_ins_left[62] ,
    \ces_0_5_io_ins_left[61] ,
    \ces_0_5_io_ins_left[60] ,
    \ces_0_5_io_ins_left[59] ,
    \ces_0_5_io_ins_left[58] ,
    \ces_0_5_io_ins_left[57] ,
    \ces_0_5_io_ins_left[56] ,
    \ces_0_5_io_ins_left[55] ,
    \ces_0_5_io_ins_left[54] ,
    \ces_0_5_io_ins_left[53] ,
    \ces_0_5_io_ins_left[52] ,
    \ces_0_5_io_ins_left[51] ,
    \ces_0_5_io_ins_left[50] ,
    \ces_0_5_io_ins_left[49] ,
    \ces_0_5_io_ins_left[48] ,
    \ces_0_5_io_ins_left[47] ,
    \ces_0_5_io_ins_left[46] ,
    \ces_0_5_io_ins_left[45] ,
    \ces_0_5_io_ins_left[44] ,
    \ces_0_5_io_ins_left[43] ,
    \ces_0_5_io_ins_left[42] ,
    \ces_0_5_io_ins_left[41] ,
    \ces_0_5_io_ins_left[40] ,
    \ces_0_5_io_ins_left[39] ,
    \ces_0_5_io_ins_left[38] ,
    \ces_0_5_io_ins_left[37] ,
    \ces_0_5_io_ins_left[36] ,
    \ces_0_5_io_ins_left[35] ,
    \ces_0_5_io_ins_left[34] ,
    \ces_0_5_io_ins_left[33] ,
    \ces_0_5_io_ins_left[32] ,
    \ces_0_5_io_ins_left[31] ,
    \ces_0_5_io_ins_left[30] ,
    \ces_0_5_io_ins_left[29] ,
    \ces_0_5_io_ins_left[28] ,
    \ces_0_5_io_ins_left[27] ,
    \ces_0_5_io_ins_left[26] ,
    \ces_0_5_io_ins_left[25] ,
    \ces_0_5_io_ins_left[24] ,
    \ces_0_5_io_ins_left[23] ,
    \ces_0_5_io_ins_left[22] ,
    \ces_0_5_io_ins_left[21] ,
    \ces_0_5_io_ins_left[20] ,
    \ces_0_5_io_ins_left[19] ,
    \ces_0_5_io_ins_left[18] ,
    \ces_0_5_io_ins_left[17] ,
    \ces_0_5_io_ins_left[16] ,
    \ces_0_5_io_ins_left[15] ,
    \ces_0_5_io_ins_left[14] ,
    \ces_0_5_io_ins_left[13] ,
    \ces_0_5_io_ins_left[12] ,
    \ces_0_5_io_ins_left[11] ,
    \ces_0_5_io_ins_left[10] ,
    \ces_0_5_io_ins_left[9] ,
    \ces_0_5_io_ins_left[8] ,
    \ces_0_5_io_ins_left[7] ,
    \ces_0_5_io_ins_left[6] ,
    \ces_0_5_io_ins_left[5] ,
    \ces_0_5_io_ins_left[4] ,
    \ces_0_5_io_ins_left[3] ,
    \ces_0_5_io_ins_left[2] ,
    \ces_0_5_io_ins_left[1] ,
    \ces_0_5_io_ins_left[0] }),
    .io_outs_right({\ces_0_6_io_outs_right[63] ,
    \ces_0_6_io_outs_right[62] ,
    \ces_0_6_io_outs_right[61] ,
    \ces_0_6_io_outs_right[60] ,
    \ces_0_6_io_outs_right[59] ,
    \ces_0_6_io_outs_right[58] ,
    \ces_0_6_io_outs_right[57] ,
    \ces_0_6_io_outs_right[56] ,
    \ces_0_6_io_outs_right[55] ,
    \ces_0_6_io_outs_right[54] ,
    \ces_0_6_io_outs_right[53] ,
    \ces_0_6_io_outs_right[52] ,
    \ces_0_6_io_outs_right[51] ,
    \ces_0_6_io_outs_right[50] ,
    \ces_0_6_io_outs_right[49] ,
    \ces_0_6_io_outs_right[48] ,
    \ces_0_6_io_outs_right[47] ,
    \ces_0_6_io_outs_right[46] ,
    \ces_0_6_io_outs_right[45] ,
    \ces_0_6_io_outs_right[44] ,
    \ces_0_6_io_outs_right[43] ,
    \ces_0_6_io_outs_right[42] ,
    \ces_0_6_io_outs_right[41] ,
    \ces_0_6_io_outs_right[40] ,
    \ces_0_6_io_outs_right[39] ,
    \ces_0_6_io_outs_right[38] ,
    \ces_0_6_io_outs_right[37] ,
    \ces_0_6_io_outs_right[36] ,
    \ces_0_6_io_outs_right[35] ,
    \ces_0_6_io_outs_right[34] ,
    \ces_0_6_io_outs_right[33] ,
    \ces_0_6_io_outs_right[32] ,
    \ces_0_6_io_outs_right[31] ,
    \ces_0_6_io_outs_right[30] ,
    \ces_0_6_io_outs_right[29] ,
    \ces_0_6_io_outs_right[28] ,
    \ces_0_6_io_outs_right[27] ,
    \ces_0_6_io_outs_right[26] ,
    \ces_0_6_io_outs_right[25] ,
    \ces_0_6_io_outs_right[24] ,
    \ces_0_6_io_outs_right[23] ,
    \ces_0_6_io_outs_right[22] ,
    \ces_0_6_io_outs_right[21] ,
    \ces_0_6_io_outs_right[20] ,
    \ces_0_6_io_outs_right[19] ,
    \ces_0_6_io_outs_right[18] ,
    \ces_0_6_io_outs_right[17] ,
    \ces_0_6_io_outs_right[16] ,
    \ces_0_6_io_outs_right[15] ,
    \ces_0_6_io_outs_right[14] ,
    \ces_0_6_io_outs_right[13] ,
    \ces_0_6_io_outs_right[12] ,
    \ces_0_6_io_outs_right[11] ,
    \ces_0_6_io_outs_right[10] ,
    \ces_0_6_io_outs_right[9] ,
    \ces_0_6_io_outs_right[8] ,
    \ces_0_6_io_outs_right[7] ,
    \ces_0_6_io_outs_right[6] ,
    \ces_0_6_io_outs_right[5] ,
    \ces_0_6_io_outs_right[4] ,
    \ces_0_6_io_outs_right[3] ,
    \ces_0_6_io_outs_right[2] ,
    \ces_0_6_io_outs_right[1] ,
    \ces_0_6_io_outs_right[0] }),
    .io_outs_up({\ces_0_6_io_outs_up[63] ,
    \ces_0_6_io_outs_up[62] ,
    \ces_0_6_io_outs_up[61] ,
    \ces_0_6_io_outs_up[60] ,
    \ces_0_6_io_outs_up[59] ,
    \ces_0_6_io_outs_up[58] ,
    \ces_0_6_io_outs_up[57] ,
    \ces_0_6_io_outs_up[56] ,
    \ces_0_6_io_outs_up[55] ,
    \ces_0_6_io_outs_up[54] ,
    \ces_0_6_io_outs_up[53] ,
    \ces_0_6_io_outs_up[52] ,
    \ces_0_6_io_outs_up[51] ,
    \ces_0_6_io_outs_up[50] ,
    \ces_0_6_io_outs_up[49] ,
    \ces_0_6_io_outs_up[48] ,
    \ces_0_6_io_outs_up[47] ,
    \ces_0_6_io_outs_up[46] ,
    \ces_0_6_io_outs_up[45] ,
    \ces_0_6_io_outs_up[44] ,
    \ces_0_6_io_outs_up[43] ,
    \ces_0_6_io_outs_up[42] ,
    \ces_0_6_io_outs_up[41] ,
    \ces_0_6_io_outs_up[40] ,
    \ces_0_6_io_outs_up[39] ,
    \ces_0_6_io_outs_up[38] ,
    \ces_0_6_io_outs_up[37] ,
    \ces_0_6_io_outs_up[36] ,
    \ces_0_6_io_outs_up[35] ,
    \ces_0_6_io_outs_up[34] ,
    \ces_0_6_io_outs_up[33] ,
    \ces_0_6_io_outs_up[32] ,
    \ces_0_6_io_outs_up[31] ,
    \ces_0_6_io_outs_up[30] ,
    \ces_0_6_io_outs_up[29] ,
    \ces_0_6_io_outs_up[28] ,
    \ces_0_6_io_outs_up[27] ,
    \ces_0_6_io_outs_up[26] ,
    \ces_0_6_io_outs_up[25] ,
    \ces_0_6_io_outs_up[24] ,
    \ces_0_6_io_outs_up[23] ,
    \ces_0_6_io_outs_up[22] ,
    \ces_0_6_io_outs_up[21] ,
    \ces_0_6_io_outs_up[20] ,
    \ces_0_6_io_outs_up[19] ,
    \ces_0_6_io_outs_up[18] ,
    \ces_0_6_io_outs_up[17] ,
    \ces_0_6_io_outs_up[16] ,
    \ces_0_6_io_outs_up[15] ,
    \ces_0_6_io_outs_up[14] ,
    \ces_0_6_io_outs_up[13] ,
    \ces_0_6_io_outs_up[12] ,
    \ces_0_6_io_outs_up[11] ,
    \ces_0_6_io_outs_up[10] ,
    \ces_0_6_io_outs_up[9] ,
    \ces_0_6_io_outs_up[8] ,
    \ces_0_6_io_outs_up[7] ,
    \ces_0_6_io_outs_up[6] ,
    \ces_0_6_io_outs_up[5] ,
    \ces_0_6_io_outs_up[4] ,
    \ces_0_6_io_outs_up[3] ,
    \ces_0_6_io_outs_up[2] ,
    \ces_0_6_io_outs_up[1] ,
    \ces_0_6_io_outs_up[0] }));
 Element ces_0_7 (.clock(clknet_3_2_0_clock),
    .io_lsbIns_1(ces_0_6_io_lsbOuts_1),
    .io_lsbIns_2(ces_0_6_io_lsbOuts_2),
    .io_lsbIns_3(ces_0_6_io_lsbOuts_3),
    .io_lsbIns_4(ces_0_6_io_lsbOuts_4),
    .io_lsbIns_5(ces_0_6_io_lsbOuts_5),
    .io_lsbIns_6(ces_0_6_io_lsbOuts_6),
    .io_lsbIns_7(ces_0_6_io_lsbOuts_7),
    .io_lsbOuts_0(ces_0_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_0_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_0_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_0_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_0_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_0_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_0_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_0_7_io_lsbOuts_7),
    .io_ins_down({\ces_0_7_io_ins_down[63] ,
    \ces_0_7_io_ins_down[62] ,
    \ces_0_7_io_ins_down[61] ,
    \ces_0_7_io_ins_down[60] ,
    \ces_0_7_io_ins_down[59] ,
    \ces_0_7_io_ins_down[58] ,
    \ces_0_7_io_ins_down[57] ,
    \ces_0_7_io_ins_down[56] ,
    \ces_0_7_io_ins_down[55] ,
    \ces_0_7_io_ins_down[54] ,
    \ces_0_7_io_ins_down[53] ,
    \ces_0_7_io_ins_down[52] ,
    \ces_0_7_io_ins_down[51] ,
    \ces_0_7_io_ins_down[50] ,
    \ces_0_7_io_ins_down[49] ,
    \ces_0_7_io_ins_down[48] ,
    \ces_0_7_io_ins_down[47] ,
    \ces_0_7_io_ins_down[46] ,
    \ces_0_7_io_ins_down[45] ,
    \ces_0_7_io_ins_down[44] ,
    \ces_0_7_io_ins_down[43] ,
    \ces_0_7_io_ins_down[42] ,
    \ces_0_7_io_ins_down[41] ,
    \ces_0_7_io_ins_down[40] ,
    \ces_0_7_io_ins_down[39] ,
    \ces_0_7_io_ins_down[38] ,
    \ces_0_7_io_ins_down[37] ,
    \ces_0_7_io_ins_down[36] ,
    \ces_0_7_io_ins_down[35] ,
    \ces_0_7_io_ins_down[34] ,
    \ces_0_7_io_ins_down[33] ,
    \ces_0_7_io_ins_down[32] ,
    \ces_0_7_io_ins_down[31] ,
    \ces_0_7_io_ins_down[30] ,
    \ces_0_7_io_ins_down[29] ,
    \ces_0_7_io_ins_down[28] ,
    \ces_0_7_io_ins_down[27] ,
    \ces_0_7_io_ins_down[26] ,
    \ces_0_7_io_ins_down[25] ,
    \ces_0_7_io_ins_down[24] ,
    \ces_0_7_io_ins_down[23] ,
    \ces_0_7_io_ins_down[22] ,
    \ces_0_7_io_ins_down[21] ,
    \ces_0_7_io_ins_down[20] ,
    \ces_0_7_io_ins_down[19] ,
    \ces_0_7_io_ins_down[18] ,
    \ces_0_7_io_ins_down[17] ,
    \ces_0_7_io_ins_down[16] ,
    \ces_0_7_io_ins_down[15] ,
    \ces_0_7_io_ins_down[14] ,
    \ces_0_7_io_ins_down[13] ,
    \ces_0_7_io_ins_down[12] ,
    \ces_0_7_io_ins_down[11] ,
    \ces_0_7_io_ins_down[10] ,
    \ces_0_7_io_ins_down[9] ,
    \ces_0_7_io_ins_down[8] ,
    \ces_0_7_io_ins_down[7] ,
    \ces_0_7_io_ins_down[6] ,
    \ces_0_7_io_ins_down[5] ,
    \ces_0_7_io_ins_down[4] ,
    \ces_0_7_io_ins_down[3] ,
    \ces_0_7_io_ins_down[2] ,
    \ces_0_7_io_ins_down[1] ,
    \ces_0_7_io_ins_down[0] }),
    .io_ins_left({net572,
    net571,
    net570,
    net569,
    net567,
    net566,
    net565,
    net564,
    net563,
    net562,
    net561,
    net560,
    net559,
    net558,
    net556,
    net555,
    net554,
    net553,
    net552,
    net551,
    net550,
    net549,
    net548,
    net547,
    net545,
    net544,
    net543,
    net542,
    net541,
    net540,
    net539,
    net538,
    net537,
    net536,
    net534,
    net533,
    net532,
    net531,
    net530,
    net529,
    net528,
    net527,
    net526,
    net525,
    net523,
    net522,
    net521,
    net520,
    net519,
    net518,
    net517,
    net516,
    net515,
    net514,
    net576,
    net575,
    net574,
    net573,
    net568,
    net557,
    net546,
    net535,
    net524,
    net513}),
    .io_ins_right({\ces_0_6_io_outs_right[63] ,
    \ces_0_6_io_outs_right[62] ,
    \ces_0_6_io_outs_right[61] ,
    \ces_0_6_io_outs_right[60] ,
    \ces_0_6_io_outs_right[59] ,
    \ces_0_6_io_outs_right[58] ,
    \ces_0_6_io_outs_right[57] ,
    \ces_0_6_io_outs_right[56] ,
    \ces_0_6_io_outs_right[55] ,
    \ces_0_6_io_outs_right[54] ,
    \ces_0_6_io_outs_right[53] ,
    \ces_0_6_io_outs_right[52] ,
    \ces_0_6_io_outs_right[51] ,
    \ces_0_6_io_outs_right[50] ,
    \ces_0_6_io_outs_right[49] ,
    \ces_0_6_io_outs_right[48] ,
    \ces_0_6_io_outs_right[47] ,
    \ces_0_6_io_outs_right[46] ,
    \ces_0_6_io_outs_right[45] ,
    \ces_0_6_io_outs_right[44] ,
    \ces_0_6_io_outs_right[43] ,
    \ces_0_6_io_outs_right[42] ,
    \ces_0_6_io_outs_right[41] ,
    \ces_0_6_io_outs_right[40] ,
    \ces_0_6_io_outs_right[39] ,
    \ces_0_6_io_outs_right[38] ,
    \ces_0_6_io_outs_right[37] ,
    \ces_0_6_io_outs_right[36] ,
    \ces_0_6_io_outs_right[35] ,
    \ces_0_6_io_outs_right[34] ,
    \ces_0_6_io_outs_right[33] ,
    \ces_0_6_io_outs_right[32] ,
    \ces_0_6_io_outs_right[31] ,
    \ces_0_6_io_outs_right[30] ,
    \ces_0_6_io_outs_right[29] ,
    \ces_0_6_io_outs_right[28] ,
    \ces_0_6_io_outs_right[27] ,
    \ces_0_6_io_outs_right[26] ,
    \ces_0_6_io_outs_right[25] ,
    \ces_0_6_io_outs_right[24] ,
    \ces_0_6_io_outs_right[23] ,
    \ces_0_6_io_outs_right[22] ,
    \ces_0_6_io_outs_right[21] ,
    \ces_0_6_io_outs_right[20] ,
    \ces_0_6_io_outs_right[19] ,
    \ces_0_6_io_outs_right[18] ,
    \ces_0_6_io_outs_right[17] ,
    \ces_0_6_io_outs_right[16] ,
    \ces_0_6_io_outs_right[15] ,
    \ces_0_6_io_outs_right[14] ,
    \ces_0_6_io_outs_right[13] ,
    \ces_0_6_io_outs_right[12] ,
    \ces_0_6_io_outs_right[11] ,
    \ces_0_6_io_outs_right[10] ,
    \ces_0_6_io_outs_right[9] ,
    \ces_0_6_io_outs_right[8] ,
    \ces_0_6_io_outs_right[7] ,
    \ces_0_6_io_outs_right[6] ,
    \ces_0_6_io_outs_right[5] ,
    \ces_0_6_io_outs_right[4] ,
    \ces_0_6_io_outs_right[3] ,
    \ces_0_6_io_outs_right[2] ,
    \ces_0_6_io_outs_right[1] ,
    \ces_0_6_io_outs_right[0] }),
    .io_ins_up({net2044,
    net2043,
    net2042,
    net2041,
    net2039,
    net2038,
    net2037,
    net2036,
    net2035,
    net2034,
    net2033,
    net2032,
    net2031,
    net2030,
    net2028,
    net2027,
    net2026,
    net2025,
    net2024,
    net2023,
    net2022,
    net2021,
    net2020,
    net2019,
    net2017,
    net2016,
    net2015,
    net2014,
    net2013,
    net2012,
    net2011,
    net2010,
    net2009,
    net2008,
    net2006,
    net2005,
    net2004,
    net2003,
    net2002,
    net2001,
    net2000,
    net1999,
    net1998,
    net1997,
    net1995,
    net1994,
    net1993,
    net1992,
    net1991,
    net1990,
    net1989,
    net1988,
    net1987,
    net1986,
    net2048,
    net2047,
    net2046,
    net2045,
    net2040,
    net2029,
    net2018,
    net2007,
    net1996,
    net1985}),
    .io_outs_down({net2620,
    net2619,
    net2618,
    net2617,
    net2615,
    net2614,
    net2613,
    net2612,
    net2611,
    net2610,
    net2609,
    net2608,
    net2607,
    net2606,
    net2604,
    net2603,
    net2602,
    net2601,
    net2600,
    net2599,
    net2598,
    net2597,
    net2596,
    net2595,
    net2593,
    net2592,
    net2591,
    net2590,
    net2589,
    net2588,
    net2587,
    net2586,
    net2585,
    net2584,
    net2582,
    net2581,
    net2580,
    net2579,
    net2578,
    net2577,
    net2576,
    net2575,
    net2574,
    net2573,
    net2571,
    net2570,
    net2569,
    net2568,
    net2567,
    net2566,
    net2565,
    net2564,
    net2563,
    net2562,
    net2624,
    net2623,
    net2622,
    net2621,
    net2616,
    net2605,
    net2594,
    net2583,
    net2572,
    net2561}),
    .io_outs_left({\ces_0_6_io_ins_left[63] ,
    \ces_0_6_io_ins_left[62] ,
    \ces_0_6_io_ins_left[61] ,
    \ces_0_6_io_ins_left[60] ,
    \ces_0_6_io_ins_left[59] ,
    \ces_0_6_io_ins_left[58] ,
    \ces_0_6_io_ins_left[57] ,
    \ces_0_6_io_ins_left[56] ,
    \ces_0_6_io_ins_left[55] ,
    \ces_0_6_io_ins_left[54] ,
    \ces_0_6_io_ins_left[53] ,
    \ces_0_6_io_ins_left[52] ,
    \ces_0_6_io_ins_left[51] ,
    \ces_0_6_io_ins_left[50] ,
    \ces_0_6_io_ins_left[49] ,
    \ces_0_6_io_ins_left[48] ,
    \ces_0_6_io_ins_left[47] ,
    \ces_0_6_io_ins_left[46] ,
    \ces_0_6_io_ins_left[45] ,
    \ces_0_6_io_ins_left[44] ,
    \ces_0_6_io_ins_left[43] ,
    \ces_0_6_io_ins_left[42] ,
    \ces_0_6_io_ins_left[41] ,
    \ces_0_6_io_ins_left[40] ,
    \ces_0_6_io_ins_left[39] ,
    \ces_0_6_io_ins_left[38] ,
    \ces_0_6_io_ins_left[37] ,
    \ces_0_6_io_ins_left[36] ,
    \ces_0_6_io_ins_left[35] ,
    \ces_0_6_io_ins_left[34] ,
    \ces_0_6_io_ins_left[33] ,
    \ces_0_6_io_ins_left[32] ,
    \ces_0_6_io_ins_left[31] ,
    \ces_0_6_io_ins_left[30] ,
    \ces_0_6_io_ins_left[29] ,
    \ces_0_6_io_ins_left[28] ,
    \ces_0_6_io_ins_left[27] ,
    \ces_0_6_io_ins_left[26] ,
    \ces_0_6_io_ins_left[25] ,
    \ces_0_6_io_ins_left[24] ,
    \ces_0_6_io_ins_left[23] ,
    \ces_0_6_io_ins_left[22] ,
    \ces_0_6_io_ins_left[21] ,
    \ces_0_6_io_ins_left[20] ,
    \ces_0_6_io_ins_left[19] ,
    \ces_0_6_io_ins_left[18] ,
    \ces_0_6_io_ins_left[17] ,
    \ces_0_6_io_ins_left[16] ,
    \ces_0_6_io_ins_left[15] ,
    \ces_0_6_io_ins_left[14] ,
    \ces_0_6_io_ins_left[13] ,
    \ces_0_6_io_ins_left[12] ,
    \ces_0_6_io_ins_left[11] ,
    \ces_0_6_io_ins_left[10] ,
    \ces_0_6_io_ins_left[9] ,
    \ces_0_6_io_ins_left[8] ,
    \ces_0_6_io_ins_left[7] ,
    \ces_0_6_io_ins_left[6] ,
    \ces_0_6_io_ins_left[5] ,
    \ces_0_6_io_ins_left[4] ,
    \ces_0_6_io_ins_left[3] ,
    \ces_0_6_io_ins_left[2] ,
    \ces_0_6_io_ins_left[1] ,
    \ces_0_6_io_ins_left[0] }),
    .io_outs_right({net3196,
    net3195,
    net3194,
    net3193,
    net3191,
    net3190,
    net3189,
    net3188,
    net3187,
    net3186,
    net3185,
    net3184,
    net3183,
    net3182,
    net3180,
    net3179,
    net3178,
    net3177,
    net3176,
    net3175,
    net3174,
    net3173,
    net3172,
    net3171,
    net3169,
    net3168,
    net3167,
    net3166,
    net3165,
    net3164,
    net3163,
    net3162,
    net3161,
    net3160,
    net3158,
    net3157,
    net3156,
    net3155,
    net3154,
    net3153,
    net3152,
    net3151,
    net3150,
    net3149,
    net3147,
    net3146,
    net3145,
    net3144,
    net3143,
    net3142,
    net3141,
    net3140,
    net3139,
    net3138,
    net3200,
    net3199,
    net3198,
    net3197,
    net3192,
    net3181,
    net3170,
    net3159,
    net3148,
    net3137}),
    .io_outs_up({\ces_0_7_io_outs_up[63] ,
    \ces_0_7_io_outs_up[62] ,
    \ces_0_7_io_outs_up[61] ,
    \ces_0_7_io_outs_up[60] ,
    \ces_0_7_io_outs_up[59] ,
    \ces_0_7_io_outs_up[58] ,
    \ces_0_7_io_outs_up[57] ,
    \ces_0_7_io_outs_up[56] ,
    \ces_0_7_io_outs_up[55] ,
    \ces_0_7_io_outs_up[54] ,
    \ces_0_7_io_outs_up[53] ,
    \ces_0_7_io_outs_up[52] ,
    \ces_0_7_io_outs_up[51] ,
    \ces_0_7_io_outs_up[50] ,
    \ces_0_7_io_outs_up[49] ,
    \ces_0_7_io_outs_up[48] ,
    \ces_0_7_io_outs_up[47] ,
    \ces_0_7_io_outs_up[46] ,
    \ces_0_7_io_outs_up[45] ,
    \ces_0_7_io_outs_up[44] ,
    \ces_0_7_io_outs_up[43] ,
    \ces_0_7_io_outs_up[42] ,
    \ces_0_7_io_outs_up[41] ,
    \ces_0_7_io_outs_up[40] ,
    \ces_0_7_io_outs_up[39] ,
    \ces_0_7_io_outs_up[38] ,
    \ces_0_7_io_outs_up[37] ,
    \ces_0_7_io_outs_up[36] ,
    \ces_0_7_io_outs_up[35] ,
    \ces_0_7_io_outs_up[34] ,
    \ces_0_7_io_outs_up[33] ,
    \ces_0_7_io_outs_up[32] ,
    \ces_0_7_io_outs_up[31] ,
    \ces_0_7_io_outs_up[30] ,
    \ces_0_7_io_outs_up[29] ,
    \ces_0_7_io_outs_up[28] ,
    \ces_0_7_io_outs_up[27] ,
    \ces_0_7_io_outs_up[26] ,
    \ces_0_7_io_outs_up[25] ,
    \ces_0_7_io_outs_up[24] ,
    \ces_0_7_io_outs_up[23] ,
    \ces_0_7_io_outs_up[22] ,
    \ces_0_7_io_outs_up[21] ,
    \ces_0_7_io_outs_up[20] ,
    \ces_0_7_io_outs_up[19] ,
    \ces_0_7_io_outs_up[18] ,
    \ces_0_7_io_outs_up[17] ,
    \ces_0_7_io_outs_up[16] ,
    \ces_0_7_io_outs_up[15] ,
    \ces_0_7_io_outs_up[14] ,
    \ces_0_7_io_outs_up[13] ,
    \ces_0_7_io_outs_up[12] ,
    \ces_0_7_io_outs_up[11] ,
    \ces_0_7_io_outs_up[10] ,
    \ces_0_7_io_outs_up[9] ,
    \ces_0_7_io_outs_up[8] ,
    \ces_0_7_io_outs_up[7] ,
    \ces_0_7_io_outs_up[6] ,
    \ces_0_7_io_outs_up[5] ,
    \ces_0_7_io_outs_up[4] ,
    \ces_0_7_io_outs_up[3] ,
    \ces_0_7_io_outs_up[2] ,
    \ces_0_7_io_outs_up[1] ,
    \ces_0_7_io_outs_up[0] }));
 Element ces_1_0 (.clock(clknet_3_0_0_clock),
    .io_lsbIns_1(net4168),
    .io_lsbIns_2(net4169),
    .io_lsbIns_3(net4170),
    .io_lsbIns_4(net4171),
    .io_lsbIns_5(net4172),
    .io_lsbIns_6(net4173),
    .io_lsbIns_7(net4174),
    .io_lsbOuts_0(ces_1_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_0_io_lsbOuts_7),
    .io_ins_down({\ces_1_0_io_ins_down[63] ,
    \ces_1_0_io_ins_down[62] ,
    \ces_1_0_io_ins_down[61] ,
    \ces_1_0_io_ins_down[60] ,
    \ces_1_0_io_ins_down[59] ,
    \ces_1_0_io_ins_down[58] ,
    \ces_1_0_io_ins_down[57] ,
    \ces_1_0_io_ins_down[56] ,
    \ces_1_0_io_ins_down[55] ,
    \ces_1_0_io_ins_down[54] ,
    \ces_1_0_io_ins_down[53] ,
    \ces_1_0_io_ins_down[52] ,
    \ces_1_0_io_ins_down[51] ,
    \ces_1_0_io_ins_down[50] ,
    \ces_1_0_io_ins_down[49] ,
    \ces_1_0_io_ins_down[48] ,
    \ces_1_0_io_ins_down[47] ,
    \ces_1_0_io_ins_down[46] ,
    \ces_1_0_io_ins_down[45] ,
    \ces_1_0_io_ins_down[44] ,
    \ces_1_0_io_ins_down[43] ,
    \ces_1_0_io_ins_down[42] ,
    \ces_1_0_io_ins_down[41] ,
    \ces_1_0_io_ins_down[40] ,
    \ces_1_0_io_ins_down[39] ,
    \ces_1_0_io_ins_down[38] ,
    \ces_1_0_io_ins_down[37] ,
    \ces_1_0_io_ins_down[36] ,
    \ces_1_0_io_ins_down[35] ,
    \ces_1_0_io_ins_down[34] ,
    \ces_1_0_io_ins_down[33] ,
    \ces_1_0_io_ins_down[32] ,
    \ces_1_0_io_ins_down[31] ,
    \ces_1_0_io_ins_down[30] ,
    \ces_1_0_io_ins_down[29] ,
    \ces_1_0_io_ins_down[28] ,
    \ces_1_0_io_ins_down[27] ,
    \ces_1_0_io_ins_down[26] ,
    \ces_1_0_io_ins_down[25] ,
    \ces_1_0_io_ins_down[24] ,
    \ces_1_0_io_ins_down[23] ,
    \ces_1_0_io_ins_down[22] ,
    \ces_1_0_io_ins_down[21] ,
    \ces_1_0_io_ins_down[20] ,
    \ces_1_0_io_ins_down[19] ,
    \ces_1_0_io_ins_down[18] ,
    \ces_1_0_io_ins_down[17] ,
    \ces_1_0_io_ins_down[16] ,
    \ces_1_0_io_ins_down[15] ,
    \ces_1_0_io_ins_down[14] ,
    \ces_1_0_io_ins_down[13] ,
    \ces_1_0_io_ins_down[12] ,
    \ces_1_0_io_ins_down[11] ,
    \ces_1_0_io_ins_down[10] ,
    \ces_1_0_io_ins_down[9] ,
    \ces_1_0_io_ins_down[8] ,
    \ces_1_0_io_ins_down[7] ,
    \ces_1_0_io_ins_down[6] ,
    \ces_1_0_io_ins_down[5] ,
    \ces_1_0_io_ins_down[4] ,
    \ces_1_0_io_ins_down[3] ,
    \ces_1_0_io_ins_down[2] ,
    \ces_1_0_io_ins_down[1] ,
    \ces_1_0_io_ins_down[0] }),
    .io_ins_left({\ces_1_0_io_ins_left[63] ,
    \ces_1_0_io_ins_left[62] ,
    \ces_1_0_io_ins_left[61] ,
    \ces_1_0_io_ins_left[60] ,
    \ces_1_0_io_ins_left[59] ,
    \ces_1_0_io_ins_left[58] ,
    \ces_1_0_io_ins_left[57] ,
    \ces_1_0_io_ins_left[56] ,
    \ces_1_0_io_ins_left[55] ,
    \ces_1_0_io_ins_left[54] ,
    \ces_1_0_io_ins_left[53] ,
    \ces_1_0_io_ins_left[52] ,
    \ces_1_0_io_ins_left[51] ,
    \ces_1_0_io_ins_left[50] ,
    \ces_1_0_io_ins_left[49] ,
    \ces_1_0_io_ins_left[48] ,
    \ces_1_0_io_ins_left[47] ,
    \ces_1_0_io_ins_left[46] ,
    \ces_1_0_io_ins_left[45] ,
    \ces_1_0_io_ins_left[44] ,
    \ces_1_0_io_ins_left[43] ,
    \ces_1_0_io_ins_left[42] ,
    \ces_1_0_io_ins_left[41] ,
    \ces_1_0_io_ins_left[40] ,
    \ces_1_0_io_ins_left[39] ,
    \ces_1_0_io_ins_left[38] ,
    \ces_1_0_io_ins_left[37] ,
    \ces_1_0_io_ins_left[36] ,
    \ces_1_0_io_ins_left[35] ,
    \ces_1_0_io_ins_left[34] ,
    \ces_1_0_io_ins_left[33] ,
    \ces_1_0_io_ins_left[32] ,
    \ces_1_0_io_ins_left[31] ,
    \ces_1_0_io_ins_left[30] ,
    \ces_1_0_io_ins_left[29] ,
    \ces_1_0_io_ins_left[28] ,
    \ces_1_0_io_ins_left[27] ,
    \ces_1_0_io_ins_left[26] ,
    \ces_1_0_io_ins_left[25] ,
    \ces_1_0_io_ins_left[24] ,
    \ces_1_0_io_ins_left[23] ,
    \ces_1_0_io_ins_left[22] ,
    \ces_1_0_io_ins_left[21] ,
    \ces_1_0_io_ins_left[20] ,
    \ces_1_0_io_ins_left[19] ,
    \ces_1_0_io_ins_left[18] ,
    \ces_1_0_io_ins_left[17] ,
    \ces_1_0_io_ins_left[16] ,
    \ces_1_0_io_ins_left[15] ,
    \ces_1_0_io_ins_left[14] ,
    \ces_1_0_io_ins_left[13] ,
    \ces_1_0_io_ins_left[12] ,
    \ces_1_0_io_ins_left[11] ,
    \ces_1_0_io_ins_left[10] ,
    \ces_1_0_io_ins_left[9] ,
    \ces_1_0_io_ins_left[8] ,
    \ces_1_0_io_ins_left[7] ,
    \ces_1_0_io_ins_left[6] ,
    \ces_1_0_io_ins_left[5] ,
    \ces_1_0_io_ins_left[4] ,
    \ces_1_0_io_ins_left[3] ,
    \ces_1_0_io_ins_left[2] ,
    \ces_1_0_io_ins_left[1] ,
    \ces_1_0_io_ins_left[0] }),
    .io_ins_right({net1148,
    net1147,
    net1146,
    net1145,
    net1143,
    net1142,
    net1141,
    net1140,
    net1139,
    net1138,
    net1137,
    net1136,
    net1135,
    net1134,
    net1132,
    net1131,
    net1130,
    net1129,
    net1128,
    net1127,
    net1126,
    net1125,
    net1124,
    net1123,
    net1121,
    net1120,
    net1119,
    net1118,
    net1117,
    net1116,
    net1115,
    net1114,
    net1113,
    net1112,
    net1110,
    net1109,
    net1108,
    net1107,
    net1106,
    net1105,
    net1104,
    net1103,
    net1102,
    net1101,
    net1099,
    net1098,
    net1097,
    net1096,
    net1095,
    net1094,
    net1093,
    net1092,
    net1091,
    net1090,
    net1152,
    net1151,
    net1150,
    net1149,
    net1144,
    net1133,
    net1122,
    net1111,
    net1100,
    net1089}),
    .io_ins_up({\ces_0_0_io_outs_up[63] ,
    \ces_0_0_io_outs_up[62] ,
    \ces_0_0_io_outs_up[61] ,
    \ces_0_0_io_outs_up[60] ,
    \ces_0_0_io_outs_up[59] ,
    \ces_0_0_io_outs_up[58] ,
    \ces_0_0_io_outs_up[57] ,
    \ces_0_0_io_outs_up[56] ,
    \ces_0_0_io_outs_up[55] ,
    \ces_0_0_io_outs_up[54] ,
    \ces_0_0_io_outs_up[53] ,
    \ces_0_0_io_outs_up[52] ,
    \ces_0_0_io_outs_up[51] ,
    \ces_0_0_io_outs_up[50] ,
    \ces_0_0_io_outs_up[49] ,
    \ces_0_0_io_outs_up[48] ,
    \ces_0_0_io_outs_up[47] ,
    \ces_0_0_io_outs_up[46] ,
    \ces_0_0_io_outs_up[45] ,
    \ces_0_0_io_outs_up[44] ,
    \ces_0_0_io_outs_up[43] ,
    \ces_0_0_io_outs_up[42] ,
    \ces_0_0_io_outs_up[41] ,
    \ces_0_0_io_outs_up[40] ,
    \ces_0_0_io_outs_up[39] ,
    \ces_0_0_io_outs_up[38] ,
    \ces_0_0_io_outs_up[37] ,
    \ces_0_0_io_outs_up[36] ,
    \ces_0_0_io_outs_up[35] ,
    \ces_0_0_io_outs_up[34] ,
    \ces_0_0_io_outs_up[33] ,
    \ces_0_0_io_outs_up[32] ,
    \ces_0_0_io_outs_up[31] ,
    \ces_0_0_io_outs_up[30] ,
    \ces_0_0_io_outs_up[29] ,
    \ces_0_0_io_outs_up[28] ,
    \ces_0_0_io_outs_up[27] ,
    \ces_0_0_io_outs_up[26] ,
    \ces_0_0_io_outs_up[25] ,
    \ces_0_0_io_outs_up[24] ,
    \ces_0_0_io_outs_up[23] ,
    \ces_0_0_io_outs_up[22] ,
    \ces_0_0_io_outs_up[21] ,
    \ces_0_0_io_outs_up[20] ,
    \ces_0_0_io_outs_up[19] ,
    \ces_0_0_io_outs_up[18] ,
    \ces_0_0_io_outs_up[17] ,
    \ces_0_0_io_outs_up[16] ,
    \ces_0_0_io_outs_up[15] ,
    \ces_0_0_io_outs_up[14] ,
    \ces_0_0_io_outs_up[13] ,
    \ces_0_0_io_outs_up[12] ,
    \ces_0_0_io_outs_up[11] ,
    \ces_0_0_io_outs_up[10] ,
    \ces_0_0_io_outs_up[9] ,
    \ces_0_0_io_outs_up[8] ,
    \ces_0_0_io_outs_up[7] ,
    \ces_0_0_io_outs_up[6] ,
    \ces_0_0_io_outs_up[5] ,
    \ces_0_0_io_outs_up[4] ,
    \ces_0_0_io_outs_up[3] ,
    \ces_0_0_io_outs_up[2] ,
    \ces_0_0_io_outs_up[1] ,
    \ces_0_0_io_outs_up[0] }),
    .io_outs_down({\ces_0_0_io_ins_down[63] ,
    \ces_0_0_io_ins_down[62] ,
    \ces_0_0_io_ins_down[61] ,
    \ces_0_0_io_ins_down[60] ,
    \ces_0_0_io_ins_down[59] ,
    \ces_0_0_io_ins_down[58] ,
    \ces_0_0_io_ins_down[57] ,
    \ces_0_0_io_ins_down[56] ,
    \ces_0_0_io_ins_down[55] ,
    \ces_0_0_io_ins_down[54] ,
    \ces_0_0_io_ins_down[53] ,
    \ces_0_0_io_ins_down[52] ,
    \ces_0_0_io_ins_down[51] ,
    \ces_0_0_io_ins_down[50] ,
    \ces_0_0_io_ins_down[49] ,
    \ces_0_0_io_ins_down[48] ,
    \ces_0_0_io_ins_down[47] ,
    \ces_0_0_io_ins_down[46] ,
    \ces_0_0_io_ins_down[45] ,
    \ces_0_0_io_ins_down[44] ,
    \ces_0_0_io_ins_down[43] ,
    \ces_0_0_io_ins_down[42] ,
    \ces_0_0_io_ins_down[41] ,
    \ces_0_0_io_ins_down[40] ,
    \ces_0_0_io_ins_down[39] ,
    \ces_0_0_io_ins_down[38] ,
    \ces_0_0_io_ins_down[37] ,
    \ces_0_0_io_ins_down[36] ,
    \ces_0_0_io_ins_down[35] ,
    \ces_0_0_io_ins_down[34] ,
    \ces_0_0_io_ins_down[33] ,
    \ces_0_0_io_ins_down[32] ,
    \ces_0_0_io_ins_down[31] ,
    \ces_0_0_io_ins_down[30] ,
    \ces_0_0_io_ins_down[29] ,
    \ces_0_0_io_ins_down[28] ,
    \ces_0_0_io_ins_down[27] ,
    \ces_0_0_io_ins_down[26] ,
    \ces_0_0_io_ins_down[25] ,
    \ces_0_0_io_ins_down[24] ,
    \ces_0_0_io_ins_down[23] ,
    \ces_0_0_io_ins_down[22] ,
    \ces_0_0_io_ins_down[21] ,
    \ces_0_0_io_ins_down[20] ,
    \ces_0_0_io_ins_down[19] ,
    \ces_0_0_io_ins_down[18] ,
    \ces_0_0_io_ins_down[17] ,
    \ces_0_0_io_ins_down[16] ,
    \ces_0_0_io_ins_down[15] ,
    \ces_0_0_io_ins_down[14] ,
    \ces_0_0_io_ins_down[13] ,
    \ces_0_0_io_ins_down[12] ,
    \ces_0_0_io_ins_down[11] ,
    \ces_0_0_io_ins_down[10] ,
    \ces_0_0_io_ins_down[9] ,
    \ces_0_0_io_ins_down[8] ,
    \ces_0_0_io_ins_down[7] ,
    \ces_0_0_io_ins_down[6] ,
    \ces_0_0_io_ins_down[5] ,
    \ces_0_0_io_ins_down[4] ,
    \ces_0_0_io_ins_down[3] ,
    \ces_0_0_io_ins_down[2] ,
    \ces_0_0_io_ins_down[1] ,
    \ces_0_0_io_ins_down[0] }),
    .io_outs_left({net2748,
    net2747,
    net2746,
    net2745,
    net2743,
    net2742,
    net2741,
    net2740,
    net2739,
    net2738,
    net2737,
    net2736,
    net2735,
    net2734,
    net2732,
    net2731,
    net2730,
    net2729,
    net2728,
    net2727,
    net2726,
    net2725,
    net2724,
    net2723,
    net2721,
    net2720,
    net2719,
    net2718,
    net2717,
    net2716,
    net2715,
    net2714,
    net2713,
    net2712,
    net2710,
    net2709,
    net2708,
    net2707,
    net2706,
    net2705,
    net2704,
    net2703,
    net2702,
    net2701,
    net2699,
    net2698,
    net2697,
    net2696,
    net2695,
    net2694,
    net2693,
    net2692,
    net2691,
    net2690,
    net2752,
    net2751,
    net2750,
    net2749,
    net2744,
    net2733,
    net2722,
    net2711,
    net2700,
    net2689}),
    .io_outs_right({\ces_1_0_io_outs_right[63] ,
    \ces_1_0_io_outs_right[62] ,
    \ces_1_0_io_outs_right[61] ,
    \ces_1_0_io_outs_right[60] ,
    \ces_1_0_io_outs_right[59] ,
    \ces_1_0_io_outs_right[58] ,
    \ces_1_0_io_outs_right[57] ,
    \ces_1_0_io_outs_right[56] ,
    \ces_1_0_io_outs_right[55] ,
    \ces_1_0_io_outs_right[54] ,
    \ces_1_0_io_outs_right[53] ,
    \ces_1_0_io_outs_right[52] ,
    \ces_1_0_io_outs_right[51] ,
    \ces_1_0_io_outs_right[50] ,
    \ces_1_0_io_outs_right[49] ,
    \ces_1_0_io_outs_right[48] ,
    \ces_1_0_io_outs_right[47] ,
    \ces_1_0_io_outs_right[46] ,
    \ces_1_0_io_outs_right[45] ,
    \ces_1_0_io_outs_right[44] ,
    \ces_1_0_io_outs_right[43] ,
    \ces_1_0_io_outs_right[42] ,
    \ces_1_0_io_outs_right[41] ,
    \ces_1_0_io_outs_right[40] ,
    \ces_1_0_io_outs_right[39] ,
    \ces_1_0_io_outs_right[38] ,
    \ces_1_0_io_outs_right[37] ,
    \ces_1_0_io_outs_right[36] ,
    \ces_1_0_io_outs_right[35] ,
    \ces_1_0_io_outs_right[34] ,
    \ces_1_0_io_outs_right[33] ,
    \ces_1_0_io_outs_right[32] ,
    \ces_1_0_io_outs_right[31] ,
    \ces_1_0_io_outs_right[30] ,
    \ces_1_0_io_outs_right[29] ,
    \ces_1_0_io_outs_right[28] ,
    \ces_1_0_io_outs_right[27] ,
    \ces_1_0_io_outs_right[26] ,
    \ces_1_0_io_outs_right[25] ,
    \ces_1_0_io_outs_right[24] ,
    \ces_1_0_io_outs_right[23] ,
    \ces_1_0_io_outs_right[22] ,
    \ces_1_0_io_outs_right[21] ,
    \ces_1_0_io_outs_right[20] ,
    \ces_1_0_io_outs_right[19] ,
    \ces_1_0_io_outs_right[18] ,
    \ces_1_0_io_outs_right[17] ,
    \ces_1_0_io_outs_right[16] ,
    \ces_1_0_io_outs_right[15] ,
    \ces_1_0_io_outs_right[14] ,
    \ces_1_0_io_outs_right[13] ,
    \ces_1_0_io_outs_right[12] ,
    \ces_1_0_io_outs_right[11] ,
    \ces_1_0_io_outs_right[10] ,
    \ces_1_0_io_outs_right[9] ,
    \ces_1_0_io_outs_right[8] ,
    \ces_1_0_io_outs_right[7] ,
    \ces_1_0_io_outs_right[6] ,
    \ces_1_0_io_outs_right[5] ,
    \ces_1_0_io_outs_right[4] ,
    \ces_1_0_io_outs_right[3] ,
    \ces_1_0_io_outs_right[2] ,
    \ces_1_0_io_outs_right[1] ,
    \ces_1_0_io_outs_right[0] }),
    .io_outs_up({\ces_1_0_io_outs_up[63] ,
    \ces_1_0_io_outs_up[62] ,
    \ces_1_0_io_outs_up[61] ,
    \ces_1_0_io_outs_up[60] ,
    \ces_1_0_io_outs_up[59] ,
    \ces_1_0_io_outs_up[58] ,
    \ces_1_0_io_outs_up[57] ,
    \ces_1_0_io_outs_up[56] ,
    \ces_1_0_io_outs_up[55] ,
    \ces_1_0_io_outs_up[54] ,
    \ces_1_0_io_outs_up[53] ,
    \ces_1_0_io_outs_up[52] ,
    \ces_1_0_io_outs_up[51] ,
    \ces_1_0_io_outs_up[50] ,
    \ces_1_0_io_outs_up[49] ,
    \ces_1_0_io_outs_up[48] ,
    \ces_1_0_io_outs_up[47] ,
    \ces_1_0_io_outs_up[46] ,
    \ces_1_0_io_outs_up[45] ,
    \ces_1_0_io_outs_up[44] ,
    \ces_1_0_io_outs_up[43] ,
    \ces_1_0_io_outs_up[42] ,
    \ces_1_0_io_outs_up[41] ,
    \ces_1_0_io_outs_up[40] ,
    \ces_1_0_io_outs_up[39] ,
    \ces_1_0_io_outs_up[38] ,
    \ces_1_0_io_outs_up[37] ,
    \ces_1_0_io_outs_up[36] ,
    \ces_1_0_io_outs_up[35] ,
    \ces_1_0_io_outs_up[34] ,
    \ces_1_0_io_outs_up[33] ,
    \ces_1_0_io_outs_up[32] ,
    \ces_1_0_io_outs_up[31] ,
    \ces_1_0_io_outs_up[30] ,
    \ces_1_0_io_outs_up[29] ,
    \ces_1_0_io_outs_up[28] ,
    \ces_1_0_io_outs_up[27] ,
    \ces_1_0_io_outs_up[26] ,
    \ces_1_0_io_outs_up[25] ,
    \ces_1_0_io_outs_up[24] ,
    \ces_1_0_io_outs_up[23] ,
    \ces_1_0_io_outs_up[22] ,
    \ces_1_0_io_outs_up[21] ,
    \ces_1_0_io_outs_up[20] ,
    \ces_1_0_io_outs_up[19] ,
    \ces_1_0_io_outs_up[18] ,
    \ces_1_0_io_outs_up[17] ,
    \ces_1_0_io_outs_up[16] ,
    \ces_1_0_io_outs_up[15] ,
    \ces_1_0_io_outs_up[14] ,
    \ces_1_0_io_outs_up[13] ,
    \ces_1_0_io_outs_up[12] ,
    \ces_1_0_io_outs_up[11] ,
    \ces_1_0_io_outs_up[10] ,
    \ces_1_0_io_outs_up[9] ,
    \ces_1_0_io_outs_up[8] ,
    \ces_1_0_io_outs_up[7] ,
    \ces_1_0_io_outs_up[6] ,
    \ces_1_0_io_outs_up[5] ,
    \ces_1_0_io_outs_up[4] ,
    \ces_1_0_io_outs_up[3] ,
    \ces_1_0_io_outs_up[2] ,
    \ces_1_0_io_outs_up[1] ,
    \ces_1_0_io_outs_up[0] }));
 Element ces_1_1 (.clock(clknet_3_0_0_clock),
    .io_lsbIns_1(ces_1_0_io_lsbOuts_1),
    .io_lsbIns_2(ces_1_0_io_lsbOuts_2),
    .io_lsbIns_3(ces_1_0_io_lsbOuts_3),
    .io_lsbIns_4(ces_1_0_io_lsbOuts_4),
    .io_lsbIns_5(ces_1_0_io_lsbOuts_5),
    .io_lsbIns_6(ces_1_0_io_lsbOuts_6),
    .io_lsbIns_7(ces_1_0_io_lsbOuts_7),
    .io_lsbOuts_0(ces_1_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_1_io_lsbOuts_7),
    .io_ins_down({\ces_1_1_io_ins_down[63] ,
    \ces_1_1_io_ins_down[62] ,
    \ces_1_1_io_ins_down[61] ,
    \ces_1_1_io_ins_down[60] ,
    \ces_1_1_io_ins_down[59] ,
    \ces_1_1_io_ins_down[58] ,
    \ces_1_1_io_ins_down[57] ,
    \ces_1_1_io_ins_down[56] ,
    \ces_1_1_io_ins_down[55] ,
    \ces_1_1_io_ins_down[54] ,
    \ces_1_1_io_ins_down[53] ,
    \ces_1_1_io_ins_down[52] ,
    \ces_1_1_io_ins_down[51] ,
    \ces_1_1_io_ins_down[50] ,
    \ces_1_1_io_ins_down[49] ,
    \ces_1_1_io_ins_down[48] ,
    \ces_1_1_io_ins_down[47] ,
    \ces_1_1_io_ins_down[46] ,
    \ces_1_1_io_ins_down[45] ,
    \ces_1_1_io_ins_down[44] ,
    \ces_1_1_io_ins_down[43] ,
    \ces_1_1_io_ins_down[42] ,
    \ces_1_1_io_ins_down[41] ,
    \ces_1_1_io_ins_down[40] ,
    \ces_1_1_io_ins_down[39] ,
    \ces_1_1_io_ins_down[38] ,
    \ces_1_1_io_ins_down[37] ,
    \ces_1_1_io_ins_down[36] ,
    \ces_1_1_io_ins_down[35] ,
    \ces_1_1_io_ins_down[34] ,
    \ces_1_1_io_ins_down[33] ,
    \ces_1_1_io_ins_down[32] ,
    \ces_1_1_io_ins_down[31] ,
    \ces_1_1_io_ins_down[30] ,
    \ces_1_1_io_ins_down[29] ,
    \ces_1_1_io_ins_down[28] ,
    \ces_1_1_io_ins_down[27] ,
    \ces_1_1_io_ins_down[26] ,
    \ces_1_1_io_ins_down[25] ,
    \ces_1_1_io_ins_down[24] ,
    \ces_1_1_io_ins_down[23] ,
    \ces_1_1_io_ins_down[22] ,
    \ces_1_1_io_ins_down[21] ,
    \ces_1_1_io_ins_down[20] ,
    \ces_1_1_io_ins_down[19] ,
    \ces_1_1_io_ins_down[18] ,
    \ces_1_1_io_ins_down[17] ,
    \ces_1_1_io_ins_down[16] ,
    \ces_1_1_io_ins_down[15] ,
    \ces_1_1_io_ins_down[14] ,
    \ces_1_1_io_ins_down[13] ,
    \ces_1_1_io_ins_down[12] ,
    \ces_1_1_io_ins_down[11] ,
    \ces_1_1_io_ins_down[10] ,
    \ces_1_1_io_ins_down[9] ,
    \ces_1_1_io_ins_down[8] ,
    \ces_1_1_io_ins_down[7] ,
    \ces_1_1_io_ins_down[6] ,
    \ces_1_1_io_ins_down[5] ,
    \ces_1_1_io_ins_down[4] ,
    \ces_1_1_io_ins_down[3] ,
    \ces_1_1_io_ins_down[2] ,
    \ces_1_1_io_ins_down[1] ,
    \ces_1_1_io_ins_down[0] }),
    .io_ins_left({\ces_1_1_io_ins_left[63] ,
    \ces_1_1_io_ins_left[62] ,
    \ces_1_1_io_ins_left[61] ,
    \ces_1_1_io_ins_left[60] ,
    \ces_1_1_io_ins_left[59] ,
    \ces_1_1_io_ins_left[58] ,
    \ces_1_1_io_ins_left[57] ,
    \ces_1_1_io_ins_left[56] ,
    \ces_1_1_io_ins_left[55] ,
    \ces_1_1_io_ins_left[54] ,
    \ces_1_1_io_ins_left[53] ,
    \ces_1_1_io_ins_left[52] ,
    \ces_1_1_io_ins_left[51] ,
    \ces_1_1_io_ins_left[50] ,
    \ces_1_1_io_ins_left[49] ,
    \ces_1_1_io_ins_left[48] ,
    \ces_1_1_io_ins_left[47] ,
    \ces_1_1_io_ins_left[46] ,
    \ces_1_1_io_ins_left[45] ,
    \ces_1_1_io_ins_left[44] ,
    \ces_1_1_io_ins_left[43] ,
    \ces_1_1_io_ins_left[42] ,
    \ces_1_1_io_ins_left[41] ,
    \ces_1_1_io_ins_left[40] ,
    \ces_1_1_io_ins_left[39] ,
    \ces_1_1_io_ins_left[38] ,
    \ces_1_1_io_ins_left[37] ,
    \ces_1_1_io_ins_left[36] ,
    \ces_1_1_io_ins_left[35] ,
    \ces_1_1_io_ins_left[34] ,
    \ces_1_1_io_ins_left[33] ,
    \ces_1_1_io_ins_left[32] ,
    \ces_1_1_io_ins_left[31] ,
    \ces_1_1_io_ins_left[30] ,
    \ces_1_1_io_ins_left[29] ,
    \ces_1_1_io_ins_left[28] ,
    \ces_1_1_io_ins_left[27] ,
    \ces_1_1_io_ins_left[26] ,
    \ces_1_1_io_ins_left[25] ,
    \ces_1_1_io_ins_left[24] ,
    \ces_1_1_io_ins_left[23] ,
    \ces_1_1_io_ins_left[22] ,
    \ces_1_1_io_ins_left[21] ,
    \ces_1_1_io_ins_left[20] ,
    \ces_1_1_io_ins_left[19] ,
    \ces_1_1_io_ins_left[18] ,
    \ces_1_1_io_ins_left[17] ,
    \ces_1_1_io_ins_left[16] ,
    \ces_1_1_io_ins_left[15] ,
    \ces_1_1_io_ins_left[14] ,
    \ces_1_1_io_ins_left[13] ,
    \ces_1_1_io_ins_left[12] ,
    \ces_1_1_io_ins_left[11] ,
    \ces_1_1_io_ins_left[10] ,
    \ces_1_1_io_ins_left[9] ,
    \ces_1_1_io_ins_left[8] ,
    \ces_1_1_io_ins_left[7] ,
    \ces_1_1_io_ins_left[6] ,
    \ces_1_1_io_ins_left[5] ,
    \ces_1_1_io_ins_left[4] ,
    \ces_1_1_io_ins_left[3] ,
    \ces_1_1_io_ins_left[2] ,
    \ces_1_1_io_ins_left[1] ,
    \ces_1_1_io_ins_left[0] }),
    .io_ins_right({\ces_1_0_io_outs_right[63] ,
    \ces_1_0_io_outs_right[62] ,
    \ces_1_0_io_outs_right[61] ,
    \ces_1_0_io_outs_right[60] ,
    \ces_1_0_io_outs_right[59] ,
    \ces_1_0_io_outs_right[58] ,
    \ces_1_0_io_outs_right[57] ,
    \ces_1_0_io_outs_right[56] ,
    \ces_1_0_io_outs_right[55] ,
    \ces_1_0_io_outs_right[54] ,
    \ces_1_0_io_outs_right[53] ,
    \ces_1_0_io_outs_right[52] ,
    \ces_1_0_io_outs_right[51] ,
    \ces_1_0_io_outs_right[50] ,
    \ces_1_0_io_outs_right[49] ,
    \ces_1_0_io_outs_right[48] ,
    \ces_1_0_io_outs_right[47] ,
    \ces_1_0_io_outs_right[46] ,
    \ces_1_0_io_outs_right[45] ,
    \ces_1_0_io_outs_right[44] ,
    \ces_1_0_io_outs_right[43] ,
    \ces_1_0_io_outs_right[42] ,
    \ces_1_0_io_outs_right[41] ,
    \ces_1_0_io_outs_right[40] ,
    \ces_1_0_io_outs_right[39] ,
    \ces_1_0_io_outs_right[38] ,
    \ces_1_0_io_outs_right[37] ,
    \ces_1_0_io_outs_right[36] ,
    \ces_1_0_io_outs_right[35] ,
    \ces_1_0_io_outs_right[34] ,
    \ces_1_0_io_outs_right[33] ,
    \ces_1_0_io_outs_right[32] ,
    \ces_1_0_io_outs_right[31] ,
    \ces_1_0_io_outs_right[30] ,
    \ces_1_0_io_outs_right[29] ,
    \ces_1_0_io_outs_right[28] ,
    \ces_1_0_io_outs_right[27] ,
    \ces_1_0_io_outs_right[26] ,
    \ces_1_0_io_outs_right[25] ,
    \ces_1_0_io_outs_right[24] ,
    \ces_1_0_io_outs_right[23] ,
    \ces_1_0_io_outs_right[22] ,
    \ces_1_0_io_outs_right[21] ,
    \ces_1_0_io_outs_right[20] ,
    \ces_1_0_io_outs_right[19] ,
    \ces_1_0_io_outs_right[18] ,
    \ces_1_0_io_outs_right[17] ,
    \ces_1_0_io_outs_right[16] ,
    \ces_1_0_io_outs_right[15] ,
    \ces_1_0_io_outs_right[14] ,
    \ces_1_0_io_outs_right[13] ,
    \ces_1_0_io_outs_right[12] ,
    \ces_1_0_io_outs_right[11] ,
    \ces_1_0_io_outs_right[10] ,
    \ces_1_0_io_outs_right[9] ,
    \ces_1_0_io_outs_right[8] ,
    \ces_1_0_io_outs_right[7] ,
    \ces_1_0_io_outs_right[6] ,
    \ces_1_0_io_outs_right[5] ,
    \ces_1_0_io_outs_right[4] ,
    \ces_1_0_io_outs_right[3] ,
    \ces_1_0_io_outs_right[2] ,
    \ces_1_0_io_outs_right[1] ,
    \ces_1_0_io_outs_right[0] }),
    .io_ins_up({\ces_0_1_io_outs_up[63] ,
    \ces_0_1_io_outs_up[62] ,
    \ces_0_1_io_outs_up[61] ,
    \ces_0_1_io_outs_up[60] ,
    \ces_0_1_io_outs_up[59] ,
    \ces_0_1_io_outs_up[58] ,
    \ces_0_1_io_outs_up[57] ,
    \ces_0_1_io_outs_up[56] ,
    \ces_0_1_io_outs_up[55] ,
    \ces_0_1_io_outs_up[54] ,
    \ces_0_1_io_outs_up[53] ,
    \ces_0_1_io_outs_up[52] ,
    \ces_0_1_io_outs_up[51] ,
    \ces_0_1_io_outs_up[50] ,
    \ces_0_1_io_outs_up[49] ,
    \ces_0_1_io_outs_up[48] ,
    \ces_0_1_io_outs_up[47] ,
    \ces_0_1_io_outs_up[46] ,
    \ces_0_1_io_outs_up[45] ,
    \ces_0_1_io_outs_up[44] ,
    \ces_0_1_io_outs_up[43] ,
    \ces_0_1_io_outs_up[42] ,
    \ces_0_1_io_outs_up[41] ,
    \ces_0_1_io_outs_up[40] ,
    \ces_0_1_io_outs_up[39] ,
    \ces_0_1_io_outs_up[38] ,
    \ces_0_1_io_outs_up[37] ,
    \ces_0_1_io_outs_up[36] ,
    \ces_0_1_io_outs_up[35] ,
    \ces_0_1_io_outs_up[34] ,
    \ces_0_1_io_outs_up[33] ,
    \ces_0_1_io_outs_up[32] ,
    \ces_0_1_io_outs_up[31] ,
    \ces_0_1_io_outs_up[30] ,
    \ces_0_1_io_outs_up[29] ,
    \ces_0_1_io_outs_up[28] ,
    \ces_0_1_io_outs_up[27] ,
    \ces_0_1_io_outs_up[26] ,
    \ces_0_1_io_outs_up[25] ,
    \ces_0_1_io_outs_up[24] ,
    \ces_0_1_io_outs_up[23] ,
    \ces_0_1_io_outs_up[22] ,
    \ces_0_1_io_outs_up[21] ,
    \ces_0_1_io_outs_up[20] ,
    \ces_0_1_io_outs_up[19] ,
    \ces_0_1_io_outs_up[18] ,
    \ces_0_1_io_outs_up[17] ,
    \ces_0_1_io_outs_up[16] ,
    \ces_0_1_io_outs_up[15] ,
    \ces_0_1_io_outs_up[14] ,
    \ces_0_1_io_outs_up[13] ,
    \ces_0_1_io_outs_up[12] ,
    \ces_0_1_io_outs_up[11] ,
    \ces_0_1_io_outs_up[10] ,
    \ces_0_1_io_outs_up[9] ,
    \ces_0_1_io_outs_up[8] ,
    \ces_0_1_io_outs_up[7] ,
    \ces_0_1_io_outs_up[6] ,
    \ces_0_1_io_outs_up[5] ,
    \ces_0_1_io_outs_up[4] ,
    \ces_0_1_io_outs_up[3] ,
    \ces_0_1_io_outs_up[2] ,
    \ces_0_1_io_outs_up[1] ,
    \ces_0_1_io_outs_up[0] }),
    .io_outs_down({\ces_0_1_io_ins_down[63] ,
    \ces_0_1_io_ins_down[62] ,
    \ces_0_1_io_ins_down[61] ,
    \ces_0_1_io_ins_down[60] ,
    \ces_0_1_io_ins_down[59] ,
    \ces_0_1_io_ins_down[58] ,
    \ces_0_1_io_ins_down[57] ,
    \ces_0_1_io_ins_down[56] ,
    \ces_0_1_io_ins_down[55] ,
    \ces_0_1_io_ins_down[54] ,
    \ces_0_1_io_ins_down[53] ,
    \ces_0_1_io_ins_down[52] ,
    \ces_0_1_io_ins_down[51] ,
    \ces_0_1_io_ins_down[50] ,
    \ces_0_1_io_ins_down[49] ,
    \ces_0_1_io_ins_down[48] ,
    \ces_0_1_io_ins_down[47] ,
    \ces_0_1_io_ins_down[46] ,
    \ces_0_1_io_ins_down[45] ,
    \ces_0_1_io_ins_down[44] ,
    \ces_0_1_io_ins_down[43] ,
    \ces_0_1_io_ins_down[42] ,
    \ces_0_1_io_ins_down[41] ,
    \ces_0_1_io_ins_down[40] ,
    \ces_0_1_io_ins_down[39] ,
    \ces_0_1_io_ins_down[38] ,
    \ces_0_1_io_ins_down[37] ,
    \ces_0_1_io_ins_down[36] ,
    \ces_0_1_io_ins_down[35] ,
    \ces_0_1_io_ins_down[34] ,
    \ces_0_1_io_ins_down[33] ,
    \ces_0_1_io_ins_down[32] ,
    \ces_0_1_io_ins_down[31] ,
    \ces_0_1_io_ins_down[30] ,
    \ces_0_1_io_ins_down[29] ,
    \ces_0_1_io_ins_down[28] ,
    \ces_0_1_io_ins_down[27] ,
    \ces_0_1_io_ins_down[26] ,
    \ces_0_1_io_ins_down[25] ,
    \ces_0_1_io_ins_down[24] ,
    \ces_0_1_io_ins_down[23] ,
    \ces_0_1_io_ins_down[22] ,
    \ces_0_1_io_ins_down[21] ,
    \ces_0_1_io_ins_down[20] ,
    \ces_0_1_io_ins_down[19] ,
    \ces_0_1_io_ins_down[18] ,
    \ces_0_1_io_ins_down[17] ,
    \ces_0_1_io_ins_down[16] ,
    \ces_0_1_io_ins_down[15] ,
    \ces_0_1_io_ins_down[14] ,
    \ces_0_1_io_ins_down[13] ,
    \ces_0_1_io_ins_down[12] ,
    \ces_0_1_io_ins_down[11] ,
    \ces_0_1_io_ins_down[10] ,
    \ces_0_1_io_ins_down[9] ,
    \ces_0_1_io_ins_down[8] ,
    \ces_0_1_io_ins_down[7] ,
    \ces_0_1_io_ins_down[6] ,
    \ces_0_1_io_ins_down[5] ,
    \ces_0_1_io_ins_down[4] ,
    \ces_0_1_io_ins_down[3] ,
    \ces_0_1_io_ins_down[2] ,
    \ces_0_1_io_ins_down[1] ,
    \ces_0_1_io_ins_down[0] }),
    .io_outs_left({\ces_1_0_io_ins_left[63] ,
    \ces_1_0_io_ins_left[62] ,
    \ces_1_0_io_ins_left[61] ,
    \ces_1_0_io_ins_left[60] ,
    \ces_1_0_io_ins_left[59] ,
    \ces_1_0_io_ins_left[58] ,
    \ces_1_0_io_ins_left[57] ,
    \ces_1_0_io_ins_left[56] ,
    \ces_1_0_io_ins_left[55] ,
    \ces_1_0_io_ins_left[54] ,
    \ces_1_0_io_ins_left[53] ,
    \ces_1_0_io_ins_left[52] ,
    \ces_1_0_io_ins_left[51] ,
    \ces_1_0_io_ins_left[50] ,
    \ces_1_0_io_ins_left[49] ,
    \ces_1_0_io_ins_left[48] ,
    \ces_1_0_io_ins_left[47] ,
    \ces_1_0_io_ins_left[46] ,
    \ces_1_0_io_ins_left[45] ,
    \ces_1_0_io_ins_left[44] ,
    \ces_1_0_io_ins_left[43] ,
    \ces_1_0_io_ins_left[42] ,
    \ces_1_0_io_ins_left[41] ,
    \ces_1_0_io_ins_left[40] ,
    \ces_1_0_io_ins_left[39] ,
    \ces_1_0_io_ins_left[38] ,
    \ces_1_0_io_ins_left[37] ,
    \ces_1_0_io_ins_left[36] ,
    \ces_1_0_io_ins_left[35] ,
    \ces_1_0_io_ins_left[34] ,
    \ces_1_0_io_ins_left[33] ,
    \ces_1_0_io_ins_left[32] ,
    \ces_1_0_io_ins_left[31] ,
    \ces_1_0_io_ins_left[30] ,
    \ces_1_0_io_ins_left[29] ,
    \ces_1_0_io_ins_left[28] ,
    \ces_1_0_io_ins_left[27] ,
    \ces_1_0_io_ins_left[26] ,
    \ces_1_0_io_ins_left[25] ,
    \ces_1_0_io_ins_left[24] ,
    \ces_1_0_io_ins_left[23] ,
    \ces_1_0_io_ins_left[22] ,
    \ces_1_0_io_ins_left[21] ,
    \ces_1_0_io_ins_left[20] ,
    \ces_1_0_io_ins_left[19] ,
    \ces_1_0_io_ins_left[18] ,
    \ces_1_0_io_ins_left[17] ,
    \ces_1_0_io_ins_left[16] ,
    \ces_1_0_io_ins_left[15] ,
    \ces_1_0_io_ins_left[14] ,
    \ces_1_0_io_ins_left[13] ,
    \ces_1_0_io_ins_left[12] ,
    \ces_1_0_io_ins_left[11] ,
    \ces_1_0_io_ins_left[10] ,
    \ces_1_0_io_ins_left[9] ,
    \ces_1_0_io_ins_left[8] ,
    \ces_1_0_io_ins_left[7] ,
    \ces_1_0_io_ins_left[6] ,
    \ces_1_0_io_ins_left[5] ,
    \ces_1_0_io_ins_left[4] ,
    \ces_1_0_io_ins_left[3] ,
    \ces_1_0_io_ins_left[2] ,
    \ces_1_0_io_ins_left[1] ,
    \ces_1_0_io_ins_left[0] }),
    .io_outs_right({\ces_1_1_io_outs_right[63] ,
    \ces_1_1_io_outs_right[62] ,
    \ces_1_1_io_outs_right[61] ,
    \ces_1_1_io_outs_right[60] ,
    \ces_1_1_io_outs_right[59] ,
    \ces_1_1_io_outs_right[58] ,
    \ces_1_1_io_outs_right[57] ,
    \ces_1_1_io_outs_right[56] ,
    \ces_1_1_io_outs_right[55] ,
    \ces_1_1_io_outs_right[54] ,
    \ces_1_1_io_outs_right[53] ,
    \ces_1_1_io_outs_right[52] ,
    \ces_1_1_io_outs_right[51] ,
    \ces_1_1_io_outs_right[50] ,
    \ces_1_1_io_outs_right[49] ,
    \ces_1_1_io_outs_right[48] ,
    \ces_1_1_io_outs_right[47] ,
    \ces_1_1_io_outs_right[46] ,
    \ces_1_1_io_outs_right[45] ,
    \ces_1_1_io_outs_right[44] ,
    \ces_1_1_io_outs_right[43] ,
    \ces_1_1_io_outs_right[42] ,
    \ces_1_1_io_outs_right[41] ,
    \ces_1_1_io_outs_right[40] ,
    \ces_1_1_io_outs_right[39] ,
    \ces_1_1_io_outs_right[38] ,
    \ces_1_1_io_outs_right[37] ,
    \ces_1_1_io_outs_right[36] ,
    \ces_1_1_io_outs_right[35] ,
    \ces_1_1_io_outs_right[34] ,
    \ces_1_1_io_outs_right[33] ,
    \ces_1_1_io_outs_right[32] ,
    \ces_1_1_io_outs_right[31] ,
    \ces_1_1_io_outs_right[30] ,
    \ces_1_1_io_outs_right[29] ,
    \ces_1_1_io_outs_right[28] ,
    \ces_1_1_io_outs_right[27] ,
    \ces_1_1_io_outs_right[26] ,
    \ces_1_1_io_outs_right[25] ,
    \ces_1_1_io_outs_right[24] ,
    \ces_1_1_io_outs_right[23] ,
    \ces_1_1_io_outs_right[22] ,
    \ces_1_1_io_outs_right[21] ,
    \ces_1_1_io_outs_right[20] ,
    \ces_1_1_io_outs_right[19] ,
    \ces_1_1_io_outs_right[18] ,
    \ces_1_1_io_outs_right[17] ,
    \ces_1_1_io_outs_right[16] ,
    \ces_1_1_io_outs_right[15] ,
    \ces_1_1_io_outs_right[14] ,
    \ces_1_1_io_outs_right[13] ,
    \ces_1_1_io_outs_right[12] ,
    \ces_1_1_io_outs_right[11] ,
    \ces_1_1_io_outs_right[10] ,
    \ces_1_1_io_outs_right[9] ,
    \ces_1_1_io_outs_right[8] ,
    \ces_1_1_io_outs_right[7] ,
    \ces_1_1_io_outs_right[6] ,
    \ces_1_1_io_outs_right[5] ,
    \ces_1_1_io_outs_right[4] ,
    \ces_1_1_io_outs_right[3] ,
    \ces_1_1_io_outs_right[2] ,
    \ces_1_1_io_outs_right[1] ,
    \ces_1_1_io_outs_right[0] }),
    .io_outs_up({\ces_1_1_io_outs_up[63] ,
    \ces_1_1_io_outs_up[62] ,
    \ces_1_1_io_outs_up[61] ,
    \ces_1_1_io_outs_up[60] ,
    \ces_1_1_io_outs_up[59] ,
    \ces_1_1_io_outs_up[58] ,
    \ces_1_1_io_outs_up[57] ,
    \ces_1_1_io_outs_up[56] ,
    \ces_1_1_io_outs_up[55] ,
    \ces_1_1_io_outs_up[54] ,
    \ces_1_1_io_outs_up[53] ,
    \ces_1_1_io_outs_up[52] ,
    \ces_1_1_io_outs_up[51] ,
    \ces_1_1_io_outs_up[50] ,
    \ces_1_1_io_outs_up[49] ,
    \ces_1_1_io_outs_up[48] ,
    \ces_1_1_io_outs_up[47] ,
    \ces_1_1_io_outs_up[46] ,
    \ces_1_1_io_outs_up[45] ,
    \ces_1_1_io_outs_up[44] ,
    \ces_1_1_io_outs_up[43] ,
    \ces_1_1_io_outs_up[42] ,
    \ces_1_1_io_outs_up[41] ,
    \ces_1_1_io_outs_up[40] ,
    \ces_1_1_io_outs_up[39] ,
    \ces_1_1_io_outs_up[38] ,
    \ces_1_1_io_outs_up[37] ,
    \ces_1_1_io_outs_up[36] ,
    \ces_1_1_io_outs_up[35] ,
    \ces_1_1_io_outs_up[34] ,
    \ces_1_1_io_outs_up[33] ,
    \ces_1_1_io_outs_up[32] ,
    \ces_1_1_io_outs_up[31] ,
    \ces_1_1_io_outs_up[30] ,
    \ces_1_1_io_outs_up[29] ,
    \ces_1_1_io_outs_up[28] ,
    \ces_1_1_io_outs_up[27] ,
    \ces_1_1_io_outs_up[26] ,
    \ces_1_1_io_outs_up[25] ,
    \ces_1_1_io_outs_up[24] ,
    \ces_1_1_io_outs_up[23] ,
    \ces_1_1_io_outs_up[22] ,
    \ces_1_1_io_outs_up[21] ,
    \ces_1_1_io_outs_up[20] ,
    \ces_1_1_io_outs_up[19] ,
    \ces_1_1_io_outs_up[18] ,
    \ces_1_1_io_outs_up[17] ,
    \ces_1_1_io_outs_up[16] ,
    \ces_1_1_io_outs_up[15] ,
    \ces_1_1_io_outs_up[14] ,
    \ces_1_1_io_outs_up[13] ,
    \ces_1_1_io_outs_up[12] ,
    \ces_1_1_io_outs_up[11] ,
    \ces_1_1_io_outs_up[10] ,
    \ces_1_1_io_outs_up[9] ,
    \ces_1_1_io_outs_up[8] ,
    \ces_1_1_io_outs_up[7] ,
    \ces_1_1_io_outs_up[6] ,
    \ces_1_1_io_outs_up[5] ,
    \ces_1_1_io_outs_up[4] ,
    \ces_1_1_io_outs_up[3] ,
    \ces_1_1_io_outs_up[2] ,
    \ces_1_1_io_outs_up[1] ,
    \ces_1_1_io_outs_up[0] }));
 Element ces_1_2 (.clock(clknet_3_0_0_clock),
    .io_lsbIns_1(ces_1_1_io_lsbOuts_1),
    .io_lsbIns_2(ces_1_1_io_lsbOuts_2),
    .io_lsbIns_3(ces_1_1_io_lsbOuts_3),
    .io_lsbIns_4(ces_1_1_io_lsbOuts_4),
    .io_lsbIns_5(ces_1_1_io_lsbOuts_5),
    .io_lsbIns_6(ces_1_1_io_lsbOuts_6),
    .io_lsbIns_7(ces_1_1_io_lsbOuts_7),
    .io_lsbOuts_0(ces_1_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_2_io_lsbOuts_7),
    .io_ins_down({\ces_1_2_io_ins_down[63] ,
    \ces_1_2_io_ins_down[62] ,
    \ces_1_2_io_ins_down[61] ,
    \ces_1_2_io_ins_down[60] ,
    \ces_1_2_io_ins_down[59] ,
    \ces_1_2_io_ins_down[58] ,
    \ces_1_2_io_ins_down[57] ,
    \ces_1_2_io_ins_down[56] ,
    \ces_1_2_io_ins_down[55] ,
    \ces_1_2_io_ins_down[54] ,
    \ces_1_2_io_ins_down[53] ,
    \ces_1_2_io_ins_down[52] ,
    \ces_1_2_io_ins_down[51] ,
    \ces_1_2_io_ins_down[50] ,
    \ces_1_2_io_ins_down[49] ,
    \ces_1_2_io_ins_down[48] ,
    \ces_1_2_io_ins_down[47] ,
    \ces_1_2_io_ins_down[46] ,
    \ces_1_2_io_ins_down[45] ,
    \ces_1_2_io_ins_down[44] ,
    \ces_1_2_io_ins_down[43] ,
    \ces_1_2_io_ins_down[42] ,
    \ces_1_2_io_ins_down[41] ,
    \ces_1_2_io_ins_down[40] ,
    \ces_1_2_io_ins_down[39] ,
    \ces_1_2_io_ins_down[38] ,
    \ces_1_2_io_ins_down[37] ,
    \ces_1_2_io_ins_down[36] ,
    \ces_1_2_io_ins_down[35] ,
    \ces_1_2_io_ins_down[34] ,
    \ces_1_2_io_ins_down[33] ,
    \ces_1_2_io_ins_down[32] ,
    \ces_1_2_io_ins_down[31] ,
    \ces_1_2_io_ins_down[30] ,
    \ces_1_2_io_ins_down[29] ,
    \ces_1_2_io_ins_down[28] ,
    \ces_1_2_io_ins_down[27] ,
    \ces_1_2_io_ins_down[26] ,
    \ces_1_2_io_ins_down[25] ,
    \ces_1_2_io_ins_down[24] ,
    \ces_1_2_io_ins_down[23] ,
    \ces_1_2_io_ins_down[22] ,
    \ces_1_2_io_ins_down[21] ,
    \ces_1_2_io_ins_down[20] ,
    \ces_1_2_io_ins_down[19] ,
    \ces_1_2_io_ins_down[18] ,
    \ces_1_2_io_ins_down[17] ,
    \ces_1_2_io_ins_down[16] ,
    \ces_1_2_io_ins_down[15] ,
    \ces_1_2_io_ins_down[14] ,
    \ces_1_2_io_ins_down[13] ,
    \ces_1_2_io_ins_down[12] ,
    \ces_1_2_io_ins_down[11] ,
    \ces_1_2_io_ins_down[10] ,
    \ces_1_2_io_ins_down[9] ,
    \ces_1_2_io_ins_down[8] ,
    \ces_1_2_io_ins_down[7] ,
    \ces_1_2_io_ins_down[6] ,
    \ces_1_2_io_ins_down[5] ,
    \ces_1_2_io_ins_down[4] ,
    \ces_1_2_io_ins_down[3] ,
    \ces_1_2_io_ins_down[2] ,
    \ces_1_2_io_ins_down[1] ,
    \ces_1_2_io_ins_down[0] }),
    .io_ins_left({\ces_1_2_io_ins_left[63] ,
    \ces_1_2_io_ins_left[62] ,
    \ces_1_2_io_ins_left[61] ,
    \ces_1_2_io_ins_left[60] ,
    \ces_1_2_io_ins_left[59] ,
    \ces_1_2_io_ins_left[58] ,
    \ces_1_2_io_ins_left[57] ,
    \ces_1_2_io_ins_left[56] ,
    \ces_1_2_io_ins_left[55] ,
    \ces_1_2_io_ins_left[54] ,
    \ces_1_2_io_ins_left[53] ,
    \ces_1_2_io_ins_left[52] ,
    \ces_1_2_io_ins_left[51] ,
    \ces_1_2_io_ins_left[50] ,
    \ces_1_2_io_ins_left[49] ,
    \ces_1_2_io_ins_left[48] ,
    \ces_1_2_io_ins_left[47] ,
    \ces_1_2_io_ins_left[46] ,
    \ces_1_2_io_ins_left[45] ,
    \ces_1_2_io_ins_left[44] ,
    \ces_1_2_io_ins_left[43] ,
    \ces_1_2_io_ins_left[42] ,
    \ces_1_2_io_ins_left[41] ,
    \ces_1_2_io_ins_left[40] ,
    \ces_1_2_io_ins_left[39] ,
    \ces_1_2_io_ins_left[38] ,
    \ces_1_2_io_ins_left[37] ,
    \ces_1_2_io_ins_left[36] ,
    \ces_1_2_io_ins_left[35] ,
    \ces_1_2_io_ins_left[34] ,
    \ces_1_2_io_ins_left[33] ,
    \ces_1_2_io_ins_left[32] ,
    \ces_1_2_io_ins_left[31] ,
    \ces_1_2_io_ins_left[30] ,
    \ces_1_2_io_ins_left[29] ,
    \ces_1_2_io_ins_left[28] ,
    \ces_1_2_io_ins_left[27] ,
    \ces_1_2_io_ins_left[26] ,
    \ces_1_2_io_ins_left[25] ,
    \ces_1_2_io_ins_left[24] ,
    \ces_1_2_io_ins_left[23] ,
    \ces_1_2_io_ins_left[22] ,
    \ces_1_2_io_ins_left[21] ,
    \ces_1_2_io_ins_left[20] ,
    \ces_1_2_io_ins_left[19] ,
    \ces_1_2_io_ins_left[18] ,
    \ces_1_2_io_ins_left[17] ,
    \ces_1_2_io_ins_left[16] ,
    \ces_1_2_io_ins_left[15] ,
    \ces_1_2_io_ins_left[14] ,
    \ces_1_2_io_ins_left[13] ,
    \ces_1_2_io_ins_left[12] ,
    \ces_1_2_io_ins_left[11] ,
    \ces_1_2_io_ins_left[10] ,
    \ces_1_2_io_ins_left[9] ,
    \ces_1_2_io_ins_left[8] ,
    \ces_1_2_io_ins_left[7] ,
    \ces_1_2_io_ins_left[6] ,
    \ces_1_2_io_ins_left[5] ,
    \ces_1_2_io_ins_left[4] ,
    \ces_1_2_io_ins_left[3] ,
    \ces_1_2_io_ins_left[2] ,
    \ces_1_2_io_ins_left[1] ,
    \ces_1_2_io_ins_left[0] }),
    .io_ins_right({\ces_1_1_io_outs_right[63] ,
    \ces_1_1_io_outs_right[62] ,
    \ces_1_1_io_outs_right[61] ,
    \ces_1_1_io_outs_right[60] ,
    \ces_1_1_io_outs_right[59] ,
    \ces_1_1_io_outs_right[58] ,
    \ces_1_1_io_outs_right[57] ,
    \ces_1_1_io_outs_right[56] ,
    \ces_1_1_io_outs_right[55] ,
    \ces_1_1_io_outs_right[54] ,
    \ces_1_1_io_outs_right[53] ,
    \ces_1_1_io_outs_right[52] ,
    \ces_1_1_io_outs_right[51] ,
    \ces_1_1_io_outs_right[50] ,
    \ces_1_1_io_outs_right[49] ,
    \ces_1_1_io_outs_right[48] ,
    \ces_1_1_io_outs_right[47] ,
    \ces_1_1_io_outs_right[46] ,
    \ces_1_1_io_outs_right[45] ,
    \ces_1_1_io_outs_right[44] ,
    \ces_1_1_io_outs_right[43] ,
    \ces_1_1_io_outs_right[42] ,
    \ces_1_1_io_outs_right[41] ,
    \ces_1_1_io_outs_right[40] ,
    \ces_1_1_io_outs_right[39] ,
    \ces_1_1_io_outs_right[38] ,
    \ces_1_1_io_outs_right[37] ,
    \ces_1_1_io_outs_right[36] ,
    \ces_1_1_io_outs_right[35] ,
    \ces_1_1_io_outs_right[34] ,
    \ces_1_1_io_outs_right[33] ,
    \ces_1_1_io_outs_right[32] ,
    \ces_1_1_io_outs_right[31] ,
    \ces_1_1_io_outs_right[30] ,
    \ces_1_1_io_outs_right[29] ,
    \ces_1_1_io_outs_right[28] ,
    \ces_1_1_io_outs_right[27] ,
    \ces_1_1_io_outs_right[26] ,
    \ces_1_1_io_outs_right[25] ,
    \ces_1_1_io_outs_right[24] ,
    \ces_1_1_io_outs_right[23] ,
    \ces_1_1_io_outs_right[22] ,
    \ces_1_1_io_outs_right[21] ,
    \ces_1_1_io_outs_right[20] ,
    \ces_1_1_io_outs_right[19] ,
    \ces_1_1_io_outs_right[18] ,
    \ces_1_1_io_outs_right[17] ,
    \ces_1_1_io_outs_right[16] ,
    \ces_1_1_io_outs_right[15] ,
    \ces_1_1_io_outs_right[14] ,
    \ces_1_1_io_outs_right[13] ,
    \ces_1_1_io_outs_right[12] ,
    \ces_1_1_io_outs_right[11] ,
    \ces_1_1_io_outs_right[10] ,
    \ces_1_1_io_outs_right[9] ,
    \ces_1_1_io_outs_right[8] ,
    \ces_1_1_io_outs_right[7] ,
    \ces_1_1_io_outs_right[6] ,
    \ces_1_1_io_outs_right[5] ,
    \ces_1_1_io_outs_right[4] ,
    \ces_1_1_io_outs_right[3] ,
    \ces_1_1_io_outs_right[2] ,
    \ces_1_1_io_outs_right[1] ,
    \ces_1_1_io_outs_right[0] }),
    .io_ins_up({\ces_0_2_io_outs_up[63] ,
    \ces_0_2_io_outs_up[62] ,
    \ces_0_2_io_outs_up[61] ,
    \ces_0_2_io_outs_up[60] ,
    \ces_0_2_io_outs_up[59] ,
    \ces_0_2_io_outs_up[58] ,
    \ces_0_2_io_outs_up[57] ,
    \ces_0_2_io_outs_up[56] ,
    \ces_0_2_io_outs_up[55] ,
    \ces_0_2_io_outs_up[54] ,
    \ces_0_2_io_outs_up[53] ,
    \ces_0_2_io_outs_up[52] ,
    \ces_0_2_io_outs_up[51] ,
    \ces_0_2_io_outs_up[50] ,
    \ces_0_2_io_outs_up[49] ,
    \ces_0_2_io_outs_up[48] ,
    \ces_0_2_io_outs_up[47] ,
    \ces_0_2_io_outs_up[46] ,
    \ces_0_2_io_outs_up[45] ,
    \ces_0_2_io_outs_up[44] ,
    \ces_0_2_io_outs_up[43] ,
    \ces_0_2_io_outs_up[42] ,
    \ces_0_2_io_outs_up[41] ,
    \ces_0_2_io_outs_up[40] ,
    \ces_0_2_io_outs_up[39] ,
    \ces_0_2_io_outs_up[38] ,
    \ces_0_2_io_outs_up[37] ,
    \ces_0_2_io_outs_up[36] ,
    \ces_0_2_io_outs_up[35] ,
    \ces_0_2_io_outs_up[34] ,
    \ces_0_2_io_outs_up[33] ,
    \ces_0_2_io_outs_up[32] ,
    \ces_0_2_io_outs_up[31] ,
    \ces_0_2_io_outs_up[30] ,
    \ces_0_2_io_outs_up[29] ,
    \ces_0_2_io_outs_up[28] ,
    \ces_0_2_io_outs_up[27] ,
    \ces_0_2_io_outs_up[26] ,
    \ces_0_2_io_outs_up[25] ,
    \ces_0_2_io_outs_up[24] ,
    \ces_0_2_io_outs_up[23] ,
    \ces_0_2_io_outs_up[22] ,
    \ces_0_2_io_outs_up[21] ,
    \ces_0_2_io_outs_up[20] ,
    \ces_0_2_io_outs_up[19] ,
    \ces_0_2_io_outs_up[18] ,
    \ces_0_2_io_outs_up[17] ,
    \ces_0_2_io_outs_up[16] ,
    \ces_0_2_io_outs_up[15] ,
    \ces_0_2_io_outs_up[14] ,
    \ces_0_2_io_outs_up[13] ,
    \ces_0_2_io_outs_up[12] ,
    \ces_0_2_io_outs_up[11] ,
    \ces_0_2_io_outs_up[10] ,
    \ces_0_2_io_outs_up[9] ,
    \ces_0_2_io_outs_up[8] ,
    \ces_0_2_io_outs_up[7] ,
    \ces_0_2_io_outs_up[6] ,
    \ces_0_2_io_outs_up[5] ,
    \ces_0_2_io_outs_up[4] ,
    \ces_0_2_io_outs_up[3] ,
    \ces_0_2_io_outs_up[2] ,
    \ces_0_2_io_outs_up[1] ,
    \ces_0_2_io_outs_up[0] }),
    .io_outs_down({\ces_0_2_io_ins_down[63] ,
    \ces_0_2_io_ins_down[62] ,
    \ces_0_2_io_ins_down[61] ,
    \ces_0_2_io_ins_down[60] ,
    \ces_0_2_io_ins_down[59] ,
    \ces_0_2_io_ins_down[58] ,
    \ces_0_2_io_ins_down[57] ,
    \ces_0_2_io_ins_down[56] ,
    \ces_0_2_io_ins_down[55] ,
    \ces_0_2_io_ins_down[54] ,
    \ces_0_2_io_ins_down[53] ,
    \ces_0_2_io_ins_down[52] ,
    \ces_0_2_io_ins_down[51] ,
    \ces_0_2_io_ins_down[50] ,
    \ces_0_2_io_ins_down[49] ,
    \ces_0_2_io_ins_down[48] ,
    \ces_0_2_io_ins_down[47] ,
    \ces_0_2_io_ins_down[46] ,
    \ces_0_2_io_ins_down[45] ,
    \ces_0_2_io_ins_down[44] ,
    \ces_0_2_io_ins_down[43] ,
    \ces_0_2_io_ins_down[42] ,
    \ces_0_2_io_ins_down[41] ,
    \ces_0_2_io_ins_down[40] ,
    \ces_0_2_io_ins_down[39] ,
    \ces_0_2_io_ins_down[38] ,
    \ces_0_2_io_ins_down[37] ,
    \ces_0_2_io_ins_down[36] ,
    \ces_0_2_io_ins_down[35] ,
    \ces_0_2_io_ins_down[34] ,
    \ces_0_2_io_ins_down[33] ,
    \ces_0_2_io_ins_down[32] ,
    \ces_0_2_io_ins_down[31] ,
    \ces_0_2_io_ins_down[30] ,
    \ces_0_2_io_ins_down[29] ,
    \ces_0_2_io_ins_down[28] ,
    \ces_0_2_io_ins_down[27] ,
    \ces_0_2_io_ins_down[26] ,
    \ces_0_2_io_ins_down[25] ,
    \ces_0_2_io_ins_down[24] ,
    \ces_0_2_io_ins_down[23] ,
    \ces_0_2_io_ins_down[22] ,
    \ces_0_2_io_ins_down[21] ,
    \ces_0_2_io_ins_down[20] ,
    \ces_0_2_io_ins_down[19] ,
    \ces_0_2_io_ins_down[18] ,
    \ces_0_2_io_ins_down[17] ,
    \ces_0_2_io_ins_down[16] ,
    \ces_0_2_io_ins_down[15] ,
    \ces_0_2_io_ins_down[14] ,
    \ces_0_2_io_ins_down[13] ,
    \ces_0_2_io_ins_down[12] ,
    \ces_0_2_io_ins_down[11] ,
    \ces_0_2_io_ins_down[10] ,
    \ces_0_2_io_ins_down[9] ,
    \ces_0_2_io_ins_down[8] ,
    \ces_0_2_io_ins_down[7] ,
    \ces_0_2_io_ins_down[6] ,
    \ces_0_2_io_ins_down[5] ,
    \ces_0_2_io_ins_down[4] ,
    \ces_0_2_io_ins_down[3] ,
    \ces_0_2_io_ins_down[2] ,
    \ces_0_2_io_ins_down[1] ,
    \ces_0_2_io_ins_down[0] }),
    .io_outs_left({\ces_1_1_io_ins_left[63] ,
    \ces_1_1_io_ins_left[62] ,
    \ces_1_1_io_ins_left[61] ,
    \ces_1_1_io_ins_left[60] ,
    \ces_1_1_io_ins_left[59] ,
    \ces_1_1_io_ins_left[58] ,
    \ces_1_1_io_ins_left[57] ,
    \ces_1_1_io_ins_left[56] ,
    \ces_1_1_io_ins_left[55] ,
    \ces_1_1_io_ins_left[54] ,
    \ces_1_1_io_ins_left[53] ,
    \ces_1_1_io_ins_left[52] ,
    \ces_1_1_io_ins_left[51] ,
    \ces_1_1_io_ins_left[50] ,
    \ces_1_1_io_ins_left[49] ,
    \ces_1_1_io_ins_left[48] ,
    \ces_1_1_io_ins_left[47] ,
    \ces_1_1_io_ins_left[46] ,
    \ces_1_1_io_ins_left[45] ,
    \ces_1_1_io_ins_left[44] ,
    \ces_1_1_io_ins_left[43] ,
    \ces_1_1_io_ins_left[42] ,
    \ces_1_1_io_ins_left[41] ,
    \ces_1_1_io_ins_left[40] ,
    \ces_1_1_io_ins_left[39] ,
    \ces_1_1_io_ins_left[38] ,
    \ces_1_1_io_ins_left[37] ,
    \ces_1_1_io_ins_left[36] ,
    \ces_1_1_io_ins_left[35] ,
    \ces_1_1_io_ins_left[34] ,
    \ces_1_1_io_ins_left[33] ,
    \ces_1_1_io_ins_left[32] ,
    \ces_1_1_io_ins_left[31] ,
    \ces_1_1_io_ins_left[30] ,
    \ces_1_1_io_ins_left[29] ,
    \ces_1_1_io_ins_left[28] ,
    \ces_1_1_io_ins_left[27] ,
    \ces_1_1_io_ins_left[26] ,
    \ces_1_1_io_ins_left[25] ,
    \ces_1_1_io_ins_left[24] ,
    \ces_1_1_io_ins_left[23] ,
    \ces_1_1_io_ins_left[22] ,
    \ces_1_1_io_ins_left[21] ,
    \ces_1_1_io_ins_left[20] ,
    \ces_1_1_io_ins_left[19] ,
    \ces_1_1_io_ins_left[18] ,
    \ces_1_1_io_ins_left[17] ,
    \ces_1_1_io_ins_left[16] ,
    \ces_1_1_io_ins_left[15] ,
    \ces_1_1_io_ins_left[14] ,
    \ces_1_1_io_ins_left[13] ,
    \ces_1_1_io_ins_left[12] ,
    \ces_1_1_io_ins_left[11] ,
    \ces_1_1_io_ins_left[10] ,
    \ces_1_1_io_ins_left[9] ,
    \ces_1_1_io_ins_left[8] ,
    \ces_1_1_io_ins_left[7] ,
    \ces_1_1_io_ins_left[6] ,
    \ces_1_1_io_ins_left[5] ,
    \ces_1_1_io_ins_left[4] ,
    \ces_1_1_io_ins_left[3] ,
    \ces_1_1_io_ins_left[2] ,
    \ces_1_1_io_ins_left[1] ,
    \ces_1_1_io_ins_left[0] }),
    .io_outs_right({\ces_1_2_io_outs_right[63] ,
    \ces_1_2_io_outs_right[62] ,
    \ces_1_2_io_outs_right[61] ,
    \ces_1_2_io_outs_right[60] ,
    \ces_1_2_io_outs_right[59] ,
    \ces_1_2_io_outs_right[58] ,
    \ces_1_2_io_outs_right[57] ,
    \ces_1_2_io_outs_right[56] ,
    \ces_1_2_io_outs_right[55] ,
    \ces_1_2_io_outs_right[54] ,
    \ces_1_2_io_outs_right[53] ,
    \ces_1_2_io_outs_right[52] ,
    \ces_1_2_io_outs_right[51] ,
    \ces_1_2_io_outs_right[50] ,
    \ces_1_2_io_outs_right[49] ,
    \ces_1_2_io_outs_right[48] ,
    \ces_1_2_io_outs_right[47] ,
    \ces_1_2_io_outs_right[46] ,
    \ces_1_2_io_outs_right[45] ,
    \ces_1_2_io_outs_right[44] ,
    \ces_1_2_io_outs_right[43] ,
    \ces_1_2_io_outs_right[42] ,
    \ces_1_2_io_outs_right[41] ,
    \ces_1_2_io_outs_right[40] ,
    \ces_1_2_io_outs_right[39] ,
    \ces_1_2_io_outs_right[38] ,
    \ces_1_2_io_outs_right[37] ,
    \ces_1_2_io_outs_right[36] ,
    \ces_1_2_io_outs_right[35] ,
    \ces_1_2_io_outs_right[34] ,
    \ces_1_2_io_outs_right[33] ,
    \ces_1_2_io_outs_right[32] ,
    \ces_1_2_io_outs_right[31] ,
    \ces_1_2_io_outs_right[30] ,
    \ces_1_2_io_outs_right[29] ,
    \ces_1_2_io_outs_right[28] ,
    \ces_1_2_io_outs_right[27] ,
    \ces_1_2_io_outs_right[26] ,
    \ces_1_2_io_outs_right[25] ,
    \ces_1_2_io_outs_right[24] ,
    \ces_1_2_io_outs_right[23] ,
    \ces_1_2_io_outs_right[22] ,
    \ces_1_2_io_outs_right[21] ,
    \ces_1_2_io_outs_right[20] ,
    \ces_1_2_io_outs_right[19] ,
    \ces_1_2_io_outs_right[18] ,
    \ces_1_2_io_outs_right[17] ,
    \ces_1_2_io_outs_right[16] ,
    \ces_1_2_io_outs_right[15] ,
    \ces_1_2_io_outs_right[14] ,
    \ces_1_2_io_outs_right[13] ,
    \ces_1_2_io_outs_right[12] ,
    \ces_1_2_io_outs_right[11] ,
    \ces_1_2_io_outs_right[10] ,
    \ces_1_2_io_outs_right[9] ,
    \ces_1_2_io_outs_right[8] ,
    \ces_1_2_io_outs_right[7] ,
    \ces_1_2_io_outs_right[6] ,
    \ces_1_2_io_outs_right[5] ,
    \ces_1_2_io_outs_right[4] ,
    \ces_1_2_io_outs_right[3] ,
    \ces_1_2_io_outs_right[2] ,
    \ces_1_2_io_outs_right[1] ,
    \ces_1_2_io_outs_right[0] }),
    .io_outs_up({\ces_1_2_io_outs_up[63] ,
    \ces_1_2_io_outs_up[62] ,
    \ces_1_2_io_outs_up[61] ,
    \ces_1_2_io_outs_up[60] ,
    \ces_1_2_io_outs_up[59] ,
    \ces_1_2_io_outs_up[58] ,
    \ces_1_2_io_outs_up[57] ,
    \ces_1_2_io_outs_up[56] ,
    \ces_1_2_io_outs_up[55] ,
    \ces_1_2_io_outs_up[54] ,
    \ces_1_2_io_outs_up[53] ,
    \ces_1_2_io_outs_up[52] ,
    \ces_1_2_io_outs_up[51] ,
    \ces_1_2_io_outs_up[50] ,
    \ces_1_2_io_outs_up[49] ,
    \ces_1_2_io_outs_up[48] ,
    \ces_1_2_io_outs_up[47] ,
    \ces_1_2_io_outs_up[46] ,
    \ces_1_2_io_outs_up[45] ,
    \ces_1_2_io_outs_up[44] ,
    \ces_1_2_io_outs_up[43] ,
    \ces_1_2_io_outs_up[42] ,
    \ces_1_2_io_outs_up[41] ,
    \ces_1_2_io_outs_up[40] ,
    \ces_1_2_io_outs_up[39] ,
    \ces_1_2_io_outs_up[38] ,
    \ces_1_2_io_outs_up[37] ,
    \ces_1_2_io_outs_up[36] ,
    \ces_1_2_io_outs_up[35] ,
    \ces_1_2_io_outs_up[34] ,
    \ces_1_2_io_outs_up[33] ,
    \ces_1_2_io_outs_up[32] ,
    \ces_1_2_io_outs_up[31] ,
    \ces_1_2_io_outs_up[30] ,
    \ces_1_2_io_outs_up[29] ,
    \ces_1_2_io_outs_up[28] ,
    \ces_1_2_io_outs_up[27] ,
    \ces_1_2_io_outs_up[26] ,
    \ces_1_2_io_outs_up[25] ,
    \ces_1_2_io_outs_up[24] ,
    \ces_1_2_io_outs_up[23] ,
    \ces_1_2_io_outs_up[22] ,
    \ces_1_2_io_outs_up[21] ,
    \ces_1_2_io_outs_up[20] ,
    \ces_1_2_io_outs_up[19] ,
    \ces_1_2_io_outs_up[18] ,
    \ces_1_2_io_outs_up[17] ,
    \ces_1_2_io_outs_up[16] ,
    \ces_1_2_io_outs_up[15] ,
    \ces_1_2_io_outs_up[14] ,
    \ces_1_2_io_outs_up[13] ,
    \ces_1_2_io_outs_up[12] ,
    \ces_1_2_io_outs_up[11] ,
    \ces_1_2_io_outs_up[10] ,
    \ces_1_2_io_outs_up[9] ,
    \ces_1_2_io_outs_up[8] ,
    \ces_1_2_io_outs_up[7] ,
    \ces_1_2_io_outs_up[6] ,
    \ces_1_2_io_outs_up[5] ,
    \ces_1_2_io_outs_up[4] ,
    \ces_1_2_io_outs_up[3] ,
    \ces_1_2_io_outs_up[2] ,
    \ces_1_2_io_outs_up[1] ,
    \ces_1_2_io_outs_up[0] }));
 Element ces_1_3 (.clock(clknet_3_0_0_clock),
    .io_lsbIns_1(ces_1_2_io_lsbOuts_1),
    .io_lsbIns_2(ces_1_2_io_lsbOuts_2),
    .io_lsbIns_3(ces_1_2_io_lsbOuts_3),
    .io_lsbIns_4(ces_1_2_io_lsbOuts_4),
    .io_lsbIns_5(ces_1_2_io_lsbOuts_5),
    .io_lsbIns_6(ces_1_2_io_lsbOuts_6),
    .io_lsbIns_7(ces_1_2_io_lsbOuts_7),
    .io_lsbOuts_0(ces_1_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_3_io_lsbOuts_7),
    .io_ins_down({\ces_1_3_io_ins_down[63] ,
    \ces_1_3_io_ins_down[62] ,
    \ces_1_3_io_ins_down[61] ,
    \ces_1_3_io_ins_down[60] ,
    \ces_1_3_io_ins_down[59] ,
    \ces_1_3_io_ins_down[58] ,
    \ces_1_3_io_ins_down[57] ,
    \ces_1_3_io_ins_down[56] ,
    \ces_1_3_io_ins_down[55] ,
    \ces_1_3_io_ins_down[54] ,
    \ces_1_3_io_ins_down[53] ,
    \ces_1_3_io_ins_down[52] ,
    \ces_1_3_io_ins_down[51] ,
    \ces_1_3_io_ins_down[50] ,
    \ces_1_3_io_ins_down[49] ,
    \ces_1_3_io_ins_down[48] ,
    \ces_1_3_io_ins_down[47] ,
    \ces_1_3_io_ins_down[46] ,
    \ces_1_3_io_ins_down[45] ,
    \ces_1_3_io_ins_down[44] ,
    \ces_1_3_io_ins_down[43] ,
    \ces_1_3_io_ins_down[42] ,
    \ces_1_3_io_ins_down[41] ,
    \ces_1_3_io_ins_down[40] ,
    \ces_1_3_io_ins_down[39] ,
    \ces_1_3_io_ins_down[38] ,
    \ces_1_3_io_ins_down[37] ,
    \ces_1_3_io_ins_down[36] ,
    \ces_1_3_io_ins_down[35] ,
    \ces_1_3_io_ins_down[34] ,
    \ces_1_3_io_ins_down[33] ,
    \ces_1_3_io_ins_down[32] ,
    \ces_1_3_io_ins_down[31] ,
    \ces_1_3_io_ins_down[30] ,
    \ces_1_3_io_ins_down[29] ,
    \ces_1_3_io_ins_down[28] ,
    \ces_1_3_io_ins_down[27] ,
    \ces_1_3_io_ins_down[26] ,
    \ces_1_3_io_ins_down[25] ,
    \ces_1_3_io_ins_down[24] ,
    \ces_1_3_io_ins_down[23] ,
    \ces_1_3_io_ins_down[22] ,
    \ces_1_3_io_ins_down[21] ,
    \ces_1_3_io_ins_down[20] ,
    \ces_1_3_io_ins_down[19] ,
    \ces_1_3_io_ins_down[18] ,
    \ces_1_3_io_ins_down[17] ,
    \ces_1_3_io_ins_down[16] ,
    \ces_1_3_io_ins_down[15] ,
    \ces_1_3_io_ins_down[14] ,
    \ces_1_3_io_ins_down[13] ,
    \ces_1_3_io_ins_down[12] ,
    \ces_1_3_io_ins_down[11] ,
    \ces_1_3_io_ins_down[10] ,
    \ces_1_3_io_ins_down[9] ,
    \ces_1_3_io_ins_down[8] ,
    \ces_1_3_io_ins_down[7] ,
    \ces_1_3_io_ins_down[6] ,
    \ces_1_3_io_ins_down[5] ,
    \ces_1_3_io_ins_down[4] ,
    \ces_1_3_io_ins_down[3] ,
    \ces_1_3_io_ins_down[2] ,
    \ces_1_3_io_ins_down[1] ,
    \ces_1_3_io_ins_down[0] }),
    .io_ins_left({\ces_1_3_io_ins_left[63] ,
    \ces_1_3_io_ins_left[62] ,
    \ces_1_3_io_ins_left[61] ,
    \ces_1_3_io_ins_left[60] ,
    \ces_1_3_io_ins_left[59] ,
    \ces_1_3_io_ins_left[58] ,
    \ces_1_3_io_ins_left[57] ,
    \ces_1_3_io_ins_left[56] ,
    \ces_1_3_io_ins_left[55] ,
    \ces_1_3_io_ins_left[54] ,
    \ces_1_3_io_ins_left[53] ,
    \ces_1_3_io_ins_left[52] ,
    \ces_1_3_io_ins_left[51] ,
    \ces_1_3_io_ins_left[50] ,
    \ces_1_3_io_ins_left[49] ,
    \ces_1_3_io_ins_left[48] ,
    \ces_1_3_io_ins_left[47] ,
    \ces_1_3_io_ins_left[46] ,
    \ces_1_3_io_ins_left[45] ,
    \ces_1_3_io_ins_left[44] ,
    \ces_1_3_io_ins_left[43] ,
    \ces_1_3_io_ins_left[42] ,
    \ces_1_3_io_ins_left[41] ,
    \ces_1_3_io_ins_left[40] ,
    \ces_1_3_io_ins_left[39] ,
    \ces_1_3_io_ins_left[38] ,
    \ces_1_3_io_ins_left[37] ,
    \ces_1_3_io_ins_left[36] ,
    \ces_1_3_io_ins_left[35] ,
    \ces_1_3_io_ins_left[34] ,
    \ces_1_3_io_ins_left[33] ,
    \ces_1_3_io_ins_left[32] ,
    \ces_1_3_io_ins_left[31] ,
    \ces_1_3_io_ins_left[30] ,
    \ces_1_3_io_ins_left[29] ,
    \ces_1_3_io_ins_left[28] ,
    \ces_1_3_io_ins_left[27] ,
    \ces_1_3_io_ins_left[26] ,
    \ces_1_3_io_ins_left[25] ,
    \ces_1_3_io_ins_left[24] ,
    \ces_1_3_io_ins_left[23] ,
    \ces_1_3_io_ins_left[22] ,
    \ces_1_3_io_ins_left[21] ,
    \ces_1_3_io_ins_left[20] ,
    \ces_1_3_io_ins_left[19] ,
    \ces_1_3_io_ins_left[18] ,
    \ces_1_3_io_ins_left[17] ,
    \ces_1_3_io_ins_left[16] ,
    \ces_1_3_io_ins_left[15] ,
    \ces_1_3_io_ins_left[14] ,
    \ces_1_3_io_ins_left[13] ,
    \ces_1_3_io_ins_left[12] ,
    \ces_1_3_io_ins_left[11] ,
    \ces_1_3_io_ins_left[10] ,
    \ces_1_3_io_ins_left[9] ,
    \ces_1_3_io_ins_left[8] ,
    \ces_1_3_io_ins_left[7] ,
    \ces_1_3_io_ins_left[6] ,
    \ces_1_3_io_ins_left[5] ,
    \ces_1_3_io_ins_left[4] ,
    \ces_1_3_io_ins_left[3] ,
    \ces_1_3_io_ins_left[2] ,
    \ces_1_3_io_ins_left[1] ,
    \ces_1_3_io_ins_left[0] }),
    .io_ins_right({\ces_1_2_io_outs_right[63] ,
    \ces_1_2_io_outs_right[62] ,
    \ces_1_2_io_outs_right[61] ,
    \ces_1_2_io_outs_right[60] ,
    \ces_1_2_io_outs_right[59] ,
    \ces_1_2_io_outs_right[58] ,
    \ces_1_2_io_outs_right[57] ,
    \ces_1_2_io_outs_right[56] ,
    \ces_1_2_io_outs_right[55] ,
    \ces_1_2_io_outs_right[54] ,
    \ces_1_2_io_outs_right[53] ,
    \ces_1_2_io_outs_right[52] ,
    \ces_1_2_io_outs_right[51] ,
    \ces_1_2_io_outs_right[50] ,
    \ces_1_2_io_outs_right[49] ,
    \ces_1_2_io_outs_right[48] ,
    \ces_1_2_io_outs_right[47] ,
    \ces_1_2_io_outs_right[46] ,
    \ces_1_2_io_outs_right[45] ,
    \ces_1_2_io_outs_right[44] ,
    \ces_1_2_io_outs_right[43] ,
    \ces_1_2_io_outs_right[42] ,
    \ces_1_2_io_outs_right[41] ,
    \ces_1_2_io_outs_right[40] ,
    \ces_1_2_io_outs_right[39] ,
    \ces_1_2_io_outs_right[38] ,
    \ces_1_2_io_outs_right[37] ,
    \ces_1_2_io_outs_right[36] ,
    \ces_1_2_io_outs_right[35] ,
    \ces_1_2_io_outs_right[34] ,
    \ces_1_2_io_outs_right[33] ,
    \ces_1_2_io_outs_right[32] ,
    \ces_1_2_io_outs_right[31] ,
    \ces_1_2_io_outs_right[30] ,
    \ces_1_2_io_outs_right[29] ,
    \ces_1_2_io_outs_right[28] ,
    \ces_1_2_io_outs_right[27] ,
    \ces_1_2_io_outs_right[26] ,
    \ces_1_2_io_outs_right[25] ,
    \ces_1_2_io_outs_right[24] ,
    \ces_1_2_io_outs_right[23] ,
    \ces_1_2_io_outs_right[22] ,
    \ces_1_2_io_outs_right[21] ,
    \ces_1_2_io_outs_right[20] ,
    \ces_1_2_io_outs_right[19] ,
    \ces_1_2_io_outs_right[18] ,
    \ces_1_2_io_outs_right[17] ,
    \ces_1_2_io_outs_right[16] ,
    \ces_1_2_io_outs_right[15] ,
    \ces_1_2_io_outs_right[14] ,
    \ces_1_2_io_outs_right[13] ,
    \ces_1_2_io_outs_right[12] ,
    \ces_1_2_io_outs_right[11] ,
    \ces_1_2_io_outs_right[10] ,
    \ces_1_2_io_outs_right[9] ,
    \ces_1_2_io_outs_right[8] ,
    \ces_1_2_io_outs_right[7] ,
    \ces_1_2_io_outs_right[6] ,
    \ces_1_2_io_outs_right[5] ,
    \ces_1_2_io_outs_right[4] ,
    \ces_1_2_io_outs_right[3] ,
    \ces_1_2_io_outs_right[2] ,
    \ces_1_2_io_outs_right[1] ,
    \ces_1_2_io_outs_right[0] }),
    .io_ins_up({\ces_0_3_io_outs_up[63] ,
    \ces_0_3_io_outs_up[62] ,
    \ces_0_3_io_outs_up[61] ,
    \ces_0_3_io_outs_up[60] ,
    \ces_0_3_io_outs_up[59] ,
    \ces_0_3_io_outs_up[58] ,
    \ces_0_3_io_outs_up[57] ,
    \ces_0_3_io_outs_up[56] ,
    \ces_0_3_io_outs_up[55] ,
    \ces_0_3_io_outs_up[54] ,
    \ces_0_3_io_outs_up[53] ,
    \ces_0_3_io_outs_up[52] ,
    \ces_0_3_io_outs_up[51] ,
    \ces_0_3_io_outs_up[50] ,
    \ces_0_3_io_outs_up[49] ,
    \ces_0_3_io_outs_up[48] ,
    \ces_0_3_io_outs_up[47] ,
    \ces_0_3_io_outs_up[46] ,
    \ces_0_3_io_outs_up[45] ,
    \ces_0_3_io_outs_up[44] ,
    \ces_0_3_io_outs_up[43] ,
    \ces_0_3_io_outs_up[42] ,
    \ces_0_3_io_outs_up[41] ,
    \ces_0_3_io_outs_up[40] ,
    \ces_0_3_io_outs_up[39] ,
    \ces_0_3_io_outs_up[38] ,
    \ces_0_3_io_outs_up[37] ,
    \ces_0_3_io_outs_up[36] ,
    \ces_0_3_io_outs_up[35] ,
    \ces_0_3_io_outs_up[34] ,
    \ces_0_3_io_outs_up[33] ,
    \ces_0_3_io_outs_up[32] ,
    \ces_0_3_io_outs_up[31] ,
    \ces_0_3_io_outs_up[30] ,
    \ces_0_3_io_outs_up[29] ,
    \ces_0_3_io_outs_up[28] ,
    \ces_0_3_io_outs_up[27] ,
    \ces_0_3_io_outs_up[26] ,
    \ces_0_3_io_outs_up[25] ,
    \ces_0_3_io_outs_up[24] ,
    \ces_0_3_io_outs_up[23] ,
    \ces_0_3_io_outs_up[22] ,
    \ces_0_3_io_outs_up[21] ,
    \ces_0_3_io_outs_up[20] ,
    \ces_0_3_io_outs_up[19] ,
    \ces_0_3_io_outs_up[18] ,
    \ces_0_3_io_outs_up[17] ,
    \ces_0_3_io_outs_up[16] ,
    \ces_0_3_io_outs_up[15] ,
    \ces_0_3_io_outs_up[14] ,
    \ces_0_3_io_outs_up[13] ,
    \ces_0_3_io_outs_up[12] ,
    \ces_0_3_io_outs_up[11] ,
    \ces_0_3_io_outs_up[10] ,
    \ces_0_3_io_outs_up[9] ,
    \ces_0_3_io_outs_up[8] ,
    \ces_0_3_io_outs_up[7] ,
    \ces_0_3_io_outs_up[6] ,
    \ces_0_3_io_outs_up[5] ,
    \ces_0_3_io_outs_up[4] ,
    \ces_0_3_io_outs_up[3] ,
    \ces_0_3_io_outs_up[2] ,
    \ces_0_3_io_outs_up[1] ,
    \ces_0_3_io_outs_up[0] }),
    .io_outs_down({\ces_0_3_io_ins_down[63] ,
    \ces_0_3_io_ins_down[62] ,
    \ces_0_3_io_ins_down[61] ,
    \ces_0_3_io_ins_down[60] ,
    \ces_0_3_io_ins_down[59] ,
    \ces_0_3_io_ins_down[58] ,
    \ces_0_3_io_ins_down[57] ,
    \ces_0_3_io_ins_down[56] ,
    \ces_0_3_io_ins_down[55] ,
    \ces_0_3_io_ins_down[54] ,
    \ces_0_3_io_ins_down[53] ,
    \ces_0_3_io_ins_down[52] ,
    \ces_0_3_io_ins_down[51] ,
    \ces_0_3_io_ins_down[50] ,
    \ces_0_3_io_ins_down[49] ,
    \ces_0_3_io_ins_down[48] ,
    \ces_0_3_io_ins_down[47] ,
    \ces_0_3_io_ins_down[46] ,
    \ces_0_3_io_ins_down[45] ,
    \ces_0_3_io_ins_down[44] ,
    \ces_0_3_io_ins_down[43] ,
    \ces_0_3_io_ins_down[42] ,
    \ces_0_3_io_ins_down[41] ,
    \ces_0_3_io_ins_down[40] ,
    \ces_0_3_io_ins_down[39] ,
    \ces_0_3_io_ins_down[38] ,
    \ces_0_3_io_ins_down[37] ,
    \ces_0_3_io_ins_down[36] ,
    \ces_0_3_io_ins_down[35] ,
    \ces_0_3_io_ins_down[34] ,
    \ces_0_3_io_ins_down[33] ,
    \ces_0_3_io_ins_down[32] ,
    \ces_0_3_io_ins_down[31] ,
    \ces_0_3_io_ins_down[30] ,
    \ces_0_3_io_ins_down[29] ,
    \ces_0_3_io_ins_down[28] ,
    \ces_0_3_io_ins_down[27] ,
    \ces_0_3_io_ins_down[26] ,
    \ces_0_3_io_ins_down[25] ,
    \ces_0_3_io_ins_down[24] ,
    \ces_0_3_io_ins_down[23] ,
    \ces_0_3_io_ins_down[22] ,
    \ces_0_3_io_ins_down[21] ,
    \ces_0_3_io_ins_down[20] ,
    \ces_0_3_io_ins_down[19] ,
    \ces_0_3_io_ins_down[18] ,
    \ces_0_3_io_ins_down[17] ,
    \ces_0_3_io_ins_down[16] ,
    \ces_0_3_io_ins_down[15] ,
    \ces_0_3_io_ins_down[14] ,
    \ces_0_3_io_ins_down[13] ,
    \ces_0_3_io_ins_down[12] ,
    \ces_0_3_io_ins_down[11] ,
    \ces_0_3_io_ins_down[10] ,
    \ces_0_3_io_ins_down[9] ,
    \ces_0_3_io_ins_down[8] ,
    \ces_0_3_io_ins_down[7] ,
    \ces_0_3_io_ins_down[6] ,
    \ces_0_3_io_ins_down[5] ,
    \ces_0_3_io_ins_down[4] ,
    \ces_0_3_io_ins_down[3] ,
    \ces_0_3_io_ins_down[2] ,
    \ces_0_3_io_ins_down[1] ,
    \ces_0_3_io_ins_down[0] }),
    .io_outs_left({\ces_1_2_io_ins_left[63] ,
    \ces_1_2_io_ins_left[62] ,
    \ces_1_2_io_ins_left[61] ,
    \ces_1_2_io_ins_left[60] ,
    \ces_1_2_io_ins_left[59] ,
    \ces_1_2_io_ins_left[58] ,
    \ces_1_2_io_ins_left[57] ,
    \ces_1_2_io_ins_left[56] ,
    \ces_1_2_io_ins_left[55] ,
    \ces_1_2_io_ins_left[54] ,
    \ces_1_2_io_ins_left[53] ,
    \ces_1_2_io_ins_left[52] ,
    \ces_1_2_io_ins_left[51] ,
    \ces_1_2_io_ins_left[50] ,
    \ces_1_2_io_ins_left[49] ,
    \ces_1_2_io_ins_left[48] ,
    \ces_1_2_io_ins_left[47] ,
    \ces_1_2_io_ins_left[46] ,
    \ces_1_2_io_ins_left[45] ,
    \ces_1_2_io_ins_left[44] ,
    \ces_1_2_io_ins_left[43] ,
    \ces_1_2_io_ins_left[42] ,
    \ces_1_2_io_ins_left[41] ,
    \ces_1_2_io_ins_left[40] ,
    \ces_1_2_io_ins_left[39] ,
    \ces_1_2_io_ins_left[38] ,
    \ces_1_2_io_ins_left[37] ,
    \ces_1_2_io_ins_left[36] ,
    \ces_1_2_io_ins_left[35] ,
    \ces_1_2_io_ins_left[34] ,
    \ces_1_2_io_ins_left[33] ,
    \ces_1_2_io_ins_left[32] ,
    \ces_1_2_io_ins_left[31] ,
    \ces_1_2_io_ins_left[30] ,
    \ces_1_2_io_ins_left[29] ,
    \ces_1_2_io_ins_left[28] ,
    \ces_1_2_io_ins_left[27] ,
    \ces_1_2_io_ins_left[26] ,
    \ces_1_2_io_ins_left[25] ,
    \ces_1_2_io_ins_left[24] ,
    \ces_1_2_io_ins_left[23] ,
    \ces_1_2_io_ins_left[22] ,
    \ces_1_2_io_ins_left[21] ,
    \ces_1_2_io_ins_left[20] ,
    \ces_1_2_io_ins_left[19] ,
    \ces_1_2_io_ins_left[18] ,
    \ces_1_2_io_ins_left[17] ,
    \ces_1_2_io_ins_left[16] ,
    \ces_1_2_io_ins_left[15] ,
    \ces_1_2_io_ins_left[14] ,
    \ces_1_2_io_ins_left[13] ,
    \ces_1_2_io_ins_left[12] ,
    \ces_1_2_io_ins_left[11] ,
    \ces_1_2_io_ins_left[10] ,
    \ces_1_2_io_ins_left[9] ,
    \ces_1_2_io_ins_left[8] ,
    \ces_1_2_io_ins_left[7] ,
    \ces_1_2_io_ins_left[6] ,
    \ces_1_2_io_ins_left[5] ,
    \ces_1_2_io_ins_left[4] ,
    \ces_1_2_io_ins_left[3] ,
    \ces_1_2_io_ins_left[2] ,
    \ces_1_2_io_ins_left[1] ,
    \ces_1_2_io_ins_left[0] }),
    .io_outs_right({\ces_1_3_io_outs_right[63] ,
    \ces_1_3_io_outs_right[62] ,
    \ces_1_3_io_outs_right[61] ,
    \ces_1_3_io_outs_right[60] ,
    \ces_1_3_io_outs_right[59] ,
    \ces_1_3_io_outs_right[58] ,
    \ces_1_3_io_outs_right[57] ,
    \ces_1_3_io_outs_right[56] ,
    \ces_1_3_io_outs_right[55] ,
    \ces_1_3_io_outs_right[54] ,
    \ces_1_3_io_outs_right[53] ,
    \ces_1_3_io_outs_right[52] ,
    \ces_1_3_io_outs_right[51] ,
    \ces_1_3_io_outs_right[50] ,
    \ces_1_3_io_outs_right[49] ,
    \ces_1_3_io_outs_right[48] ,
    \ces_1_3_io_outs_right[47] ,
    \ces_1_3_io_outs_right[46] ,
    \ces_1_3_io_outs_right[45] ,
    \ces_1_3_io_outs_right[44] ,
    \ces_1_3_io_outs_right[43] ,
    \ces_1_3_io_outs_right[42] ,
    \ces_1_3_io_outs_right[41] ,
    \ces_1_3_io_outs_right[40] ,
    \ces_1_3_io_outs_right[39] ,
    \ces_1_3_io_outs_right[38] ,
    \ces_1_3_io_outs_right[37] ,
    \ces_1_3_io_outs_right[36] ,
    \ces_1_3_io_outs_right[35] ,
    \ces_1_3_io_outs_right[34] ,
    \ces_1_3_io_outs_right[33] ,
    \ces_1_3_io_outs_right[32] ,
    \ces_1_3_io_outs_right[31] ,
    \ces_1_3_io_outs_right[30] ,
    \ces_1_3_io_outs_right[29] ,
    \ces_1_3_io_outs_right[28] ,
    \ces_1_3_io_outs_right[27] ,
    \ces_1_3_io_outs_right[26] ,
    \ces_1_3_io_outs_right[25] ,
    \ces_1_3_io_outs_right[24] ,
    \ces_1_3_io_outs_right[23] ,
    \ces_1_3_io_outs_right[22] ,
    \ces_1_3_io_outs_right[21] ,
    \ces_1_3_io_outs_right[20] ,
    \ces_1_3_io_outs_right[19] ,
    \ces_1_3_io_outs_right[18] ,
    \ces_1_3_io_outs_right[17] ,
    \ces_1_3_io_outs_right[16] ,
    \ces_1_3_io_outs_right[15] ,
    \ces_1_3_io_outs_right[14] ,
    \ces_1_3_io_outs_right[13] ,
    \ces_1_3_io_outs_right[12] ,
    \ces_1_3_io_outs_right[11] ,
    \ces_1_3_io_outs_right[10] ,
    \ces_1_3_io_outs_right[9] ,
    \ces_1_3_io_outs_right[8] ,
    \ces_1_3_io_outs_right[7] ,
    \ces_1_3_io_outs_right[6] ,
    \ces_1_3_io_outs_right[5] ,
    \ces_1_3_io_outs_right[4] ,
    \ces_1_3_io_outs_right[3] ,
    \ces_1_3_io_outs_right[2] ,
    \ces_1_3_io_outs_right[1] ,
    \ces_1_3_io_outs_right[0] }),
    .io_outs_up({\ces_1_3_io_outs_up[63] ,
    \ces_1_3_io_outs_up[62] ,
    \ces_1_3_io_outs_up[61] ,
    \ces_1_3_io_outs_up[60] ,
    \ces_1_3_io_outs_up[59] ,
    \ces_1_3_io_outs_up[58] ,
    \ces_1_3_io_outs_up[57] ,
    \ces_1_3_io_outs_up[56] ,
    \ces_1_3_io_outs_up[55] ,
    \ces_1_3_io_outs_up[54] ,
    \ces_1_3_io_outs_up[53] ,
    \ces_1_3_io_outs_up[52] ,
    \ces_1_3_io_outs_up[51] ,
    \ces_1_3_io_outs_up[50] ,
    \ces_1_3_io_outs_up[49] ,
    \ces_1_3_io_outs_up[48] ,
    \ces_1_3_io_outs_up[47] ,
    \ces_1_3_io_outs_up[46] ,
    \ces_1_3_io_outs_up[45] ,
    \ces_1_3_io_outs_up[44] ,
    \ces_1_3_io_outs_up[43] ,
    \ces_1_3_io_outs_up[42] ,
    \ces_1_3_io_outs_up[41] ,
    \ces_1_3_io_outs_up[40] ,
    \ces_1_3_io_outs_up[39] ,
    \ces_1_3_io_outs_up[38] ,
    \ces_1_3_io_outs_up[37] ,
    \ces_1_3_io_outs_up[36] ,
    \ces_1_3_io_outs_up[35] ,
    \ces_1_3_io_outs_up[34] ,
    \ces_1_3_io_outs_up[33] ,
    \ces_1_3_io_outs_up[32] ,
    \ces_1_3_io_outs_up[31] ,
    \ces_1_3_io_outs_up[30] ,
    \ces_1_3_io_outs_up[29] ,
    \ces_1_3_io_outs_up[28] ,
    \ces_1_3_io_outs_up[27] ,
    \ces_1_3_io_outs_up[26] ,
    \ces_1_3_io_outs_up[25] ,
    \ces_1_3_io_outs_up[24] ,
    \ces_1_3_io_outs_up[23] ,
    \ces_1_3_io_outs_up[22] ,
    \ces_1_3_io_outs_up[21] ,
    \ces_1_3_io_outs_up[20] ,
    \ces_1_3_io_outs_up[19] ,
    \ces_1_3_io_outs_up[18] ,
    \ces_1_3_io_outs_up[17] ,
    \ces_1_3_io_outs_up[16] ,
    \ces_1_3_io_outs_up[15] ,
    \ces_1_3_io_outs_up[14] ,
    \ces_1_3_io_outs_up[13] ,
    \ces_1_3_io_outs_up[12] ,
    \ces_1_3_io_outs_up[11] ,
    \ces_1_3_io_outs_up[10] ,
    \ces_1_3_io_outs_up[9] ,
    \ces_1_3_io_outs_up[8] ,
    \ces_1_3_io_outs_up[7] ,
    \ces_1_3_io_outs_up[6] ,
    \ces_1_3_io_outs_up[5] ,
    \ces_1_3_io_outs_up[4] ,
    \ces_1_3_io_outs_up[3] ,
    \ces_1_3_io_outs_up[2] ,
    \ces_1_3_io_outs_up[1] ,
    \ces_1_3_io_outs_up[0] }));
 Element ces_1_4 (.clock(clknet_3_2_0_clock),
    .io_lsbIns_1(ces_1_3_io_lsbOuts_1),
    .io_lsbIns_2(ces_1_3_io_lsbOuts_2),
    .io_lsbIns_3(ces_1_3_io_lsbOuts_3),
    .io_lsbIns_4(ces_1_3_io_lsbOuts_4),
    .io_lsbIns_5(ces_1_3_io_lsbOuts_5),
    .io_lsbIns_6(ces_1_3_io_lsbOuts_6),
    .io_lsbIns_7(ces_1_3_io_lsbOuts_7),
    .io_lsbOuts_0(ces_1_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_4_io_lsbOuts_7),
    .io_ins_down({\ces_1_4_io_ins_down[63] ,
    \ces_1_4_io_ins_down[62] ,
    \ces_1_4_io_ins_down[61] ,
    \ces_1_4_io_ins_down[60] ,
    \ces_1_4_io_ins_down[59] ,
    \ces_1_4_io_ins_down[58] ,
    \ces_1_4_io_ins_down[57] ,
    \ces_1_4_io_ins_down[56] ,
    \ces_1_4_io_ins_down[55] ,
    \ces_1_4_io_ins_down[54] ,
    \ces_1_4_io_ins_down[53] ,
    \ces_1_4_io_ins_down[52] ,
    \ces_1_4_io_ins_down[51] ,
    \ces_1_4_io_ins_down[50] ,
    \ces_1_4_io_ins_down[49] ,
    \ces_1_4_io_ins_down[48] ,
    \ces_1_4_io_ins_down[47] ,
    \ces_1_4_io_ins_down[46] ,
    \ces_1_4_io_ins_down[45] ,
    \ces_1_4_io_ins_down[44] ,
    \ces_1_4_io_ins_down[43] ,
    \ces_1_4_io_ins_down[42] ,
    \ces_1_4_io_ins_down[41] ,
    \ces_1_4_io_ins_down[40] ,
    \ces_1_4_io_ins_down[39] ,
    \ces_1_4_io_ins_down[38] ,
    \ces_1_4_io_ins_down[37] ,
    \ces_1_4_io_ins_down[36] ,
    \ces_1_4_io_ins_down[35] ,
    \ces_1_4_io_ins_down[34] ,
    \ces_1_4_io_ins_down[33] ,
    \ces_1_4_io_ins_down[32] ,
    \ces_1_4_io_ins_down[31] ,
    \ces_1_4_io_ins_down[30] ,
    \ces_1_4_io_ins_down[29] ,
    \ces_1_4_io_ins_down[28] ,
    \ces_1_4_io_ins_down[27] ,
    \ces_1_4_io_ins_down[26] ,
    \ces_1_4_io_ins_down[25] ,
    \ces_1_4_io_ins_down[24] ,
    \ces_1_4_io_ins_down[23] ,
    \ces_1_4_io_ins_down[22] ,
    \ces_1_4_io_ins_down[21] ,
    \ces_1_4_io_ins_down[20] ,
    \ces_1_4_io_ins_down[19] ,
    \ces_1_4_io_ins_down[18] ,
    \ces_1_4_io_ins_down[17] ,
    \ces_1_4_io_ins_down[16] ,
    \ces_1_4_io_ins_down[15] ,
    \ces_1_4_io_ins_down[14] ,
    \ces_1_4_io_ins_down[13] ,
    \ces_1_4_io_ins_down[12] ,
    \ces_1_4_io_ins_down[11] ,
    \ces_1_4_io_ins_down[10] ,
    \ces_1_4_io_ins_down[9] ,
    \ces_1_4_io_ins_down[8] ,
    \ces_1_4_io_ins_down[7] ,
    \ces_1_4_io_ins_down[6] ,
    \ces_1_4_io_ins_down[5] ,
    \ces_1_4_io_ins_down[4] ,
    \ces_1_4_io_ins_down[3] ,
    \ces_1_4_io_ins_down[2] ,
    \ces_1_4_io_ins_down[1] ,
    \ces_1_4_io_ins_down[0] }),
    .io_ins_left({\ces_1_4_io_ins_left[63] ,
    \ces_1_4_io_ins_left[62] ,
    \ces_1_4_io_ins_left[61] ,
    \ces_1_4_io_ins_left[60] ,
    \ces_1_4_io_ins_left[59] ,
    \ces_1_4_io_ins_left[58] ,
    \ces_1_4_io_ins_left[57] ,
    \ces_1_4_io_ins_left[56] ,
    \ces_1_4_io_ins_left[55] ,
    \ces_1_4_io_ins_left[54] ,
    \ces_1_4_io_ins_left[53] ,
    \ces_1_4_io_ins_left[52] ,
    \ces_1_4_io_ins_left[51] ,
    \ces_1_4_io_ins_left[50] ,
    \ces_1_4_io_ins_left[49] ,
    \ces_1_4_io_ins_left[48] ,
    \ces_1_4_io_ins_left[47] ,
    \ces_1_4_io_ins_left[46] ,
    \ces_1_4_io_ins_left[45] ,
    \ces_1_4_io_ins_left[44] ,
    \ces_1_4_io_ins_left[43] ,
    \ces_1_4_io_ins_left[42] ,
    \ces_1_4_io_ins_left[41] ,
    \ces_1_4_io_ins_left[40] ,
    \ces_1_4_io_ins_left[39] ,
    \ces_1_4_io_ins_left[38] ,
    \ces_1_4_io_ins_left[37] ,
    \ces_1_4_io_ins_left[36] ,
    \ces_1_4_io_ins_left[35] ,
    \ces_1_4_io_ins_left[34] ,
    \ces_1_4_io_ins_left[33] ,
    \ces_1_4_io_ins_left[32] ,
    \ces_1_4_io_ins_left[31] ,
    \ces_1_4_io_ins_left[30] ,
    \ces_1_4_io_ins_left[29] ,
    \ces_1_4_io_ins_left[28] ,
    \ces_1_4_io_ins_left[27] ,
    \ces_1_4_io_ins_left[26] ,
    \ces_1_4_io_ins_left[25] ,
    \ces_1_4_io_ins_left[24] ,
    \ces_1_4_io_ins_left[23] ,
    \ces_1_4_io_ins_left[22] ,
    \ces_1_4_io_ins_left[21] ,
    \ces_1_4_io_ins_left[20] ,
    \ces_1_4_io_ins_left[19] ,
    \ces_1_4_io_ins_left[18] ,
    \ces_1_4_io_ins_left[17] ,
    \ces_1_4_io_ins_left[16] ,
    \ces_1_4_io_ins_left[15] ,
    \ces_1_4_io_ins_left[14] ,
    \ces_1_4_io_ins_left[13] ,
    \ces_1_4_io_ins_left[12] ,
    \ces_1_4_io_ins_left[11] ,
    \ces_1_4_io_ins_left[10] ,
    \ces_1_4_io_ins_left[9] ,
    \ces_1_4_io_ins_left[8] ,
    \ces_1_4_io_ins_left[7] ,
    \ces_1_4_io_ins_left[6] ,
    \ces_1_4_io_ins_left[5] ,
    \ces_1_4_io_ins_left[4] ,
    \ces_1_4_io_ins_left[3] ,
    \ces_1_4_io_ins_left[2] ,
    \ces_1_4_io_ins_left[1] ,
    \ces_1_4_io_ins_left[0] }),
    .io_ins_right({\ces_1_3_io_outs_right[63] ,
    \ces_1_3_io_outs_right[62] ,
    \ces_1_3_io_outs_right[61] ,
    \ces_1_3_io_outs_right[60] ,
    \ces_1_3_io_outs_right[59] ,
    \ces_1_3_io_outs_right[58] ,
    \ces_1_3_io_outs_right[57] ,
    \ces_1_3_io_outs_right[56] ,
    \ces_1_3_io_outs_right[55] ,
    \ces_1_3_io_outs_right[54] ,
    \ces_1_3_io_outs_right[53] ,
    \ces_1_3_io_outs_right[52] ,
    \ces_1_3_io_outs_right[51] ,
    \ces_1_3_io_outs_right[50] ,
    \ces_1_3_io_outs_right[49] ,
    \ces_1_3_io_outs_right[48] ,
    \ces_1_3_io_outs_right[47] ,
    \ces_1_3_io_outs_right[46] ,
    \ces_1_3_io_outs_right[45] ,
    \ces_1_3_io_outs_right[44] ,
    \ces_1_3_io_outs_right[43] ,
    \ces_1_3_io_outs_right[42] ,
    \ces_1_3_io_outs_right[41] ,
    \ces_1_3_io_outs_right[40] ,
    \ces_1_3_io_outs_right[39] ,
    \ces_1_3_io_outs_right[38] ,
    \ces_1_3_io_outs_right[37] ,
    \ces_1_3_io_outs_right[36] ,
    \ces_1_3_io_outs_right[35] ,
    \ces_1_3_io_outs_right[34] ,
    \ces_1_3_io_outs_right[33] ,
    \ces_1_3_io_outs_right[32] ,
    \ces_1_3_io_outs_right[31] ,
    \ces_1_3_io_outs_right[30] ,
    \ces_1_3_io_outs_right[29] ,
    \ces_1_3_io_outs_right[28] ,
    \ces_1_3_io_outs_right[27] ,
    \ces_1_3_io_outs_right[26] ,
    \ces_1_3_io_outs_right[25] ,
    \ces_1_3_io_outs_right[24] ,
    \ces_1_3_io_outs_right[23] ,
    \ces_1_3_io_outs_right[22] ,
    \ces_1_3_io_outs_right[21] ,
    \ces_1_3_io_outs_right[20] ,
    \ces_1_3_io_outs_right[19] ,
    \ces_1_3_io_outs_right[18] ,
    \ces_1_3_io_outs_right[17] ,
    \ces_1_3_io_outs_right[16] ,
    \ces_1_3_io_outs_right[15] ,
    \ces_1_3_io_outs_right[14] ,
    \ces_1_3_io_outs_right[13] ,
    \ces_1_3_io_outs_right[12] ,
    \ces_1_3_io_outs_right[11] ,
    \ces_1_3_io_outs_right[10] ,
    \ces_1_3_io_outs_right[9] ,
    \ces_1_3_io_outs_right[8] ,
    \ces_1_3_io_outs_right[7] ,
    \ces_1_3_io_outs_right[6] ,
    \ces_1_3_io_outs_right[5] ,
    \ces_1_3_io_outs_right[4] ,
    \ces_1_3_io_outs_right[3] ,
    \ces_1_3_io_outs_right[2] ,
    \ces_1_3_io_outs_right[1] ,
    \ces_1_3_io_outs_right[0] }),
    .io_ins_up({\ces_0_4_io_outs_up[63] ,
    \ces_0_4_io_outs_up[62] ,
    \ces_0_4_io_outs_up[61] ,
    \ces_0_4_io_outs_up[60] ,
    \ces_0_4_io_outs_up[59] ,
    \ces_0_4_io_outs_up[58] ,
    \ces_0_4_io_outs_up[57] ,
    \ces_0_4_io_outs_up[56] ,
    \ces_0_4_io_outs_up[55] ,
    \ces_0_4_io_outs_up[54] ,
    \ces_0_4_io_outs_up[53] ,
    \ces_0_4_io_outs_up[52] ,
    \ces_0_4_io_outs_up[51] ,
    \ces_0_4_io_outs_up[50] ,
    \ces_0_4_io_outs_up[49] ,
    \ces_0_4_io_outs_up[48] ,
    \ces_0_4_io_outs_up[47] ,
    \ces_0_4_io_outs_up[46] ,
    \ces_0_4_io_outs_up[45] ,
    \ces_0_4_io_outs_up[44] ,
    \ces_0_4_io_outs_up[43] ,
    \ces_0_4_io_outs_up[42] ,
    \ces_0_4_io_outs_up[41] ,
    \ces_0_4_io_outs_up[40] ,
    \ces_0_4_io_outs_up[39] ,
    \ces_0_4_io_outs_up[38] ,
    \ces_0_4_io_outs_up[37] ,
    \ces_0_4_io_outs_up[36] ,
    \ces_0_4_io_outs_up[35] ,
    \ces_0_4_io_outs_up[34] ,
    \ces_0_4_io_outs_up[33] ,
    \ces_0_4_io_outs_up[32] ,
    \ces_0_4_io_outs_up[31] ,
    \ces_0_4_io_outs_up[30] ,
    \ces_0_4_io_outs_up[29] ,
    \ces_0_4_io_outs_up[28] ,
    \ces_0_4_io_outs_up[27] ,
    \ces_0_4_io_outs_up[26] ,
    \ces_0_4_io_outs_up[25] ,
    \ces_0_4_io_outs_up[24] ,
    \ces_0_4_io_outs_up[23] ,
    \ces_0_4_io_outs_up[22] ,
    \ces_0_4_io_outs_up[21] ,
    \ces_0_4_io_outs_up[20] ,
    \ces_0_4_io_outs_up[19] ,
    \ces_0_4_io_outs_up[18] ,
    \ces_0_4_io_outs_up[17] ,
    \ces_0_4_io_outs_up[16] ,
    \ces_0_4_io_outs_up[15] ,
    \ces_0_4_io_outs_up[14] ,
    \ces_0_4_io_outs_up[13] ,
    \ces_0_4_io_outs_up[12] ,
    \ces_0_4_io_outs_up[11] ,
    \ces_0_4_io_outs_up[10] ,
    \ces_0_4_io_outs_up[9] ,
    \ces_0_4_io_outs_up[8] ,
    \ces_0_4_io_outs_up[7] ,
    \ces_0_4_io_outs_up[6] ,
    \ces_0_4_io_outs_up[5] ,
    \ces_0_4_io_outs_up[4] ,
    \ces_0_4_io_outs_up[3] ,
    \ces_0_4_io_outs_up[2] ,
    \ces_0_4_io_outs_up[1] ,
    \ces_0_4_io_outs_up[0] }),
    .io_outs_down({\ces_0_4_io_ins_down[63] ,
    \ces_0_4_io_ins_down[62] ,
    \ces_0_4_io_ins_down[61] ,
    \ces_0_4_io_ins_down[60] ,
    \ces_0_4_io_ins_down[59] ,
    \ces_0_4_io_ins_down[58] ,
    \ces_0_4_io_ins_down[57] ,
    \ces_0_4_io_ins_down[56] ,
    \ces_0_4_io_ins_down[55] ,
    \ces_0_4_io_ins_down[54] ,
    \ces_0_4_io_ins_down[53] ,
    \ces_0_4_io_ins_down[52] ,
    \ces_0_4_io_ins_down[51] ,
    \ces_0_4_io_ins_down[50] ,
    \ces_0_4_io_ins_down[49] ,
    \ces_0_4_io_ins_down[48] ,
    \ces_0_4_io_ins_down[47] ,
    \ces_0_4_io_ins_down[46] ,
    \ces_0_4_io_ins_down[45] ,
    \ces_0_4_io_ins_down[44] ,
    \ces_0_4_io_ins_down[43] ,
    \ces_0_4_io_ins_down[42] ,
    \ces_0_4_io_ins_down[41] ,
    \ces_0_4_io_ins_down[40] ,
    \ces_0_4_io_ins_down[39] ,
    \ces_0_4_io_ins_down[38] ,
    \ces_0_4_io_ins_down[37] ,
    \ces_0_4_io_ins_down[36] ,
    \ces_0_4_io_ins_down[35] ,
    \ces_0_4_io_ins_down[34] ,
    \ces_0_4_io_ins_down[33] ,
    \ces_0_4_io_ins_down[32] ,
    \ces_0_4_io_ins_down[31] ,
    \ces_0_4_io_ins_down[30] ,
    \ces_0_4_io_ins_down[29] ,
    \ces_0_4_io_ins_down[28] ,
    \ces_0_4_io_ins_down[27] ,
    \ces_0_4_io_ins_down[26] ,
    \ces_0_4_io_ins_down[25] ,
    \ces_0_4_io_ins_down[24] ,
    \ces_0_4_io_ins_down[23] ,
    \ces_0_4_io_ins_down[22] ,
    \ces_0_4_io_ins_down[21] ,
    \ces_0_4_io_ins_down[20] ,
    \ces_0_4_io_ins_down[19] ,
    \ces_0_4_io_ins_down[18] ,
    \ces_0_4_io_ins_down[17] ,
    \ces_0_4_io_ins_down[16] ,
    \ces_0_4_io_ins_down[15] ,
    \ces_0_4_io_ins_down[14] ,
    \ces_0_4_io_ins_down[13] ,
    \ces_0_4_io_ins_down[12] ,
    \ces_0_4_io_ins_down[11] ,
    \ces_0_4_io_ins_down[10] ,
    \ces_0_4_io_ins_down[9] ,
    \ces_0_4_io_ins_down[8] ,
    \ces_0_4_io_ins_down[7] ,
    \ces_0_4_io_ins_down[6] ,
    \ces_0_4_io_ins_down[5] ,
    \ces_0_4_io_ins_down[4] ,
    \ces_0_4_io_ins_down[3] ,
    \ces_0_4_io_ins_down[2] ,
    \ces_0_4_io_ins_down[1] ,
    \ces_0_4_io_ins_down[0] }),
    .io_outs_left({\ces_1_3_io_ins_left[63] ,
    \ces_1_3_io_ins_left[62] ,
    \ces_1_3_io_ins_left[61] ,
    \ces_1_3_io_ins_left[60] ,
    \ces_1_3_io_ins_left[59] ,
    \ces_1_3_io_ins_left[58] ,
    \ces_1_3_io_ins_left[57] ,
    \ces_1_3_io_ins_left[56] ,
    \ces_1_3_io_ins_left[55] ,
    \ces_1_3_io_ins_left[54] ,
    \ces_1_3_io_ins_left[53] ,
    \ces_1_3_io_ins_left[52] ,
    \ces_1_3_io_ins_left[51] ,
    \ces_1_3_io_ins_left[50] ,
    \ces_1_3_io_ins_left[49] ,
    \ces_1_3_io_ins_left[48] ,
    \ces_1_3_io_ins_left[47] ,
    \ces_1_3_io_ins_left[46] ,
    \ces_1_3_io_ins_left[45] ,
    \ces_1_3_io_ins_left[44] ,
    \ces_1_3_io_ins_left[43] ,
    \ces_1_3_io_ins_left[42] ,
    \ces_1_3_io_ins_left[41] ,
    \ces_1_3_io_ins_left[40] ,
    \ces_1_3_io_ins_left[39] ,
    \ces_1_3_io_ins_left[38] ,
    \ces_1_3_io_ins_left[37] ,
    \ces_1_3_io_ins_left[36] ,
    \ces_1_3_io_ins_left[35] ,
    \ces_1_3_io_ins_left[34] ,
    \ces_1_3_io_ins_left[33] ,
    \ces_1_3_io_ins_left[32] ,
    \ces_1_3_io_ins_left[31] ,
    \ces_1_3_io_ins_left[30] ,
    \ces_1_3_io_ins_left[29] ,
    \ces_1_3_io_ins_left[28] ,
    \ces_1_3_io_ins_left[27] ,
    \ces_1_3_io_ins_left[26] ,
    \ces_1_3_io_ins_left[25] ,
    \ces_1_3_io_ins_left[24] ,
    \ces_1_3_io_ins_left[23] ,
    \ces_1_3_io_ins_left[22] ,
    \ces_1_3_io_ins_left[21] ,
    \ces_1_3_io_ins_left[20] ,
    \ces_1_3_io_ins_left[19] ,
    \ces_1_3_io_ins_left[18] ,
    \ces_1_3_io_ins_left[17] ,
    \ces_1_3_io_ins_left[16] ,
    \ces_1_3_io_ins_left[15] ,
    \ces_1_3_io_ins_left[14] ,
    \ces_1_3_io_ins_left[13] ,
    \ces_1_3_io_ins_left[12] ,
    \ces_1_3_io_ins_left[11] ,
    \ces_1_3_io_ins_left[10] ,
    \ces_1_3_io_ins_left[9] ,
    \ces_1_3_io_ins_left[8] ,
    \ces_1_3_io_ins_left[7] ,
    \ces_1_3_io_ins_left[6] ,
    \ces_1_3_io_ins_left[5] ,
    \ces_1_3_io_ins_left[4] ,
    \ces_1_3_io_ins_left[3] ,
    \ces_1_3_io_ins_left[2] ,
    \ces_1_3_io_ins_left[1] ,
    \ces_1_3_io_ins_left[0] }),
    .io_outs_right({\ces_1_4_io_outs_right[63] ,
    \ces_1_4_io_outs_right[62] ,
    \ces_1_4_io_outs_right[61] ,
    \ces_1_4_io_outs_right[60] ,
    \ces_1_4_io_outs_right[59] ,
    \ces_1_4_io_outs_right[58] ,
    \ces_1_4_io_outs_right[57] ,
    \ces_1_4_io_outs_right[56] ,
    \ces_1_4_io_outs_right[55] ,
    \ces_1_4_io_outs_right[54] ,
    \ces_1_4_io_outs_right[53] ,
    \ces_1_4_io_outs_right[52] ,
    \ces_1_4_io_outs_right[51] ,
    \ces_1_4_io_outs_right[50] ,
    \ces_1_4_io_outs_right[49] ,
    \ces_1_4_io_outs_right[48] ,
    \ces_1_4_io_outs_right[47] ,
    \ces_1_4_io_outs_right[46] ,
    \ces_1_4_io_outs_right[45] ,
    \ces_1_4_io_outs_right[44] ,
    \ces_1_4_io_outs_right[43] ,
    \ces_1_4_io_outs_right[42] ,
    \ces_1_4_io_outs_right[41] ,
    \ces_1_4_io_outs_right[40] ,
    \ces_1_4_io_outs_right[39] ,
    \ces_1_4_io_outs_right[38] ,
    \ces_1_4_io_outs_right[37] ,
    \ces_1_4_io_outs_right[36] ,
    \ces_1_4_io_outs_right[35] ,
    \ces_1_4_io_outs_right[34] ,
    \ces_1_4_io_outs_right[33] ,
    \ces_1_4_io_outs_right[32] ,
    \ces_1_4_io_outs_right[31] ,
    \ces_1_4_io_outs_right[30] ,
    \ces_1_4_io_outs_right[29] ,
    \ces_1_4_io_outs_right[28] ,
    \ces_1_4_io_outs_right[27] ,
    \ces_1_4_io_outs_right[26] ,
    \ces_1_4_io_outs_right[25] ,
    \ces_1_4_io_outs_right[24] ,
    \ces_1_4_io_outs_right[23] ,
    \ces_1_4_io_outs_right[22] ,
    \ces_1_4_io_outs_right[21] ,
    \ces_1_4_io_outs_right[20] ,
    \ces_1_4_io_outs_right[19] ,
    \ces_1_4_io_outs_right[18] ,
    \ces_1_4_io_outs_right[17] ,
    \ces_1_4_io_outs_right[16] ,
    \ces_1_4_io_outs_right[15] ,
    \ces_1_4_io_outs_right[14] ,
    \ces_1_4_io_outs_right[13] ,
    \ces_1_4_io_outs_right[12] ,
    \ces_1_4_io_outs_right[11] ,
    \ces_1_4_io_outs_right[10] ,
    \ces_1_4_io_outs_right[9] ,
    \ces_1_4_io_outs_right[8] ,
    \ces_1_4_io_outs_right[7] ,
    \ces_1_4_io_outs_right[6] ,
    \ces_1_4_io_outs_right[5] ,
    \ces_1_4_io_outs_right[4] ,
    \ces_1_4_io_outs_right[3] ,
    \ces_1_4_io_outs_right[2] ,
    \ces_1_4_io_outs_right[1] ,
    \ces_1_4_io_outs_right[0] }),
    .io_outs_up({\ces_1_4_io_outs_up[63] ,
    \ces_1_4_io_outs_up[62] ,
    \ces_1_4_io_outs_up[61] ,
    \ces_1_4_io_outs_up[60] ,
    \ces_1_4_io_outs_up[59] ,
    \ces_1_4_io_outs_up[58] ,
    \ces_1_4_io_outs_up[57] ,
    \ces_1_4_io_outs_up[56] ,
    \ces_1_4_io_outs_up[55] ,
    \ces_1_4_io_outs_up[54] ,
    \ces_1_4_io_outs_up[53] ,
    \ces_1_4_io_outs_up[52] ,
    \ces_1_4_io_outs_up[51] ,
    \ces_1_4_io_outs_up[50] ,
    \ces_1_4_io_outs_up[49] ,
    \ces_1_4_io_outs_up[48] ,
    \ces_1_4_io_outs_up[47] ,
    \ces_1_4_io_outs_up[46] ,
    \ces_1_4_io_outs_up[45] ,
    \ces_1_4_io_outs_up[44] ,
    \ces_1_4_io_outs_up[43] ,
    \ces_1_4_io_outs_up[42] ,
    \ces_1_4_io_outs_up[41] ,
    \ces_1_4_io_outs_up[40] ,
    \ces_1_4_io_outs_up[39] ,
    \ces_1_4_io_outs_up[38] ,
    \ces_1_4_io_outs_up[37] ,
    \ces_1_4_io_outs_up[36] ,
    \ces_1_4_io_outs_up[35] ,
    \ces_1_4_io_outs_up[34] ,
    \ces_1_4_io_outs_up[33] ,
    \ces_1_4_io_outs_up[32] ,
    \ces_1_4_io_outs_up[31] ,
    \ces_1_4_io_outs_up[30] ,
    \ces_1_4_io_outs_up[29] ,
    \ces_1_4_io_outs_up[28] ,
    \ces_1_4_io_outs_up[27] ,
    \ces_1_4_io_outs_up[26] ,
    \ces_1_4_io_outs_up[25] ,
    \ces_1_4_io_outs_up[24] ,
    \ces_1_4_io_outs_up[23] ,
    \ces_1_4_io_outs_up[22] ,
    \ces_1_4_io_outs_up[21] ,
    \ces_1_4_io_outs_up[20] ,
    \ces_1_4_io_outs_up[19] ,
    \ces_1_4_io_outs_up[18] ,
    \ces_1_4_io_outs_up[17] ,
    \ces_1_4_io_outs_up[16] ,
    \ces_1_4_io_outs_up[15] ,
    \ces_1_4_io_outs_up[14] ,
    \ces_1_4_io_outs_up[13] ,
    \ces_1_4_io_outs_up[12] ,
    \ces_1_4_io_outs_up[11] ,
    \ces_1_4_io_outs_up[10] ,
    \ces_1_4_io_outs_up[9] ,
    \ces_1_4_io_outs_up[8] ,
    \ces_1_4_io_outs_up[7] ,
    \ces_1_4_io_outs_up[6] ,
    \ces_1_4_io_outs_up[5] ,
    \ces_1_4_io_outs_up[4] ,
    \ces_1_4_io_outs_up[3] ,
    \ces_1_4_io_outs_up[2] ,
    \ces_1_4_io_outs_up[1] ,
    \ces_1_4_io_outs_up[0] }));
 Element ces_1_5 (.clock(clknet_3_2_0_clock),
    .io_lsbIns_1(ces_1_4_io_lsbOuts_1),
    .io_lsbIns_2(ces_1_4_io_lsbOuts_2),
    .io_lsbIns_3(ces_1_4_io_lsbOuts_3),
    .io_lsbIns_4(ces_1_4_io_lsbOuts_4),
    .io_lsbIns_5(ces_1_4_io_lsbOuts_5),
    .io_lsbIns_6(ces_1_4_io_lsbOuts_6),
    .io_lsbIns_7(ces_1_4_io_lsbOuts_7),
    .io_lsbOuts_0(ces_1_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_5_io_lsbOuts_7),
    .io_ins_down({\ces_1_5_io_ins_down[63] ,
    \ces_1_5_io_ins_down[62] ,
    \ces_1_5_io_ins_down[61] ,
    \ces_1_5_io_ins_down[60] ,
    \ces_1_5_io_ins_down[59] ,
    \ces_1_5_io_ins_down[58] ,
    \ces_1_5_io_ins_down[57] ,
    \ces_1_5_io_ins_down[56] ,
    \ces_1_5_io_ins_down[55] ,
    \ces_1_5_io_ins_down[54] ,
    \ces_1_5_io_ins_down[53] ,
    \ces_1_5_io_ins_down[52] ,
    \ces_1_5_io_ins_down[51] ,
    \ces_1_5_io_ins_down[50] ,
    \ces_1_5_io_ins_down[49] ,
    \ces_1_5_io_ins_down[48] ,
    \ces_1_5_io_ins_down[47] ,
    \ces_1_5_io_ins_down[46] ,
    \ces_1_5_io_ins_down[45] ,
    \ces_1_5_io_ins_down[44] ,
    \ces_1_5_io_ins_down[43] ,
    \ces_1_5_io_ins_down[42] ,
    \ces_1_5_io_ins_down[41] ,
    \ces_1_5_io_ins_down[40] ,
    \ces_1_5_io_ins_down[39] ,
    \ces_1_5_io_ins_down[38] ,
    \ces_1_5_io_ins_down[37] ,
    \ces_1_5_io_ins_down[36] ,
    \ces_1_5_io_ins_down[35] ,
    \ces_1_5_io_ins_down[34] ,
    \ces_1_5_io_ins_down[33] ,
    \ces_1_5_io_ins_down[32] ,
    \ces_1_5_io_ins_down[31] ,
    \ces_1_5_io_ins_down[30] ,
    \ces_1_5_io_ins_down[29] ,
    \ces_1_5_io_ins_down[28] ,
    \ces_1_5_io_ins_down[27] ,
    \ces_1_5_io_ins_down[26] ,
    \ces_1_5_io_ins_down[25] ,
    \ces_1_5_io_ins_down[24] ,
    \ces_1_5_io_ins_down[23] ,
    \ces_1_5_io_ins_down[22] ,
    \ces_1_5_io_ins_down[21] ,
    \ces_1_5_io_ins_down[20] ,
    \ces_1_5_io_ins_down[19] ,
    \ces_1_5_io_ins_down[18] ,
    \ces_1_5_io_ins_down[17] ,
    \ces_1_5_io_ins_down[16] ,
    \ces_1_5_io_ins_down[15] ,
    \ces_1_5_io_ins_down[14] ,
    \ces_1_5_io_ins_down[13] ,
    \ces_1_5_io_ins_down[12] ,
    \ces_1_5_io_ins_down[11] ,
    \ces_1_5_io_ins_down[10] ,
    \ces_1_5_io_ins_down[9] ,
    \ces_1_5_io_ins_down[8] ,
    \ces_1_5_io_ins_down[7] ,
    \ces_1_5_io_ins_down[6] ,
    \ces_1_5_io_ins_down[5] ,
    \ces_1_5_io_ins_down[4] ,
    \ces_1_5_io_ins_down[3] ,
    \ces_1_5_io_ins_down[2] ,
    \ces_1_5_io_ins_down[1] ,
    \ces_1_5_io_ins_down[0] }),
    .io_ins_left({\ces_1_5_io_ins_left[63] ,
    \ces_1_5_io_ins_left[62] ,
    \ces_1_5_io_ins_left[61] ,
    \ces_1_5_io_ins_left[60] ,
    \ces_1_5_io_ins_left[59] ,
    \ces_1_5_io_ins_left[58] ,
    \ces_1_5_io_ins_left[57] ,
    \ces_1_5_io_ins_left[56] ,
    \ces_1_5_io_ins_left[55] ,
    \ces_1_5_io_ins_left[54] ,
    \ces_1_5_io_ins_left[53] ,
    \ces_1_5_io_ins_left[52] ,
    \ces_1_5_io_ins_left[51] ,
    \ces_1_5_io_ins_left[50] ,
    \ces_1_5_io_ins_left[49] ,
    \ces_1_5_io_ins_left[48] ,
    \ces_1_5_io_ins_left[47] ,
    \ces_1_5_io_ins_left[46] ,
    \ces_1_5_io_ins_left[45] ,
    \ces_1_5_io_ins_left[44] ,
    \ces_1_5_io_ins_left[43] ,
    \ces_1_5_io_ins_left[42] ,
    \ces_1_5_io_ins_left[41] ,
    \ces_1_5_io_ins_left[40] ,
    \ces_1_5_io_ins_left[39] ,
    \ces_1_5_io_ins_left[38] ,
    \ces_1_5_io_ins_left[37] ,
    \ces_1_5_io_ins_left[36] ,
    \ces_1_5_io_ins_left[35] ,
    \ces_1_5_io_ins_left[34] ,
    \ces_1_5_io_ins_left[33] ,
    \ces_1_5_io_ins_left[32] ,
    \ces_1_5_io_ins_left[31] ,
    \ces_1_5_io_ins_left[30] ,
    \ces_1_5_io_ins_left[29] ,
    \ces_1_5_io_ins_left[28] ,
    \ces_1_5_io_ins_left[27] ,
    \ces_1_5_io_ins_left[26] ,
    \ces_1_5_io_ins_left[25] ,
    \ces_1_5_io_ins_left[24] ,
    \ces_1_5_io_ins_left[23] ,
    \ces_1_5_io_ins_left[22] ,
    \ces_1_5_io_ins_left[21] ,
    \ces_1_5_io_ins_left[20] ,
    \ces_1_5_io_ins_left[19] ,
    \ces_1_5_io_ins_left[18] ,
    \ces_1_5_io_ins_left[17] ,
    \ces_1_5_io_ins_left[16] ,
    \ces_1_5_io_ins_left[15] ,
    \ces_1_5_io_ins_left[14] ,
    \ces_1_5_io_ins_left[13] ,
    \ces_1_5_io_ins_left[12] ,
    \ces_1_5_io_ins_left[11] ,
    \ces_1_5_io_ins_left[10] ,
    \ces_1_5_io_ins_left[9] ,
    \ces_1_5_io_ins_left[8] ,
    \ces_1_5_io_ins_left[7] ,
    \ces_1_5_io_ins_left[6] ,
    \ces_1_5_io_ins_left[5] ,
    \ces_1_5_io_ins_left[4] ,
    \ces_1_5_io_ins_left[3] ,
    \ces_1_5_io_ins_left[2] ,
    \ces_1_5_io_ins_left[1] ,
    \ces_1_5_io_ins_left[0] }),
    .io_ins_right({\ces_1_4_io_outs_right[63] ,
    \ces_1_4_io_outs_right[62] ,
    \ces_1_4_io_outs_right[61] ,
    \ces_1_4_io_outs_right[60] ,
    \ces_1_4_io_outs_right[59] ,
    \ces_1_4_io_outs_right[58] ,
    \ces_1_4_io_outs_right[57] ,
    \ces_1_4_io_outs_right[56] ,
    \ces_1_4_io_outs_right[55] ,
    \ces_1_4_io_outs_right[54] ,
    \ces_1_4_io_outs_right[53] ,
    \ces_1_4_io_outs_right[52] ,
    \ces_1_4_io_outs_right[51] ,
    \ces_1_4_io_outs_right[50] ,
    \ces_1_4_io_outs_right[49] ,
    \ces_1_4_io_outs_right[48] ,
    \ces_1_4_io_outs_right[47] ,
    \ces_1_4_io_outs_right[46] ,
    \ces_1_4_io_outs_right[45] ,
    \ces_1_4_io_outs_right[44] ,
    \ces_1_4_io_outs_right[43] ,
    \ces_1_4_io_outs_right[42] ,
    \ces_1_4_io_outs_right[41] ,
    \ces_1_4_io_outs_right[40] ,
    \ces_1_4_io_outs_right[39] ,
    \ces_1_4_io_outs_right[38] ,
    \ces_1_4_io_outs_right[37] ,
    \ces_1_4_io_outs_right[36] ,
    \ces_1_4_io_outs_right[35] ,
    \ces_1_4_io_outs_right[34] ,
    \ces_1_4_io_outs_right[33] ,
    \ces_1_4_io_outs_right[32] ,
    \ces_1_4_io_outs_right[31] ,
    \ces_1_4_io_outs_right[30] ,
    \ces_1_4_io_outs_right[29] ,
    \ces_1_4_io_outs_right[28] ,
    \ces_1_4_io_outs_right[27] ,
    \ces_1_4_io_outs_right[26] ,
    \ces_1_4_io_outs_right[25] ,
    \ces_1_4_io_outs_right[24] ,
    \ces_1_4_io_outs_right[23] ,
    \ces_1_4_io_outs_right[22] ,
    \ces_1_4_io_outs_right[21] ,
    \ces_1_4_io_outs_right[20] ,
    \ces_1_4_io_outs_right[19] ,
    \ces_1_4_io_outs_right[18] ,
    \ces_1_4_io_outs_right[17] ,
    \ces_1_4_io_outs_right[16] ,
    \ces_1_4_io_outs_right[15] ,
    \ces_1_4_io_outs_right[14] ,
    \ces_1_4_io_outs_right[13] ,
    \ces_1_4_io_outs_right[12] ,
    \ces_1_4_io_outs_right[11] ,
    \ces_1_4_io_outs_right[10] ,
    \ces_1_4_io_outs_right[9] ,
    \ces_1_4_io_outs_right[8] ,
    \ces_1_4_io_outs_right[7] ,
    \ces_1_4_io_outs_right[6] ,
    \ces_1_4_io_outs_right[5] ,
    \ces_1_4_io_outs_right[4] ,
    \ces_1_4_io_outs_right[3] ,
    \ces_1_4_io_outs_right[2] ,
    \ces_1_4_io_outs_right[1] ,
    \ces_1_4_io_outs_right[0] }),
    .io_ins_up({\ces_0_5_io_outs_up[63] ,
    \ces_0_5_io_outs_up[62] ,
    \ces_0_5_io_outs_up[61] ,
    \ces_0_5_io_outs_up[60] ,
    \ces_0_5_io_outs_up[59] ,
    \ces_0_5_io_outs_up[58] ,
    \ces_0_5_io_outs_up[57] ,
    \ces_0_5_io_outs_up[56] ,
    \ces_0_5_io_outs_up[55] ,
    \ces_0_5_io_outs_up[54] ,
    \ces_0_5_io_outs_up[53] ,
    \ces_0_5_io_outs_up[52] ,
    \ces_0_5_io_outs_up[51] ,
    \ces_0_5_io_outs_up[50] ,
    \ces_0_5_io_outs_up[49] ,
    \ces_0_5_io_outs_up[48] ,
    \ces_0_5_io_outs_up[47] ,
    \ces_0_5_io_outs_up[46] ,
    \ces_0_5_io_outs_up[45] ,
    \ces_0_5_io_outs_up[44] ,
    \ces_0_5_io_outs_up[43] ,
    \ces_0_5_io_outs_up[42] ,
    \ces_0_5_io_outs_up[41] ,
    \ces_0_5_io_outs_up[40] ,
    \ces_0_5_io_outs_up[39] ,
    \ces_0_5_io_outs_up[38] ,
    \ces_0_5_io_outs_up[37] ,
    \ces_0_5_io_outs_up[36] ,
    \ces_0_5_io_outs_up[35] ,
    \ces_0_5_io_outs_up[34] ,
    \ces_0_5_io_outs_up[33] ,
    \ces_0_5_io_outs_up[32] ,
    \ces_0_5_io_outs_up[31] ,
    \ces_0_5_io_outs_up[30] ,
    \ces_0_5_io_outs_up[29] ,
    \ces_0_5_io_outs_up[28] ,
    \ces_0_5_io_outs_up[27] ,
    \ces_0_5_io_outs_up[26] ,
    \ces_0_5_io_outs_up[25] ,
    \ces_0_5_io_outs_up[24] ,
    \ces_0_5_io_outs_up[23] ,
    \ces_0_5_io_outs_up[22] ,
    \ces_0_5_io_outs_up[21] ,
    \ces_0_5_io_outs_up[20] ,
    \ces_0_5_io_outs_up[19] ,
    \ces_0_5_io_outs_up[18] ,
    \ces_0_5_io_outs_up[17] ,
    \ces_0_5_io_outs_up[16] ,
    \ces_0_5_io_outs_up[15] ,
    \ces_0_5_io_outs_up[14] ,
    \ces_0_5_io_outs_up[13] ,
    \ces_0_5_io_outs_up[12] ,
    \ces_0_5_io_outs_up[11] ,
    \ces_0_5_io_outs_up[10] ,
    \ces_0_5_io_outs_up[9] ,
    \ces_0_5_io_outs_up[8] ,
    \ces_0_5_io_outs_up[7] ,
    \ces_0_5_io_outs_up[6] ,
    \ces_0_5_io_outs_up[5] ,
    \ces_0_5_io_outs_up[4] ,
    \ces_0_5_io_outs_up[3] ,
    \ces_0_5_io_outs_up[2] ,
    \ces_0_5_io_outs_up[1] ,
    \ces_0_5_io_outs_up[0] }),
    .io_outs_down({\ces_0_5_io_ins_down[63] ,
    \ces_0_5_io_ins_down[62] ,
    \ces_0_5_io_ins_down[61] ,
    \ces_0_5_io_ins_down[60] ,
    \ces_0_5_io_ins_down[59] ,
    \ces_0_5_io_ins_down[58] ,
    \ces_0_5_io_ins_down[57] ,
    \ces_0_5_io_ins_down[56] ,
    \ces_0_5_io_ins_down[55] ,
    \ces_0_5_io_ins_down[54] ,
    \ces_0_5_io_ins_down[53] ,
    \ces_0_5_io_ins_down[52] ,
    \ces_0_5_io_ins_down[51] ,
    \ces_0_5_io_ins_down[50] ,
    \ces_0_5_io_ins_down[49] ,
    \ces_0_5_io_ins_down[48] ,
    \ces_0_5_io_ins_down[47] ,
    \ces_0_5_io_ins_down[46] ,
    \ces_0_5_io_ins_down[45] ,
    \ces_0_5_io_ins_down[44] ,
    \ces_0_5_io_ins_down[43] ,
    \ces_0_5_io_ins_down[42] ,
    \ces_0_5_io_ins_down[41] ,
    \ces_0_5_io_ins_down[40] ,
    \ces_0_5_io_ins_down[39] ,
    \ces_0_5_io_ins_down[38] ,
    \ces_0_5_io_ins_down[37] ,
    \ces_0_5_io_ins_down[36] ,
    \ces_0_5_io_ins_down[35] ,
    \ces_0_5_io_ins_down[34] ,
    \ces_0_5_io_ins_down[33] ,
    \ces_0_5_io_ins_down[32] ,
    \ces_0_5_io_ins_down[31] ,
    \ces_0_5_io_ins_down[30] ,
    \ces_0_5_io_ins_down[29] ,
    \ces_0_5_io_ins_down[28] ,
    \ces_0_5_io_ins_down[27] ,
    \ces_0_5_io_ins_down[26] ,
    \ces_0_5_io_ins_down[25] ,
    \ces_0_5_io_ins_down[24] ,
    \ces_0_5_io_ins_down[23] ,
    \ces_0_5_io_ins_down[22] ,
    \ces_0_5_io_ins_down[21] ,
    \ces_0_5_io_ins_down[20] ,
    \ces_0_5_io_ins_down[19] ,
    \ces_0_5_io_ins_down[18] ,
    \ces_0_5_io_ins_down[17] ,
    \ces_0_5_io_ins_down[16] ,
    \ces_0_5_io_ins_down[15] ,
    \ces_0_5_io_ins_down[14] ,
    \ces_0_5_io_ins_down[13] ,
    \ces_0_5_io_ins_down[12] ,
    \ces_0_5_io_ins_down[11] ,
    \ces_0_5_io_ins_down[10] ,
    \ces_0_5_io_ins_down[9] ,
    \ces_0_5_io_ins_down[8] ,
    \ces_0_5_io_ins_down[7] ,
    \ces_0_5_io_ins_down[6] ,
    \ces_0_5_io_ins_down[5] ,
    \ces_0_5_io_ins_down[4] ,
    \ces_0_5_io_ins_down[3] ,
    \ces_0_5_io_ins_down[2] ,
    \ces_0_5_io_ins_down[1] ,
    \ces_0_5_io_ins_down[0] }),
    .io_outs_left({\ces_1_4_io_ins_left[63] ,
    \ces_1_4_io_ins_left[62] ,
    \ces_1_4_io_ins_left[61] ,
    \ces_1_4_io_ins_left[60] ,
    \ces_1_4_io_ins_left[59] ,
    \ces_1_4_io_ins_left[58] ,
    \ces_1_4_io_ins_left[57] ,
    \ces_1_4_io_ins_left[56] ,
    \ces_1_4_io_ins_left[55] ,
    \ces_1_4_io_ins_left[54] ,
    \ces_1_4_io_ins_left[53] ,
    \ces_1_4_io_ins_left[52] ,
    \ces_1_4_io_ins_left[51] ,
    \ces_1_4_io_ins_left[50] ,
    \ces_1_4_io_ins_left[49] ,
    \ces_1_4_io_ins_left[48] ,
    \ces_1_4_io_ins_left[47] ,
    \ces_1_4_io_ins_left[46] ,
    \ces_1_4_io_ins_left[45] ,
    \ces_1_4_io_ins_left[44] ,
    \ces_1_4_io_ins_left[43] ,
    \ces_1_4_io_ins_left[42] ,
    \ces_1_4_io_ins_left[41] ,
    \ces_1_4_io_ins_left[40] ,
    \ces_1_4_io_ins_left[39] ,
    \ces_1_4_io_ins_left[38] ,
    \ces_1_4_io_ins_left[37] ,
    \ces_1_4_io_ins_left[36] ,
    \ces_1_4_io_ins_left[35] ,
    \ces_1_4_io_ins_left[34] ,
    \ces_1_4_io_ins_left[33] ,
    \ces_1_4_io_ins_left[32] ,
    \ces_1_4_io_ins_left[31] ,
    \ces_1_4_io_ins_left[30] ,
    \ces_1_4_io_ins_left[29] ,
    \ces_1_4_io_ins_left[28] ,
    \ces_1_4_io_ins_left[27] ,
    \ces_1_4_io_ins_left[26] ,
    \ces_1_4_io_ins_left[25] ,
    \ces_1_4_io_ins_left[24] ,
    \ces_1_4_io_ins_left[23] ,
    \ces_1_4_io_ins_left[22] ,
    \ces_1_4_io_ins_left[21] ,
    \ces_1_4_io_ins_left[20] ,
    \ces_1_4_io_ins_left[19] ,
    \ces_1_4_io_ins_left[18] ,
    \ces_1_4_io_ins_left[17] ,
    \ces_1_4_io_ins_left[16] ,
    \ces_1_4_io_ins_left[15] ,
    \ces_1_4_io_ins_left[14] ,
    \ces_1_4_io_ins_left[13] ,
    \ces_1_4_io_ins_left[12] ,
    \ces_1_4_io_ins_left[11] ,
    \ces_1_4_io_ins_left[10] ,
    \ces_1_4_io_ins_left[9] ,
    \ces_1_4_io_ins_left[8] ,
    \ces_1_4_io_ins_left[7] ,
    \ces_1_4_io_ins_left[6] ,
    \ces_1_4_io_ins_left[5] ,
    \ces_1_4_io_ins_left[4] ,
    \ces_1_4_io_ins_left[3] ,
    \ces_1_4_io_ins_left[2] ,
    \ces_1_4_io_ins_left[1] ,
    \ces_1_4_io_ins_left[0] }),
    .io_outs_right({\ces_1_5_io_outs_right[63] ,
    \ces_1_5_io_outs_right[62] ,
    \ces_1_5_io_outs_right[61] ,
    \ces_1_5_io_outs_right[60] ,
    \ces_1_5_io_outs_right[59] ,
    \ces_1_5_io_outs_right[58] ,
    \ces_1_5_io_outs_right[57] ,
    \ces_1_5_io_outs_right[56] ,
    \ces_1_5_io_outs_right[55] ,
    \ces_1_5_io_outs_right[54] ,
    \ces_1_5_io_outs_right[53] ,
    \ces_1_5_io_outs_right[52] ,
    \ces_1_5_io_outs_right[51] ,
    \ces_1_5_io_outs_right[50] ,
    \ces_1_5_io_outs_right[49] ,
    \ces_1_5_io_outs_right[48] ,
    \ces_1_5_io_outs_right[47] ,
    \ces_1_5_io_outs_right[46] ,
    \ces_1_5_io_outs_right[45] ,
    \ces_1_5_io_outs_right[44] ,
    \ces_1_5_io_outs_right[43] ,
    \ces_1_5_io_outs_right[42] ,
    \ces_1_5_io_outs_right[41] ,
    \ces_1_5_io_outs_right[40] ,
    \ces_1_5_io_outs_right[39] ,
    \ces_1_5_io_outs_right[38] ,
    \ces_1_5_io_outs_right[37] ,
    \ces_1_5_io_outs_right[36] ,
    \ces_1_5_io_outs_right[35] ,
    \ces_1_5_io_outs_right[34] ,
    \ces_1_5_io_outs_right[33] ,
    \ces_1_5_io_outs_right[32] ,
    \ces_1_5_io_outs_right[31] ,
    \ces_1_5_io_outs_right[30] ,
    \ces_1_5_io_outs_right[29] ,
    \ces_1_5_io_outs_right[28] ,
    \ces_1_5_io_outs_right[27] ,
    \ces_1_5_io_outs_right[26] ,
    \ces_1_5_io_outs_right[25] ,
    \ces_1_5_io_outs_right[24] ,
    \ces_1_5_io_outs_right[23] ,
    \ces_1_5_io_outs_right[22] ,
    \ces_1_5_io_outs_right[21] ,
    \ces_1_5_io_outs_right[20] ,
    \ces_1_5_io_outs_right[19] ,
    \ces_1_5_io_outs_right[18] ,
    \ces_1_5_io_outs_right[17] ,
    \ces_1_5_io_outs_right[16] ,
    \ces_1_5_io_outs_right[15] ,
    \ces_1_5_io_outs_right[14] ,
    \ces_1_5_io_outs_right[13] ,
    \ces_1_5_io_outs_right[12] ,
    \ces_1_5_io_outs_right[11] ,
    \ces_1_5_io_outs_right[10] ,
    \ces_1_5_io_outs_right[9] ,
    \ces_1_5_io_outs_right[8] ,
    \ces_1_5_io_outs_right[7] ,
    \ces_1_5_io_outs_right[6] ,
    \ces_1_5_io_outs_right[5] ,
    \ces_1_5_io_outs_right[4] ,
    \ces_1_5_io_outs_right[3] ,
    \ces_1_5_io_outs_right[2] ,
    \ces_1_5_io_outs_right[1] ,
    \ces_1_5_io_outs_right[0] }),
    .io_outs_up({\ces_1_5_io_outs_up[63] ,
    \ces_1_5_io_outs_up[62] ,
    \ces_1_5_io_outs_up[61] ,
    \ces_1_5_io_outs_up[60] ,
    \ces_1_5_io_outs_up[59] ,
    \ces_1_5_io_outs_up[58] ,
    \ces_1_5_io_outs_up[57] ,
    \ces_1_5_io_outs_up[56] ,
    \ces_1_5_io_outs_up[55] ,
    \ces_1_5_io_outs_up[54] ,
    \ces_1_5_io_outs_up[53] ,
    \ces_1_5_io_outs_up[52] ,
    \ces_1_5_io_outs_up[51] ,
    \ces_1_5_io_outs_up[50] ,
    \ces_1_5_io_outs_up[49] ,
    \ces_1_5_io_outs_up[48] ,
    \ces_1_5_io_outs_up[47] ,
    \ces_1_5_io_outs_up[46] ,
    \ces_1_5_io_outs_up[45] ,
    \ces_1_5_io_outs_up[44] ,
    \ces_1_5_io_outs_up[43] ,
    \ces_1_5_io_outs_up[42] ,
    \ces_1_5_io_outs_up[41] ,
    \ces_1_5_io_outs_up[40] ,
    \ces_1_5_io_outs_up[39] ,
    \ces_1_5_io_outs_up[38] ,
    \ces_1_5_io_outs_up[37] ,
    \ces_1_5_io_outs_up[36] ,
    \ces_1_5_io_outs_up[35] ,
    \ces_1_5_io_outs_up[34] ,
    \ces_1_5_io_outs_up[33] ,
    \ces_1_5_io_outs_up[32] ,
    \ces_1_5_io_outs_up[31] ,
    \ces_1_5_io_outs_up[30] ,
    \ces_1_5_io_outs_up[29] ,
    \ces_1_5_io_outs_up[28] ,
    \ces_1_5_io_outs_up[27] ,
    \ces_1_5_io_outs_up[26] ,
    \ces_1_5_io_outs_up[25] ,
    \ces_1_5_io_outs_up[24] ,
    \ces_1_5_io_outs_up[23] ,
    \ces_1_5_io_outs_up[22] ,
    \ces_1_5_io_outs_up[21] ,
    \ces_1_5_io_outs_up[20] ,
    \ces_1_5_io_outs_up[19] ,
    \ces_1_5_io_outs_up[18] ,
    \ces_1_5_io_outs_up[17] ,
    \ces_1_5_io_outs_up[16] ,
    \ces_1_5_io_outs_up[15] ,
    \ces_1_5_io_outs_up[14] ,
    \ces_1_5_io_outs_up[13] ,
    \ces_1_5_io_outs_up[12] ,
    \ces_1_5_io_outs_up[11] ,
    \ces_1_5_io_outs_up[10] ,
    \ces_1_5_io_outs_up[9] ,
    \ces_1_5_io_outs_up[8] ,
    \ces_1_5_io_outs_up[7] ,
    \ces_1_5_io_outs_up[6] ,
    \ces_1_5_io_outs_up[5] ,
    \ces_1_5_io_outs_up[4] ,
    \ces_1_5_io_outs_up[3] ,
    \ces_1_5_io_outs_up[2] ,
    \ces_1_5_io_outs_up[1] ,
    \ces_1_5_io_outs_up[0] }));
 Element ces_1_6 (.clock(clknet_3_2_0_clock),
    .io_lsbIns_1(ces_1_5_io_lsbOuts_1),
    .io_lsbIns_2(ces_1_5_io_lsbOuts_2),
    .io_lsbIns_3(ces_1_5_io_lsbOuts_3),
    .io_lsbIns_4(ces_1_5_io_lsbOuts_4),
    .io_lsbIns_5(ces_1_5_io_lsbOuts_5),
    .io_lsbIns_6(ces_1_5_io_lsbOuts_6),
    .io_lsbIns_7(ces_1_5_io_lsbOuts_7),
    .io_lsbOuts_0(ces_1_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_6_io_lsbOuts_7),
    .io_ins_down({\ces_1_6_io_ins_down[63] ,
    \ces_1_6_io_ins_down[62] ,
    \ces_1_6_io_ins_down[61] ,
    \ces_1_6_io_ins_down[60] ,
    \ces_1_6_io_ins_down[59] ,
    \ces_1_6_io_ins_down[58] ,
    \ces_1_6_io_ins_down[57] ,
    \ces_1_6_io_ins_down[56] ,
    \ces_1_6_io_ins_down[55] ,
    \ces_1_6_io_ins_down[54] ,
    \ces_1_6_io_ins_down[53] ,
    \ces_1_6_io_ins_down[52] ,
    \ces_1_6_io_ins_down[51] ,
    \ces_1_6_io_ins_down[50] ,
    \ces_1_6_io_ins_down[49] ,
    \ces_1_6_io_ins_down[48] ,
    \ces_1_6_io_ins_down[47] ,
    \ces_1_6_io_ins_down[46] ,
    \ces_1_6_io_ins_down[45] ,
    \ces_1_6_io_ins_down[44] ,
    \ces_1_6_io_ins_down[43] ,
    \ces_1_6_io_ins_down[42] ,
    \ces_1_6_io_ins_down[41] ,
    \ces_1_6_io_ins_down[40] ,
    \ces_1_6_io_ins_down[39] ,
    \ces_1_6_io_ins_down[38] ,
    \ces_1_6_io_ins_down[37] ,
    \ces_1_6_io_ins_down[36] ,
    \ces_1_6_io_ins_down[35] ,
    \ces_1_6_io_ins_down[34] ,
    \ces_1_6_io_ins_down[33] ,
    \ces_1_6_io_ins_down[32] ,
    \ces_1_6_io_ins_down[31] ,
    \ces_1_6_io_ins_down[30] ,
    \ces_1_6_io_ins_down[29] ,
    \ces_1_6_io_ins_down[28] ,
    \ces_1_6_io_ins_down[27] ,
    \ces_1_6_io_ins_down[26] ,
    \ces_1_6_io_ins_down[25] ,
    \ces_1_6_io_ins_down[24] ,
    \ces_1_6_io_ins_down[23] ,
    \ces_1_6_io_ins_down[22] ,
    \ces_1_6_io_ins_down[21] ,
    \ces_1_6_io_ins_down[20] ,
    \ces_1_6_io_ins_down[19] ,
    \ces_1_6_io_ins_down[18] ,
    \ces_1_6_io_ins_down[17] ,
    \ces_1_6_io_ins_down[16] ,
    \ces_1_6_io_ins_down[15] ,
    \ces_1_6_io_ins_down[14] ,
    \ces_1_6_io_ins_down[13] ,
    \ces_1_6_io_ins_down[12] ,
    \ces_1_6_io_ins_down[11] ,
    \ces_1_6_io_ins_down[10] ,
    \ces_1_6_io_ins_down[9] ,
    \ces_1_6_io_ins_down[8] ,
    \ces_1_6_io_ins_down[7] ,
    \ces_1_6_io_ins_down[6] ,
    \ces_1_6_io_ins_down[5] ,
    \ces_1_6_io_ins_down[4] ,
    \ces_1_6_io_ins_down[3] ,
    \ces_1_6_io_ins_down[2] ,
    \ces_1_6_io_ins_down[1] ,
    \ces_1_6_io_ins_down[0] }),
    .io_ins_left({\ces_1_6_io_ins_left[63] ,
    \ces_1_6_io_ins_left[62] ,
    \ces_1_6_io_ins_left[61] ,
    \ces_1_6_io_ins_left[60] ,
    \ces_1_6_io_ins_left[59] ,
    \ces_1_6_io_ins_left[58] ,
    \ces_1_6_io_ins_left[57] ,
    \ces_1_6_io_ins_left[56] ,
    \ces_1_6_io_ins_left[55] ,
    \ces_1_6_io_ins_left[54] ,
    \ces_1_6_io_ins_left[53] ,
    \ces_1_6_io_ins_left[52] ,
    \ces_1_6_io_ins_left[51] ,
    \ces_1_6_io_ins_left[50] ,
    \ces_1_6_io_ins_left[49] ,
    \ces_1_6_io_ins_left[48] ,
    \ces_1_6_io_ins_left[47] ,
    \ces_1_6_io_ins_left[46] ,
    \ces_1_6_io_ins_left[45] ,
    \ces_1_6_io_ins_left[44] ,
    \ces_1_6_io_ins_left[43] ,
    \ces_1_6_io_ins_left[42] ,
    \ces_1_6_io_ins_left[41] ,
    \ces_1_6_io_ins_left[40] ,
    \ces_1_6_io_ins_left[39] ,
    \ces_1_6_io_ins_left[38] ,
    \ces_1_6_io_ins_left[37] ,
    \ces_1_6_io_ins_left[36] ,
    \ces_1_6_io_ins_left[35] ,
    \ces_1_6_io_ins_left[34] ,
    \ces_1_6_io_ins_left[33] ,
    \ces_1_6_io_ins_left[32] ,
    \ces_1_6_io_ins_left[31] ,
    \ces_1_6_io_ins_left[30] ,
    \ces_1_6_io_ins_left[29] ,
    \ces_1_6_io_ins_left[28] ,
    \ces_1_6_io_ins_left[27] ,
    \ces_1_6_io_ins_left[26] ,
    \ces_1_6_io_ins_left[25] ,
    \ces_1_6_io_ins_left[24] ,
    \ces_1_6_io_ins_left[23] ,
    \ces_1_6_io_ins_left[22] ,
    \ces_1_6_io_ins_left[21] ,
    \ces_1_6_io_ins_left[20] ,
    \ces_1_6_io_ins_left[19] ,
    \ces_1_6_io_ins_left[18] ,
    \ces_1_6_io_ins_left[17] ,
    \ces_1_6_io_ins_left[16] ,
    \ces_1_6_io_ins_left[15] ,
    \ces_1_6_io_ins_left[14] ,
    \ces_1_6_io_ins_left[13] ,
    \ces_1_6_io_ins_left[12] ,
    \ces_1_6_io_ins_left[11] ,
    \ces_1_6_io_ins_left[10] ,
    \ces_1_6_io_ins_left[9] ,
    \ces_1_6_io_ins_left[8] ,
    \ces_1_6_io_ins_left[7] ,
    \ces_1_6_io_ins_left[6] ,
    \ces_1_6_io_ins_left[5] ,
    \ces_1_6_io_ins_left[4] ,
    \ces_1_6_io_ins_left[3] ,
    \ces_1_6_io_ins_left[2] ,
    \ces_1_6_io_ins_left[1] ,
    \ces_1_6_io_ins_left[0] }),
    .io_ins_right({\ces_1_5_io_outs_right[63] ,
    \ces_1_5_io_outs_right[62] ,
    \ces_1_5_io_outs_right[61] ,
    \ces_1_5_io_outs_right[60] ,
    \ces_1_5_io_outs_right[59] ,
    \ces_1_5_io_outs_right[58] ,
    \ces_1_5_io_outs_right[57] ,
    \ces_1_5_io_outs_right[56] ,
    \ces_1_5_io_outs_right[55] ,
    \ces_1_5_io_outs_right[54] ,
    \ces_1_5_io_outs_right[53] ,
    \ces_1_5_io_outs_right[52] ,
    \ces_1_5_io_outs_right[51] ,
    \ces_1_5_io_outs_right[50] ,
    \ces_1_5_io_outs_right[49] ,
    \ces_1_5_io_outs_right[48] ,
    \ces_1_5_io_outs_right[47] ,
    \ces_1_5_io_outs_right[46] ,
    \ces_1_5_io_outs_right[45] ,
    \ces_1_5_io_outs_right[44] ,
    \ces_1_5_io_outs_right[43] ,
    \ces_1_5_io_outs_right[42] ,
    \ces_1_5_io_outs_right[41] ,
    \ces_1_5_io_outs_right[40] ,
    \ces_1_5_io_outs_right[39] ,
    \ces_1_5_io_outs_right[38] ,
    \ces_1_5_io_outs_right[37] ,
    \ces_1_5_io_outs_right[36] ,
    \ces_1_5_io_outs_right[35] ,
    \ces_1_5_io_outs_right[34] ,
    \ces_1_5_io_outs_right[33] ,
    \ces_1_5_io_outs_right[32] ,
    \ces_1_5_io_outs_right[31] ,
    \ces_1_5_io_outs_right[30] ,
    \ces_1_5_io_outs_right[29] ,
    \ces_1_5_io_outs_right[28] ,
    \ces_1_5_io_outs_right[27] ,
    \ces_1_5_io_outs_right[26] ,
    \ces_1_5_io_outs_right[25] ,
    \ces_1_5_io_outs_right[24] ,
    \ces_1_5_io_outs_right[23] ,
    \ces_1_5_io_outs_right[22] ,
    \ces_1_5_io_outs_right[21] ,
    \ces_1_5_io_outs_right[20] ,
    \ces_1_5_io_outs_right[19] ,
    \ces_1_5_io_outs_right[18] ,
    \ces_1_5_io_outs_right[17] ,
    \ces_1_5_io_outs_right[16] ,
    \ces_1_5_io_outs_right[15] ,
    \ces_1_5_io_outs_right[14] ,
    \ces_1_5_io_outs_right[13] ,
    \ces_1_5_io_outs_right[12] ,
    \ces_1_5_io_outs_right[11] ,
    \ces_1_5_io_outs_right[10] ,
    \ces_1_5_io_outs_right[9] ,
    \ces_1_5_io_outs_right[8] ,
    \ces_1_5_io_outs_right[7] ,
    \ces_1_5_io_outs_right[6] ,
    \ces_1_5_io_outs_right[5] ,
    \ces_1_5_io_outs_right[4] ,
    \ces_1_5_io_outs_right[3] ,
    \ces_1_5_io_outs_right[2] ,
    \ces_1_5_io_outs_right[1] ,
    \ces_1_5_io_outs_right[0] }),
    .io_ins_up({\ces_0_6_io_outs_up[63] ,
    \ces_0_6_io_outs_up[62] ,
    \ces_0_6_io_outs_up[61] ,
    \ces_0_6_io_outs_up[60] ,
    \ces_0_6_io_outs_up[59] ,
    \ces_0_6_io_outs_up[58] ,
    \ces_0_6_io_outs_up[57] ,
    \ces_0_6_io_outs_up[56] ,
    \ces_0_6_io_outs_up[55] ,
    \ces_0_6_io_outs_up[54] ,
    \ces_0_6_io_outs_up[53] ,
    \ces_0_6_io_outs_up[52] ,
    \ces_0_6_io_outs_up[51] ,
    \ces_0_6_io_outs_up[50] ,
    \ces_0_6_io_outs_up[49] ,
    \ces_0_6_io_outs_up[48] ,
    \ces_0_6_io_outs_up[47] ,
    \ces_0_6_io_outs_up[46] ,
    \ces_0_6_io_outs_up[45] ,
    \ces_0_6_io_outs_up[44] ,
    \ces_0_6_io_outs_up[43] ,
    \ces_0_6_io_outs_up[42] ,
    \ces_0_6_io_outs_up[41] ,
    \ces_0_6_io_outs_up[40] ,
    \ces_0_6_io_outs_up[39] ,
    \ces_0_6_io_outs_up[38] ,
    \ces_0_6_io_outs_up[37] ,
    \ces_0_6_io_outs_up[36] ,
    \ces_0_6_io_outs_up[35] ,
    \ces_0_6_io_outs_up[34] ,
    \ces_0_6_io_outs_up[33] ,
    \ces_0_6_io_outs_up[32] ,
    \ces_0_6_io_outs_up[31] ,
    \ces_0_6_io_outs_up[30] ,
    \ces_0_6_io_outs_up[29] ,
    \ces_0_6_io_outs_up[28] ,
    \ces_0_6_io_outs_up[27] ,
    \ces_0_6_io_outs_up[26] ,
    \ces_0_6_io_outs_up[25] ,
    \ces_0_6_io_outs_up[24] ,
    \ces_0_6_io_outs_up[23] ,
    \ces_0_6_io_outs_up[22] ,
    \ces_0_6_io_outs_up[21] ,
    \ces_0_6_io_outs_up[20] ,
    \ces_0_6_io_outs_up[19] ,
    \ces_0_6_io_outs_up[18] ,
    \ces_0_6_io_outs_up[17] ,
    \ces_0_6_io_outs_up[16] ,
    \ces_0_6_io_outs_up[15] ,
    \ces_0_6_io_outs_up[14] ,
    \ces_0_6_io_outs_up[13] ,
    \ces_0_6_io_outs_up[12] ,
    \ces_0_6_io_outs_up[11] ,
    \ces_0_6_io_outs_up[10] ,
    \ces_0_6_io_outs_up[9] ,
    \ces_0_6_io_outs_up[8] ,
    \ces_0_6_io_outs_up[7] ,
    \ces_0_6_io_outs_up[6] ,
    \ces_0_6_io_outs_up[5] ,
    \ces_0_6_io_outs_up[4] ,
    \ces_0_6_io_outs_up[3] ,
    \ces_0_6_io_outs_up[2] ,
    \ces_0_6_io_outs_up[1] ,
    \ces_0_6_io_outs_up[0] }),
    .io_outs_down({\ces_0_6_io_ins_down[63] ,
    \ces_0_6_io_ins_down[62] ,
    \ces_0_6_io_ins_down[61] ,
    \ces_0_6_io_ins_down[60] ,
    \ces_0_6_io_ins_down[59] ,
    \ces_0_6_io_ins_down[58] ,
    \ces_0_6_io_ins_down[57] ,
    \ces_0_6_io_ins_down[56] ,
    \ces_0_6_io_ins_down[55] ,
    \ces_0_6_io_ins_down[54] ,
    \ces_0_6_io_ins_down[53] ,
    \ces_0_6_io_ins_down[52] ,
    \ces_0_6_io_ins_down[51] ,
    \ces_0_6_io_ins_down[50] ,
    \ces_0_6_io_ins_down[49] ,
    \ces_0_6_io_ins_down[48] ,
    \ces_0_6_io_ins_down[47] ,
    \ces_0_6_io_ins_down[46] ,
    \ces_0_6_io_ins_down[45] ,
    \ces_0_6_io_ins_down[44] ,
    \ces_0_6_io_ins_down[43] ,
    \ces_0_6_io_ins_down[42] ,
    \ces_0_6_io_ins_down[41] ,
    \ces_0_6_io_ins_down[40] ,
    \ces_0_6_io_ins_down[39] ,
    \ces_0_6_io_ins_down[38] ,
    \ces_0_6_io_ins_down[37] ,
    \ces_0_6_io_ins_down[36] ,
    \ces_0_6_io_ins_down[35] ,
    \ces_0_6_io_ins_down[34] ,
    \ces_0_6_io_ins_down[33] ,
    \ces_0_6_io_ins_down[32] ,
    \ces_0_6_io_ins_down[31] ,
    \ces_0_6_io_ins_down[30] ,
    \ces_0_6_io_ins_down[29] ,
    \ces_0_6_io_ins_down[28] ,
    \ces_0_6_io_ins_down[27] ,
    \ces_0_6_io_ins_down[26] ,
    \ces_0_6_io_ins_down[25] ,
    \ces_0_6_io_ins_down[24] ,
    \ces_0_6_io_ins_down[23] ,
    \ces_0_6_io_ins_down[22] ,
    \ces_0_6_io_ins_down[21] ,
    \ces_0_6_io_ins_down[20] ,
    \ces_0_6_io_ins_down[19] ,
    \ces_0_6_io_ins_down[18] ,
    \ces_0_6_io_ins_down[17] ,
    \ces_0_6_io_ins_down[16] ,
    \ces_0_6_io_ins_down[15] ,
    \ces_0_6_io_ins_down[14] ,
    \ces_0_6_io_ins_down[13] ,
    \ces_0_6_io_ins_down[12] ,
    \ces_0_6_io_ins_down[11] ,
    \ces_0_6_io_ins_down[10] ,
    \ces_0_6_io_ins_down[9] ,
    \ces_0_6_io_ins_down[8] ,
    \ces_0_6_io_ins_down[7] ,
    \ces_0_6_io_ins_down[6] ,
    \ces_0_6_io_ins_down[5] ,
    \ces_0_6_io_ins_down[4] ,
    \ces_0_6_io_ins_down[3] ,
    \ces_0_6_io_ins_down[2] ,
    \ces_0_6_io_ins_down[1] ,
    \ces_0_6_io_ins_down[0] }),
    .io_outs_left({\ces_1_5_io_ins_left[63] ,
    \ces_1_5_io_ins_left[62] ,
    \ces_1_5_io_ins_left[61] ,
    \ces_1_5_io_ins_left[60] ,
    \ces_1_5_io_ins_left[59] ,
    \ces_1_5_io_ins_left[58] ,
    \ces_1_5_io_ins_left[57] ,
    \ces_1_5_io_ins_left[56] ,
    \ces_1_5_io_ins_left[55] ,
    \ces_1_5_io_ins_left[54] ,
    \ces_1_5_io_ins_left[53] ,
    \ces_1_5_io_ins_left[52] ,
    \ces_1_5_io_ins_left[51] ,
    \ces_1_5_io_ins_left[50] ,
    \ces_1_5_io_ins_left[49] ,
    \ces_1_5_io_ins_left[48] ,
    \ces_1_5_io_ins_left[47] ,
    \ces_1_5_io_ins_left[46] ,
    \ces_1_5_io_ins_left[45] ,
    \ces_1_5_io_ins_left[44] ,
    \ces_1_5_io_ins_left[43] ,
    \ces_1_5_io_ins_left[42] ,
    \ces_1_5_io_ins_left[41] ,
    \ces_1_5_io_ins_left[40] ,
    \ces_1_5_io_ins_left[39] ,
    \ces_1_5_io_ins_left[38] ,
    \ces_1_5_io_ins_left[37] ,
    \ces_1_5_io_ins_left[36] ,
    \ces_1_5_io_ins_left[35] ,
    \ces_1_5_io_ins_left[34] ,
    \ces_1_5_io_ins_left[33] ,
    \ces_1_5_io_ins_left[32] ,
    \ces_1_5_io_ins_left[31] ,
    \ces_1_5_io_ins_left[30] ,
    \ces_1_5_io_ins_left[29] ,
    \ces_1_5_io_ins_left[28] ,
    \ces_1_5_io_ins_left[27] ,
    \ces_1_5_io_ins_left[26] ,
    \ces_1_5_io_ins_left[25] ,
    \ces_1_5_io_ins_left[24] ,
    \ces_1_5_io_ins_left[23] ,
    \ces_1_5_io_ins_left[22] ,
    \ces_1_5_io_ins_left[21] ,
    \ces_1_5_io_ins_left[20] ,
    \ces_1_5_io_ins_left[19] ,
    \ces_1_5_io_ins_left[18] ,
    \ces_1_5_io_ins_left[17] ,
    \ces_1_5_io_ins_left[16] ,
    \ces_1_5_io_ins_left[15] ,
    \ces_1_5_io_ins_left[14] ,
    \ces_1_5_io_ins_left[13] ,
    \ces_1_5_io_ins_left[12] ,
    \ces_1_5_io_ins_left[11] ,
    \ces_1_5_io_ins_left[10] ,
    \ces_1_5_io_ins_left[9] ,
    \ces_1_5_io_ins_left[8] ,
    \ces_1_5_io_ins_left[7] ,
    \ces_1_5_io_ins_left[6] ,
    \ces_1_5_io_ins_left[5] ,
    \ces_1_5_io_ins_left[4] ,
    \ces_1_5_io_ins_left[3] ,
    \ces_1_5_io_ins_left[2] ,
    \ces_1_5_io_ins_left[1] ,
    \ces_1_5_io_ins_left[0] }),
    .io_outs_right({\ces_1_6_io_outs_right[63] ,
    \ces_1_6_io_outs_right[62] ,
    \ces_1_6_io_outs_right[61] ,
    \ces_1_6_io_outs_right[60] ,
    \ces_1_6_io_outs_right[59] ,
    \ces_1_6_io_outs_right[58] ,
    \ces_1_6_io_outs_right[57] ,
    \ces_1_6_io_outs_right[56] ,
    \ces_1_6_io_outs_right[55] ,
    \ces_1_6_io_outs_right[54] ,
    \ces_1_6_io_outs_right[53] ,
    \ces_1_6_io_outs_right[52] ,
    \ces_1_6_io_outs_right[51] ,
    \ces_1_6_io_outs_right[50] ,
    \ces_1_6_io_outs_right[49] ,
    \ces_1_6_io_outs_right[48] ,
    \ces_1_6_io_outs_right[47] ,
    \ces_1_6_io_outs_right[46] ,
    \ces_1_6_io_outs_right[45] ,
    \ces_1_6_io_outs_right[44] ,
    \ces_1_6_io_outs_right[43] ,
    \ces_1_6_io_outs_right[42] ,
    \ces_1_6_io_outs_right[41] ,
    \ces_1_6_io_outs_right[40] ,
    \ces_1_6_io_outs_right[39] ,
    \ces_1_6_io_outs_right[38] ,
    \ces_1_6_io_outs_right[37] ,
    \ces_1_6_io_outs_right[36] ,
    \ces_1_6_io_outs_right[35] ,
    \ces_1_6_io_outs_right[34] ,
    \ces_1_6_io_outs_right[33] ,
    \ces_1_6_io_outs_right[32] ,
    \ces_1_6_io_outs_right[31] ,
    \ces_1_6_io_outs_right[30] ,
    \ces_1_6_io_outs_right[29] ,
    \ces_1_6_io_outs_right[28] ,
    \ces_1_6_io_outs_right[27] ,
    \ces_1_6_io_outs_right[26] ,
    \ces_1_6_io_outs_right[25] ,
    \ces_1_6_io_outs_right[24] ,
    \ces_1_6_io_outs_right[23] ,
    \ces_1_6_io_outs_right[22] ,
    \ces_1_6_io_outs_right[21] ,
    \ces_1_6_io_outs_right[20] ,
    \ces_1_6_io_outs_right[19] ,
    \ces_1_6_io_outs_right[18] ,
    \ces_1_6_io_outs_right[17] ,
    \ces_1_6_io_outs_right[16] ,
    \ces_1_6_io_outs_right[15] ,
    \ces_1_6_io_outs_right[14] ,
    \ces_1_6_io_outs_right[13] ,
    \ces_1_6_io_outs_right[12] ,
    \ces_1_6_io_outs_right[11] ,
    \ces_1_6_io_outs_right[10] ,
    \ces_1_6_io_outs_right[9] ,
    \ces_1_6_io_outs_right[8] ,
    \ces_1_6_io_outs_right[7] ,
    \ces_1_6_io_outs_right[6] ,
    \ces_1_6_io_outs_right[5] ,
    \ces_1_6_io_outs_right[4] ,
    \ces_1_6_io_outs_right[3] ,
    \ces_1_6_io_outs_right[2] ,
    \ces_1_6_io_outs_right[1] ,
    \ces_1_6_io_outs_right[0] }),
    .io_outs_up({\ces_1_6_io_outs_up[63] ,
    \ces_1_6_io_outs_up[62] ,
    \ces_1_6_io_outs_up[61] ,
    \ces_1_6_io_outs_up[60] ,
    \ces_1_6_io_outs_up[59] ,
    \ces_1_6_io_outs_up[58] ,
    \ces_1_6_io_outs_up[57] ,
    \ces_1_6_io_outs_up[56] ,
    \ces_1_6_io_outs_up[55] ,
    \ces_1_6_io_outs_up[54] ,
    \ces_1_6_io_outs_up[53] ,
    \ces_1_6_io_outs_up[52] ,
    \ces_1_6_io_outs_up[51] ,
    \ces_1_6_io_outs_up[50] ,
    \ces_1_6_io_outs_up[49] ,
    \ces_1_6_io_outs_up[48] ,
    \ces_1_6_io_outs_up[47] ,
    \ces_1_6_io_outs_up[46] ,
    \ces_1_6_io_outs_up[45] ,
    \ces_1_6_io_outs_up[44] ,
    \ces_1_6_io_outs_up[43] ,
    \ces_1_6_io_outs_up[42] ,
    \ces_1_6_io_outs_up[41] ,
    \ces_1_6_io_outs_up[40] ,
    \ces_1_6_io_outs_up[39] ,
    \ces_1_6_io_outs_up[38] ,
    \ces_1_6_io_outs_up[37] ,
    \ces_1_6_io_outs_up[36] ,
    \ces_1_6_io_outs_up[35] ,
    \ces_1_6_io_outs_up[34] ,
    \ces_1_6_io_outs_up[33] ,
    \ces_1_6_io_outs_up[32] ,
    \ces_1_6_io_outs_up[31] ,
    \ces_1_6_io_outs_up[30] ,
    \ces_1_6_io_outs_up[29] ,
    \ces_1_6_io_outs_up[28] ,
    \ces_1_6_io_outs_up[27] ,
    \ces_1_6_io_outs_up[26] ,
    \ces_1_6_io_outs_up[25] ,
    \ces_1_6_io_outs_up[24] ,
    \ces_1_6_io_outs_up[23] ,
    \ces_1_6_io_outs_up[22] ,
    \ces_1_6_io_outs_up[21] ,
    \ces_1_6_io_outs_up[20] ,
    \ces_1_6_io_outs_up[19] ,
    \ces_1_6_io_outs_up[18] ,
    \ces_1_6_io_outs_up[17] ,
    \ces_1_6_io_outs_up[16] ,
    \ces_1_6_io_outs_up[15] ,
    \ces_1_6_io_outs_up[14] ,
    \ces_1_6_io_outs_up[13] ,
    \ces_1_6_io_outs_up[12] ,
    \ces_1_6_io_outs_up[11] ,
    \ces_1_6_io_outs_up[10] ,
    \ces_1_6_io_outs_up[9] ,
    \ces_1_6_io_outs_up[8] ,
    \ces_1_6_io_outs_up[7] ,
    \ces_1_6_io_outs_up[6] ,
    \ces_1_6_io_outs_up[5] ,
    \ces_1_6_io_outs_up[4] ,
    \ces_1_6_io_outs_up[3] ,
    \ces_1_6_io_outs_up[2] ,
    \ces_1_6_io_outs_up[1] ,
    \ces_1_6_io_outs_up[0] }));
 Element ces_1_7 (.clock(clknet_3_2_0_clock),
    .io_lsbIns_1(ces_1_6_io_lsbOuts_1),
    .io_lsbIns_2(ces_1_6_io_lsbOuts_2),
    .io_lsbIns_3(ces_1_6_io_lsbOuts_3),
    .io_lsbIns_4(ces_1_6_io_lsbOuts_4),
    .io_lsbIns_5(ces_1_6_io_lsbOuts_5),
    .io_lsbIns_6(ces_1_6_io_lsbOuts_6),
    .io_lsbIns_7(ces_1_6_io_lsbOuts_7),
    .io_lsbOuts_0(ces_1_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_1_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_1_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_1_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_1_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_1_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_1_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_1_7_io_lsbOuts_7),
    .io_ins_down({\ces_1_7_io_ins_down[63] ,
    \ces_1_7_io_ins_down[62] ,
    \ces_1_7_io_ins_down[61] ,
    \ces_1_7_io_ins_down[60] ,
    \ces_1_7_io_ins_down[59] ,
    \ces_1_7_io_ins_down[58] ,
    \ces_1_7_io_ins_down[57] ,
    \ces_1_7_io_ins_down[56] ,
    \ces_1_7_io_ins_down[55] ,
    \ces_1_7_io_ins_down[54] ,
    \ces_1_7_io_ins_down[53] ,
    \ces_1_7_io_ins_down[52] ,
    \ces_1_7_io_ins_down[51] ,
    \ces_1_7_io_ins_down[50] ,
    \ces_1_7_io_ins_down[49] ,
    \ces_1_7_io_ins_down[48] ,
    \ces_1_7_io_ins_down[47] ,
    \ces_1_7_io_ins_down[46] ,
    \ces_1_7_io_ins_down[45] ,
    \ces_1_7_io_ins_down[44] ,
    \ces_1_7_io_ins_down[43] ,
    \ces_1_7_io_ins_down[42] ,
    \ces_1_7_io_ins_down[41] ,
    \ces_1_7_io_ins_down[40] ,
    \ces_1_7_io_ins_down[39] ,
    \ces_1_7_io_ins_down[38] ,
    \ces_1_7_io_ins_down[37] ,
    \ces_1_7_io_ins_down[36] ,
    \ces_1_7_io_ins_down[35] ,
    \ces_1_7_io_ins_down[34] ,
    \ces_1_7_io_ins_down[33] ,
    \ces_1_7_io_ins_down[32] ,
    \ces_1_7_io_ins_down[31] ,
    \ces_1_7_io_ins_down[30] ,
    \ces_1_7_io_ins_down[29] ,
    \ces_1_7_io_ins_down[28] ,
    \ces_1_7_io_ins_down[27] ,
    \ces_1_7_io_ins_down[26] ,
    \ces_1_7_io_ins_down[25] ,
    \ces_1_7_io_ins_down[24] ,
    \ces_1_7_io_ins_down[23] ,
    \ces_1_7_io_ins_down[22] ,
    \ces_1_7_io_ins_down[21] ,
    \ces_1_7_io_ins_down[20] ,
    \ces_1_7_io_ins_down[19] ,
    \ces_1_7_io_ins_down[18] ,
    \ces_1_7_io_ins_down[17] ,
    \ces_1_7_io_ins_down[16] ,
    \ces_1_7_io_ins_down[15] ,
    \ces_1_7_io_ins_down[14] ,
    \ces_1_7_io_ins_down[13] ,
    \ces_1_7_io_ins_down[12] ,
    \ces_1_7_io_ins_down[11] ,
    \ces_1_7_io_ins_down[10] ,
    \ces_1_7_io_ins_down[9] ,
    \ces_1_7_io_ins_down[8] ,
    \ces_1_7_io_ins_down[7] ,
    \ces_1_7_io_ins_down[6] ,
    \ces_1_7_io_ins_down[5] ,
    \ces_1_7_io_ins_down[4] ,
    \ces_1_7_io_ins_down[3] ,
    \ces_1_7_io_ins_down[2] ,
    \ces_1_7_io_ins_down[1] ,
    \ces_1_7_io_ins_down[0] }),
    .io_ins_left({net636,
    net635,
    net634,
    net633,
    net631,
    net630,
    net629,
    net628,
    net627,
    net626,
    net625,
    net624,
    net623,
    net622,
    net620,
    net619,
    net618,
    net617,
    net616,
    net615,
    net614,
    net613,
    net612,
    net611,
    net609,
    net608,
    net607,
    net606,
    net605,
    net604,
    net603,
    net602,
    net601,
    net600,
    net598,
    net597,
    net596,
    net595,
    net594,
    net593,
    net592,
    net591,
    net590,
    net589,
    net587,
    net586,
    net585,
    net584,
    net583,
    net582,
    net581,
    net580,
    net579,
    net578,
    net640,
    net639,
    net638,
    net637,
    net632,
    net621,
    net610,
    net599,
    net588,
    net577}),
    .io_ins_right({\ces_1_6_io_outs_right[63] ,
    \ces_1_6_io_outs_right[62] ,
    \ces_1_6_io_outs_right[61] ,
    \ces_1_6_io_outs_right[60] ,
    \ces_1_6_io_outs_right[59] ,
    \ces_1_6_io_outs_right[58] ,
    \ces_1_6_io_outs_right[57] ,
    \ces_1_6_io_outs_right[56] ,
    \ces_1_6_io_outs_right[55] ,
    \ces_1_6_io_outs_right[54] ,
    \ces_1_6_io_outs_right[53] ,
    \ces_1_6_io_outs_right[52] ,
    \ces_1_6_io_outs_right[51] ,
    \ces_1_6_io_outs_right[50] ,
    \ces_1_6_io_outs_right[49] ,
    \ces_1_6_io_outs_right[48] ,
    \ces_1_6_io_outs_right[47] ,
    \ces_1_6_io_outs_right[46] ,
    \ces_1_6_io_outs_right[45] ,
    \ces_1_6_io_outs_right[44] ,
    \ces_1_6_io_outs_right[43] ,
    \ces_1_6_io_outs_right[42] ,
    \ces_1_6_io_outs_right[41] ,
    \ces_1_6_io_outs_right[40] ,
    \ces_1_6_io_outs_right[39] ,
    \ces_1_6_io_outs_right[38] ,
    \ces_1_6_io_outs_right[37] ,
    \ces_1_6_io_outs_right[36] ,
    \ces_1_6_io_outs_right[35] ,
    \ces_1_6_io_outs_right[34] ,
    \ces_1_6_io_outs_right[33] ,
    \ces_1_6_io_outs_right[32] ,
    \ces_1_6_io_outs_right[31] ,
    \ces_1_6_io_outs_right[30] ,
    \ces_1_6_io_outs_right[29] ,
    \ces_1_6_io_outs_right[28] ,
    \ces_1_6_io_outs_right[27] ,
    \ces_1_6_io_outs_right[26] ,
    \ces_1_6_io_outs_right[25] ,
    \ces_1_6_io_outs_right[24] ,
    \ces_1_6_io_outs_right[23] ,
    \ces_1_6_io_outs_right[22] ,
    \ces_1_6_io_outs_right[21] ,
    \ces_1_6_io_outs_right[20] ,
    \ces_1_6_io_outs_right[19] ,
    \ces_1_6_io_outs_right[18] ,
    \ces_1_6_io_outs_right[17] ,
    \ces_1_6_io_outs_right[16] ,
    \ces_1_6_io_outs_right[15] ,
    \ces_1_6_io_outs_right[14] ,
    \ces_1_6_io_outs_right[13] ,
    \ces_1_6_io_outs_right[12] ,
    \ces_1_6_io_outs_right[11] ,
    \ces_1_6_io_outs_right[10] ,
    \ces_1_6_io_outs_right[9] ,
    \ces_1_6_io_outs_right[8] ,
    \ces_1_6_io_outs_right[7] ,
    \ces_1_6_io_outs_right[6] ,
    \ces_1_6_io_outs_right[5] ,
    \ces_1_6_io_outs_right[4] ,
    \ces_1_6_io_outs_right[3] ,
    \ces_1_6_io_outs_right[2] ,
    \ces_1_6_io_outs_right[1] ,
    \ces_1_6_io_outs_right[0] }),
    .io_ins_up({\ces_0_7_io_outs_up[63] ,
    \ces_0_7_io_outs_up[62] ,
    \ces_0_7_io_outs_up[61] ,
    \ces_0_7_io_outs_up[60] ,
    \ces_0_7_io_outs_up[59] ,
    \ces_0_7_io_outs_up[58] ,
    \ces_0_7_io_outs_up[57] ,
    \ces_0_7_io_outs_up[56] ,
    \ces_0_7_io_outs_up[55] ,
    \ces_0_7_io_outs_up[54] ,
    \ces_0_7_io_outs_up[53] ,
    \ces_0_7_io_outs_up[52] ,
    \ces_0_7_io_outs_up[51] ,
    \ces_0_7_io_outs_up[50] ,
    \ces_0_7_io_outs_up[49] ,
    \ces_0_7_io_outs_up[48] ,
    \ces_0_7_io_outs_up[47] ,
    \ces_0_7_io_outs_up[46] ,
    \ces_0_7_io_outs_up[45] ,
    \ces_0_7_io_outs_up[44] ,
    \ces_0_7_io_outs_up[43] ,
    \ces_0_7_io_outs_up[42] ,
    \ces_0_7_io_outs_up[41] ,
    \ces_0_7_io_outs_up[40] ,
    \ces_0_7_io_outs_up[39] ,
    \ces_0_7_io_outs_up[38] ,
    \ces_0_7_io_outs_up[37] ,
    \ces_0_7_io_outs_up[36] ,
    \ces_0_7_io_outs_up[35] ,
    \ces_0_7_io_outs_up[34] ,
    \ces_0_7_io_outs_up[33] ,
    \ces_0_7_io_outs_up[32] ,
    \ces_0_7_io_outs_up[31] ,
    \ces_0_7_io_outs_up[30] ,
    \ces_0_7_io_outs_up[29] ,
    \ces_0_7_io_outs_up[28] ,
    \ces_0_7_io_outs_up[27] ,
    \ces_0_7_io_outs_up[26] ,
    \ces_0_7_io_outs_up[25] ,
    \ces_0_7_io_outs_up[24] ,
    \ces_0_7_io_outs_up[23] ,
    \ces_0_7_io_outs_up[22] ,
    \ces_0_7_io_outs_up[21] ,
    \ces_0_7_io_outs_up[20] ,
    \ces_0_7_io_outs_up[19] ,
    \ces_0_7_io_outs_up[18] ,
    \ces_0_7_io_outs_up[17] ,
    \ces_0_7_io_outs_up[16] ,
    \ces_0_7_io_outs_up[15] ,
    \ces_0_7_io_outs_up[14] ,
    \ces_0_7_io_outs_up[13] ,
    \ces_0_7_io_outs_up[12] ,
    \ces_0_7_io_outs_up[11] ,
    \ces_0_7_io_outs_up[10] ,
    \ces_0_7_io_outs_up[9] ,
    \ces_0_7_io_outs_up[8] ,
    \ces_0_7_io_outs_up[7] ,
    \ces_0_7_io_outs_up[6] ,
    \ces_0_7_io_outs_up[5] ,
    \ces_0_7_io_outs_up[4] ,
    \ces_0_7_io_outs_up[3] ,
    \ces_0_7_io_outs_up[2] ,
    \ces_0_7_io_outs_up[1] ,
    \ces_0_7_io_outs_up[0] }),
    .io_outs_down({\ces_0_7_io_ins_down[63] ,
    \ces_0_7_io_ins_down[62] ,
    \ces_0_7_io_ins_down[61] ,
    \ces_0_7_io_ins_down[60] ,
    \ces_0_7_io_ins_down[59] ,
    \ces_0_7_io_ins_down[58] ,
    \ces_0_7_io_ins_down[57] ,
    \ces_0_7_io_ins_down[56] ,
    \ces_0_7_io_ins_down[55] ,
    \ces_0_7_io_ins_down[54] ,
    \ces_0_7_io_ins_down[53] ,
    \ces_0_7_io_ins_down[52] ,
    \ces_0_7_io_ins_down[51] ,
    \ces_0_7_io_ins_down[50] ,
    \ces_0_7_io_ins_down[49] ,
    \ces_0_7_io_ins_down[48] ,
    \ces_0_7_io_ins_down[47] ,
    \ces_0_7_io_ins_down[46] ,
    \ces_0_7_io_ins_down[45] ,
    \ces_0_7_io_ins_down[44] ,
    \ces_0_7_io_ins_down[43] ,
    \ces_0_7_io_ins_down[42] ,
    \ces_0_7_io_ins_down[41] ,
    \ces_0_7_io_ins_down[40] ,
    \ces_0_7_io_ins_down[39] ,
    \ces_0_7_io_ins_down[38] ,
    \ces_0_7_io_ins_down[37] ,
    \ces_0_7_io_ins_down[36] ,
    \ces_0_7_io_ins_down[35] ,
    \ces_0_7_io_ins_down[34] ,
    \ces_0_7_io_ins_down[33] ,
    \ces_0_7_io_ins_down[32] ,
    \ces_0_7_io_ins_down[31] ,
    \ces_0_7_io_ins_down[30] ,
    \ces_0_7_io_ins_down[29] ,
    \ces_0_7_io_ins_down[28] ,
    \ces_0_7_io_ins_down[27] ,
    \ces_0_7_io_ins_down[26] ,
    \ces_0_7_io_ins_down[25] ,
    \ces_0_7_io_ins_down[24] ,
    \ces_0_7_io_ins_down[23] ,
    \ces_0_7_io_ins_down[22] ,
    \ces_0_7_io_ins_down[21] ,
    \ces_0_7_io_ins_down[20] ,
    \ces_0_7_io_ins_down[19] ,
    \ces_0_7_io_ins_down[18] ,
    \ces_0_7_io_ins_down[17] ,
    \ces_0_7_io_ins_down[16] ,
    \ces_0_7_io_ins_down[15] ,
    \ces_0_7_io_ins_down[14] ,
    \ces_0_7_io_ins_down[13] ,
    \ces_0_7_io_ins_down[12] ,
    \ces_0_7_io_ins_down[11] ,
    \ces_0_7_io_ins_down[10] ,
    \ces_0_7_io_ins_down[9] ,
    \ces_0_7_io_ins_down[8] ,
    \ces_0_7_io_ins_down[7] ,
    \ces_0_7_io_ins_down[6] ,
    \ces_0_7_io_ins_down[5] ,
    \ces_0_7_io_ins_down[4] ,
    \ces_0_7_io_ins_down[3] ,
    \ces_0_7_io_ins_down[2] ,
    \ces_0_7_io_ins_down[1] ,
    \ces_0_7_io_ins_down[0] }),
    .io_outs_left({\ces_1_6_io_ins_left[63] ,
    \ces_1_6_io_ins_left[62] ,
    \ces_1_6_io_ins_left[61] ,
    \ces_1_6_io_ins_left[60] ,
    \ces_1_6_io_ins_left[59] ,
    \ces_1_6_io_ins_left[58] ,
    \ces_1_6_io_ins_left[57] ,
    \ces_1_6_io_ins_left[56] ,
    \ces_1_6_io_ins_left[55] ,
    \ces_1_6_io_ins_left[54] ,
    \ces_1_6_io_ins_left[53] ,
    \ces_1_6_io_ins_left[52] ,
    \ces_1_6_io_ins_left[51] ,
    \ces_1_6_io_ins_left[50] ,
    \ces_1_6_io_ins_left[49] ,
    \ces_1_6_io_ins_left[48] ,
    \ces_1_6_io_ins_left[47] ,
    \ces_1_6_io_ins_left[46] ,
    \ces_1_6_io_ins_left[45] ,
    \ces_1_6_io_ins_left[44] ,
    \ces_1_6_io_ins_left[43] ,
    \ces_1_6_io_ins_left[42] ,
    \ces_1_6_io_ins_left[41] ,
    \ces_1_6_io_ins_left[40] ,
    \ces_1_6_io_ins_left[39] ,
    \ces_1_6_io_ins_left[38] ,
    \ces_1_6_io_ins_left[37] ,
    \ces_1_6_io_ins_left[36] ,
    \ces_1_6_io_ins_left[35] ,
    \ces_1_6_io_ins_left[34] ,
    \ces_1_6_io_ins_left[33] ,
    \ces_1_6_io_ins_left[32] ,
    \ces_1_6_io_ins_left[31] ,
    \ces_1_6_io_ins_left[30] ,
    \ces_1_6_io_ins_left[29] ,
    \ces_1_6_io_ins_left[28] ,
    \ces_1_6_io_ins_left[27] ,
    \ces_1_6_io_ins_left[26] ,
    \ces_1_6_io_ins_left[25] ,
    \ces_1_6_io_ins_left[24] ,
    \ces_1_6_io_ins_left[23] ,
    \ces_1_6_io_ins_left[22] ,
    \ces_1_6_io_ins_left[21] ,
    \ces_1_6_io_ins_left[20] ,
    \ces_1_6_io_ins_left[19] ,
    \ces_1_6_io_ins_left[18] ,
    \ces_1_6_io_ins_left[17] ,
    \ces_1_6_io_ins_left[16] ,
    \ces_1_6_io_ins_left[15] ,
    \ces_1_6_io_ins_left[14] ,
    \ces_1_6_io_ins_left[13] ,
    \ces_1_6_io_ins_left[12] ,
    \ces_1_6_io_ins_left[11] ,
    \ces_1_6_io_ins_left[10] ,
    \ces_1_6_io_ins_left[9] ,
    \ces_1_6_io_ins_left[8] ,
    \ces_1_6_io_ins_left[7] ,
    \ces_1_6_io_ins_left[6] ,
    \ces_1_6_io_ins_left[5] ,
    \ces_1_6_io_ins_left[4] ,
    \ces_1_6_io_ins_left[3] ,
    \ces_1_6_io_ins_left[2] ,
    \ces_1_6_io_ins_left[1] ,
    \ces_1_6_io_ins_left[0] }),
    .io_outs_right({net3260,
    net3259,
    net3258,
    net3257,
    net3255,
    net3254,
    net3253,
    net3252,
    net3251,
    net3250,
    net3249,
    net3248,
    net3247,
    net3246,
    net3244,
    net3243,
    net3242,
    net3241,
    net3240,
    net3239,
    net3238,
    net3237,
    net3236,
    net3235,
    net3233,
    net3232,
    net3231,
    net3230,
    net3229,
    net3228,
    net3227,
    net3226,
    net3225,
    net3224,
    net3222,
    net3221,
    net3220,
    net3219,
    net3218,
    net3217,
    net3216,
    net3215,
    net3214,
    net3213,
    net3211,
    net3210,
    net3209,
    net3208,
    net3207,
    net3206,
    net3205,
    net3204,
    net3203,
    net3202,
    net3264,
    net3263,
    net3262,
    net3261,
    net3256,
    net3245,
    net3234,
    net3223,
    net3212,
    net3201}),
    .io_outs_up({\ces_1_7_io_outs_up[63] ,
    \ces_1_7_io_outs_up[62] ,
    \ces_1_7_io_outs_up[61] ,
    \ces_1_7_io_outs_up[60] ,
    \ces_1_7_io_outs_up[59] ,
    \ces_1_7_io_outs_up[58] ,
    \ces_1_7_io_outs_up[57] ,
    \ces_1_7_io_outs_up[56] ,
    \ces_1_7_io_outs_up[55] ,
    \ces_1_7_io_outs_up[54] ,
    \ces_1_7_io_outs_up[53] ,
    \ces_1_7_io_outs_up[52] ,
    \ces_1_7_io_outs_up[51] ,
    \ces_1_7_io_outs_up[50] ,
    \ces_1_7_io_outs_up[49] ,
    \ces_1_7_io_outs_up[48] ,
    \ces_1_7_io_outs_up[47] ,
    \ces_1_7_io_outs_up[46] ,
    \ces_1_7_io_outs_up[45] ,
    \ces_1_7_io_outs_up[44] ,
    \ces_1_7_io_outs_up[43] ,
    \ces_1_7_io_outs_up[42] ,
    \ces_1_7_io_outs_up[41] ,
    \ces_1_7_io_outs_up[40] ,
    \ces_1_7_io_outs_up[39] ,
    \ces_1_7_io_outs_up[38] ,
    \ces_1_7_io_outs_up[37] ,
    \ces_1_7_io_outs_up[36] ,
    \ces_1_7_io_outs_up[35] ,
    \ces_1_7_io_outs_up[34] ,
    \ces_1_7_io_outs_up[33] ,
    \ces_1_7_io_outs_up[32] ,
    \ces_1_7_io_outs_up[31] ,
    \ces_1_7_io_outs_up[30] ,
    \ces_1_7_io_outs_up[29] ,
    \ces_1_7_io_outs_up[28] ,
    \ces_1_7_io_outs_up[27] ,
    \ces_1_7_io_outs_up[26] ,
    \ces_1_7_io_outs_up[25] ,
    \ces_1_7_io_outs_up[24] ,
    \ces_1_7_io_outs_up[23] ,
    \ces_1_7_io_outs_up[22] ,
    \ces_1_7_io_outs_up[21] ,
    \ces_1_7_io_outs_up[20] ,
    \ces_1_7_io_outs_up[19] ,
    \ces_1_7_io_outs_up[18] ,
    \ces_1_7_io_outs_up[17] ,
    \ces_1_7_io_outs_up[16] ,
    \ces_1_7_io_outs_up[15] ,
    \ces_1_7_io_outs_up[14] ,
    \ces_1_7_io_outs_up[13] ,
    \ces_1_7_io_outs_up[12] ,
    \ces_1_7_io_outs_up[11] ,
    \ces_1_7_io_outs_up[10] ,
    \ces_1_7_io_outs_up[9] ,
    \ces_1_7_io_outs_up[8] ,
    \ces_1_7_io_outs_up[7] ,
    \ces_1_7_io_outs_up[6] ,
    \ces_1_7_io_outs_up[5] ,
    \ces_1_7_io_outs_up[4] ,
    \ces_1_7_io_outs_up[3] ,
    \ces_1_7_io_outs_up[2] ,
    \ces_1_7_io_outs_up[1] ,
    \ces_1_7_io_outs_up[0] }));
 Element ces_2_0 (.clock(clknet_3_1_0_clock),
    .io_lsbIns_1(net4175),
    .io_lsbIns_2(net4176),
    .io_lsbIns_3(net4177),
    .io_lsbIns_4(net4178),
    .io_lsbIns_5(net4179),
    .io_lsbIns_6(net4180),
    .io_lsbIns_7(net4181),
    .io_lsbOuts_0(ces_2_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_0_io_lsbOuts_7),
    .io_ins_down({\ces_2_0_io_ins_down[63] ,
    \ces_2_0_io_ins_down[62] ,
    \ces_2_0_io_ins_down[61] ,
    \ces_2_0_io_ins_down[60] ,
    \ces_2_0_io_ins_down[59] ,
    \ces_2_0_io_ins_down[58] ,
    \ces_2_0_io_ins_down[57] ,
    \ces_2_0_io_ins_down[56] ,
    \ces_2_0_io_ins_down[55] ,
    \ces_2_0_io_ins_down[54] ,
    \ces_2_0_io_ins_down[53] ,
    \ces_2_0_io_ins_down[52] ,
    \ces_2_0_io_ins_down[51] ,
    \ces_2_0_io_ins_down[50] ,
    \ces_2_0_io_ins_down[49] ,
    \ces_2_0_io_ins_down[48] ,
    \ces_2_0_io_ins_down[47] ,
    \ces_2_0_io_ins_down[46] ,
    \ces_2_0_io_ins_down[45] ,
    \ces_2_0_io_ins_down[44] ,
    \ces_2_0_io_ins_down[43] ,
    \ces_2_0_io_ins_down[42] ,
    \ces_2_0_io_ins_down[41] ,
    \ces_2_0_io_ins_down[40] ,
    \ces_2_0_io_ins_down[39] ,
    \ces_2_0_io_ins_down[38] ,
    \ces_2_0_io_ins_down[37] ,
    \ces_2_0_io_ins_down[36] ,
    \ces_2_0_io_ins_down[35] ,
    \ces_2_0_io_ins_down[34] ,
    \ces_2_0_io_ins_down[33] ,
    \ces_2_0_io_ins_down[32] ,
    \ces_2_0_io_ins_down[31] ,
    \ces_2_0_io_ins_down[30] ,
    \ces_2_0_io_ins_down[29] ,
    \ces_2_0_io_ins_down[28] ,
    \ces_2_0_io_ins_down[27] ,
    \ces_2_0_io_ins_down[26] ,
    \ces_2_0_io_ins_down[25] ,
    \ces_2_0_io_ins_down[24] ,
    \ces_2_0_io_ins_down[23] ,
    \ces_2_0_io_ins_down[22] ,
    \ces_2_0_io_ins_down[21] ,
    \ces_2_0_io_ins_down[20] ,
    \ces_2_0_io_ins_down[19] ,
    \ces_2_0_io_ins_down[18] ,
    \ces_2_0_io_ins_down[17] ,
    \ces_2_0_io_ins_down[16] ,
    \ces_2_0_io_ins_down[15] ,
    \ces_2_0_io_ins_down[14] ,
    \ces_2_0_io_ins_down[13] ,
    \ces_2_0_io_ins_down[12] ,
    \ces_2_0_io_ins_down[11] ,
    \ces_2_0_io_ins_down[10] ,
    \ces_2_0_io_ins_down[9] ,
    \ces_2_0_io_ins_down[8] ,
    \ces_2_0_io_ins_down[7] ,
    \ces_2_0_io_ins_down[6] ,
    \ces_2_0_io_ins_down[5] ,
    \ces_2_0_io_ins_down[4] ,
    \ces_2_0_io_ins_down[3] ,
    \ces_2_0_io_ins_down[2] ,
    \ces_2_0_io_ins_down[1] ,
    \ces_2_0_io_ins_down[0] }),
    .io_ins_left({\ces_2_0_io_ins_left[63] ,
    \ces_2_0_io_ins_left[62] ,
    \ces_2_0_io_ins_left[61] ,
    \ces_2_0_io_ins_left[60] ,
    \ces_2_0_io_ins_left[59] ,
    \ces_2_0_io_ins_left[58] ,
    \ces_2_0_io_ins_left[57] ,
    \ces_2_0_io_ins_left[56] ,
    \ces_2_0_io_ins_left[55] ,
    \ces_2_0_io_ins_left[54] ,
    \ces_2_0_io_ins_left[53] ,
    \ces_2_0_io_ins_left[52] ,
    \ces_2_0_io_ins_left[51] ,
    \ces_2_0_io_ins_left[50] ,
    \ces_2_0_io_ins_left[49] ,
    \ces_2_0_io_ins_left[48] ,
    \ces_2_0_io_ins_left[47] ,
    \ces_2_0_io_ins_left[46] ,
    \ces_2_0_io_ins_left[45] ,
    \ces_2_0_io_ins_left[44] ,
    \ces_2_0_io_ins_left[43] ,
    \ces_2_0_io_ins_left[42] ,
    \ces_2_0_io_ins_left[41] ,
    \ces_2_0_io_ins_left[40] ,
    \ces_2_0_io_ins_left[39] ,
    \ces_2_0_io_ins_left[38] ,
    \ces_2_0_io_ins_left[37] ,
    \ces_2_0_io_ins_left[36] ,
    \ces_2_0_io_ins_left[35] ,
    \ces_2_0_io_ins_left[34] ,
    \ces_2_0_io_ins_left[33] ,
    \ces_2_0_io_ins_left[32] ,
    \ces_2_0_io_ins_left[31] ,
    \ces_2_0_io_ins_left[30] ,
    \ces_2_0_io_ins_left[29] ,
    \ces_2_0_io_ins_left[28] ,
    \ces_2_0_io_ins_left[27] ,
    \ces_2_0_io_ins_left[26] ,
    \ces_2_0_io_ins_left[25] ,
    \ces_2_0_io_ins_left[24] ,
    \ces_2_0_io_ins_left[23] ,
    \ces_2_0_io_ins_left[22] ,
    \ces_2_0_io_ins_left[21] ,
    \ces_2_0_io_ins_left[20] ,
    \ces_2_0_io_ins_left[19] ,
    \ces_2_0_io_ins_left[18] ,
    \ces_2_0_io_ins_left[17] ,
    \ces_2_0_io_ins_left[16] ,
    \ces_2_0_io_ins_left[15] ,
    \ces_2_0_io_ins_left[14] ,
    \ces_2_0_io_ins_left[13] ,
    \ces_2_0_io_ins_left[12] ,
    \ces_2_0_io_ins_left[11] ,
    \ces_2_0_io_ins_left[10] ,
    \ces_2_0_io_ins_left[9] ,
    \ces_2_0_io_ins_left[8] ,
    \ces_2_0_io_ins_left[7] ,
    \ces_2_0_io_ins_left[6] ,
    \ces_2_0_io_ins_left[5] ,
    \ces_2_0_io_ins_left[4] ,
    \ces_2_0_io_ins_left[3] ,
    \ces_2_0_io_ins_left[2] ,
    \ces_2_0_io_ins_left[1] ,
    \ces_2_0_io_ins_left[0] }),
    .io_ins_right({net1212,
    net1211,
    net1210,
    net1209,
    net1207,
    net1206,
    net1205,
    net1204,
    net1203,
    net1202,
    net1201,
    net1200,
    net1199,
    net1198,
    net1196,
    net1195,
    net1194,
    net1193,
    net1192,
    net1191,
    net1190,
    net1189,
    net1188,
    net1187,
    net1185,
    net1184,
    net1183,
    net1182,
    net1181,
    net1180,
    net1179,
    net1178,
    net1177,
    net1176,
    net1174,
    net1173,
    net1172,
    net1171,
    net1170,
    net1169,
    net1168,
    net1167,
    net1166,
    net1165,
    net1163,
    net1162,
    net1161,
    net1160,
    net1159,
    net1158,
    net1157,
    net1156,
    net1155,
    net1154,
    net1216,
    net1215,
    net1214,
    net1213,
    net1208,
    net1197,
    net1186,
    net1175,
    net1164,
    net1153}),
    .io_ins_up({\ces_1_0_io_outs_up[63] ,
    \ces_1_0_io_outs_up[62] ,
    \ces_1_0_io_outs_up[61] ,
    \ces_1_0_io_outs_up[60] ,
    \ces_1_0_io_outs_up[59] ,
    \ces_1_0_io_outs_up[58] ,
    \ces_1_0_io_outs_up[57] ,
    \ces_1_0_io_outs_up[56] ,
    \ces_1_0_io_outs_up[55] ,
    \ces_1_0_io_outs_up[54] ,
    \ces_1_0_io_outs_up[53] ,
    \ces_1_0_io_outs_up[52] ,
    \ces_1_0_io_outs_up[51] ,
    \ces_1_0_io_outs_up[50] ,
    \ces_1_0_io_outs_up[49] ,
    \ces_1_0_io_outs_up[48] ,
    \ces_1_0_io_outs_up[47] ,
    \ces_1_0_io_outs_up[46] ,
    \ces_1_0_io_outs_up[45] ,
    \ces_1_0_io_outs_up[44] ,
    \ces_1_0_io_outs_up[43] ,
    \ces_1_0_io_outs_up[42] ,
    \ces_1_0_io_outs_up[41] ,
    \ces_1_0_io_outs_up[40] ,
    \ces_1_0_io_outs_up[39] ,
    \ces_1_0_io_outs_up[38] ,
    \ces_1_0_io_outs_up[37] ,
    \ces_1_0_io_outs_up[36] ,
    \ces_1_0_io_outs_up[35] ,
    \ces_1_0_io_outs_up[34] ,
    \ces_1_0_io_outs_up[33] ,
    \ces_1_0_io_outs_up[32] ,
    \ces_1_0_io_outs_up[31] ,
    \ces_1_0_io_outs_up[30] ,
    \ces_1_0_io_outs_up[29] ,
    \ces_1_0_io_outs_up[28] ,
    \ces_1_0_io_outs_up[27] ,
    \ces_1_0_io_outs_up[26] ,
    \ces_1_0_io_outs_up[25] ,
    \ces_1_0_io_outs_up[24] ,
    \ces_1_0_io_outs_up[23] ,
    \ces_1_0_io_outs_up[22] ,
    \ces_1_0_io_outs_up[21] ,
    \ces_1_0_io_outs_up[20] ,
    \ces_1_0_io_outs_up[19] ,
    \ces_1_0_io_outs_up[18] ,
    \ces_1_0_io_outs_up[17] ,
    \ces_1_0_io_outs_up[16] ,
    \ces_1_0_io_outs_up[15] ,
    \ces_1_0_io_outs_up[14] ,
    \ces_1_0_io_outs_up[13] ,
    \ces_1_0_io_outs_up[12] ,
    \ces_1_0_io_outs_up[11] ,
    \ces_1_0_io_outs_up[10] ,
    \ces_1_0_io_outs_up[9] ,
    \ces_1_0_io_outs_up[8] ,
    \ces_1_0_io_outs_up[7] ,
    \ces_1_0_io_outs_up[6] ,
    \ces_1_0_io_outs_up[5] ,
    \ces_1_0_io_outs_up[4] ,
    \ces_1_0_io_outs_up[3] ,
    \ces_1_0_io_outs_up[2] ,
    \ces_1_0_io_outs_up[1] ,
    \ces_1_0_io_outs_up[0] }),
    .io_outs_down({\ces_1_0_io_ins_down[63] ,
    \ces_1_0_io_ins_down[62] ,
    \ces_1_0_io_ins_down[61] ,
    \ces_1_0_io_ins_down[60] ,
    \ces_1_0_io_ins_down[59] ,
    \ces_1_0_io_ins_down[58] ,
    \ces_1_0_io_ins_down[57] ,
    \ces_1_0_io_ins_down[56] ,
    \ces_1_0_io_ins_down[55] ,
    \ces_1_0_io_ins_down[54] ,
    \ces_1_0_io_ins_down[53] ,
    \ces_1_0_io_ins_down[52] ,
    \ces_1_0_io_ins_down[51] ,
    \ces_1_0_io_ins_down[50] ,
    \ces_1_0_io_ins_down[49] ,
    \ces_1_0_io_ins_down[48] ,
    \ces_1_0_io_ins_down[47] ,
    \ces_1_0_io_ins_down[46] ,
    \ces_1_0_io_ins_down[45] ,
    \ces_1_0_io_ins_down[44] ,
    \ces_1_0_io_ins_down[43] ,
    \ces_1_0_io_ins_down[42] ,
    \ces_1_0_io_ins_down[41] ,
    \ces_1_0_io_ins_down[40] ,
    \ces_1_0_io_ins_down[39] ,
    \ces_1_0_io_ins_down[38] ,
    \ces_1_0_io_ins_down[37] ,
    \ces_1_0_io_ins_down[36] ,
    \ces_1_0_io_ins_down[35] ,
    \ces_1_0_io_ins_down[34] ,
    \ces_1_0_io_ins_down[33] ,
    \ces_1_0_io_ins_down[32] ,
    \ces_1_0_io_ins_down[31] ,
    \ces_1_0_io_ins_down[30] ,
    \ces_1_0_io_ins_down[29] ,
    \ces_1_0_io_ins_down[28] ,
    \ces_1_0_io_ins_down[27] ,
    \ces_1_0_io_ins_down[26] ,
    \ces_1_0_io_ins_down[25] ,
    \ces_1_0_io_ins_down[24] ,
    \ces_1_0_io_ins_down[23] ,
    \ces_1_0_io_ins_down[22] ,
    \ces_1_0_io_ins_down[21] ,
    \ces_1_0_io_ins_down[20] ,
    \ces_1_0_io_ins_down[19] ,
    \ces_1_0_io_ins_down[18] ,
    \ces_1_0_io_ins_down[17] ,
    \ces_1_0_io_ins_down[16] ,
    \ces_1_0_io_ins_down[15] ,
    \ces_1_0_io_ins_down[14] ,
    \ces_1_0_io_ins_down[13] ,
    \ces_1_0_io_ins_down[12] ,
    \ces_1_0_io_ins_down[11] ,
    \ces_1_0_io_ins_down[10] ,
    \ces_1_0_io_ins_down[9] ,
    \ces_1_0_io_ins_down[8] ,
    \ces_1_0_io_ins_down[7] ,
    \ces_1_0_io_ins_down[6] ,
    \ces_1_0_io_ins_down[5] ,
    \ces_1_0_io_ins_down[4] ,
    \ces_1_0_io_ins_down[3] ,
    \ces_1_0_io_ins_down[2] ,
    \ces_1_0_io_ins_down[1] ,
    \ces_1_0_io_ins_down[0] }),
    .io_outs_left({net2812,
    net2811,
    net2810,
    net2809,
    net2807,
    net2806,
    net2805,
    net2804,
    net2803,
    net2802,
    net2801,
    net2800,
    net2799,
    net2798,
    net2796,
    net2795,
    net2794,
    net2793,
    net2792,
    net2791,
    net2790,
    net2789,
    net2788,
    net2787,
    net2785,
    net2784,
    net2783,
    net2782,
    net2781,
    net2780,
    net2779,
    net2778,
    net2777,
    net2776,
    net2774,
    net2773,
    net2772,
    net2771,
    net2770,
    net2769,
    net2768,
    net2767,
    net2766,
    net2765,
    net2763,
    net2762,
    net2761,
    net2760,
    net2759,
    net2758,
    net2757,
    net2756,
    net2755,
    net2754,
    net2816,
    net2815,
    net2814,
    net2813,
    net2808,
    net2797,
    net2786,
    net2775,
    net2764,
    net2753}),
    .io_outs_right({\ces_2_0_io_outs_right[63] ,
    \ces_2_0_io_outs_right[62] ,
    \ces_2_0_io_outs_right[61] ,
    \ces_2_0_io_outs_right[60] ,
    \ces_2_0_io_outs_right[59] ,
    \ces_2_0_io_outs_right[58] ,
    \ces_2_0_io_outs_right[57] ,
    \ces_2_0_io_outs_right[56] ,
    \ces_2_0_io_outs_right[55] ,
    \ces_2_0_io_outs_right[54] ,
    \ces_2_0_io_outs_right[53] ,
    \ces_2_0_io_outs_right[52] ,
    \ces_2_0_io_outs_right[51] ,
    \ces_2_0_io_outs_right[50] ,
    \ces_2_0_io_outs_right[49] ,
    \ces_2_0_io_outs_right[48] ,
    \ces_2_0_io_outs_right[47] ,
    \ces_2_0_io_outs_right[46] ,
    \ces_2_0_io_outs_right[45] ,
    \ces_2_0_io_outs_right[44] ,
    \ces_2_0_io_outs_right[43] ,
    \ces_2_0_io_outs_right[42] ,
    \ces_2_0_io_outs_right[41] ,
    \ces_2_0_io_outs_right[40] ,
    \ces_2_0_io_outs_right[39] ,
    \ces_2_0_io_outs_right[38] ,
    \ces_2_0_io_outs_right[37] ,
    \ces_2_0_io_outs_right[36] ,
    \ces_2_0_io_outs_right[35] ,
    \ces_2_0_io_outs_right[34] ,
    \ces_2_0_io_outs_right[33] ,
    \ces_2_0_io_outs_right[32] ,
    \ces_2_0_io_outs_right[31] ,
    \ces_2_0_io_outs_right[30] ,
    \ces_2_0_io_outs_right[29] ,
    \ces_2_0_io_outs_right[28] ,
    \ces_2_0_io_outs_right[27] ,
    \ces_2_0_io_outs_right[26] ,
    \ces_2_0_io_outs_right[25] ,
    \ces_2_0_io_outs_right[24] ,
    \ces_2_0_io_outs_right[23] ,
    \ces_2_0_io_outs_right[22] ,
    \ces_2_0_io_outs_right[21] ,
    \ces_2_0_io_outs_right[20] ,
    \ces_2_0_io_outs_right[19] ,
    \ces_2_0_io_outs_right[18] ,
    \ces_2_0_io_outs_right[17] ,
    \ces_2_0_io_outs_right[16] ,
    \ces_2_0_io_outs_right[15] ,
    \ces_2_0_io_outs_right[14] ,
    \ces_2_0_io_outs_right[13] ,
    \ces_2_0_io_outs_right[12] ,
    \ces_2_0_io_outs_right[11] ,
    \ces_2_0_io_outs_right[10] ,
    \ces_2_0_io_outs_right[9] ,
    \ces_2_0_io_outs_right[8] ,
    \ces_2_0_io_outs_right[7] ,
    \ces_2_0_io_outs_right[6] ,
    \ces_2_0_io_outs_right[5] ,
    \ces_2_0_io_outs_right[4] ,
    \ces_2_0_io_outs_right[3] ,
    \ces_2_0_io_outs_right[2] ,
    \ces_2_0_io_outs_right[1] ,
    \ces_2_0_io_outs_right[0] }),
    .io_outs_up({\ces_2_0_io_outs_up[63] ,
    \ces_2_0_io_outs_up[62] ,
    \ces_2_0_io_outs_up[61] ,
    \ces_2_0_io_outs_up[60] ,
    \ces_2_0_io_outs_up[59] ,
    \ces_2_0_io_outs_up[58] ,
    \ces_2_0_io_outs_up[57] ,
    \ces_2_0_io_outs_up[56] ,
    \ces_2_0_io_outs_up[55] ,
    \ces_2_0_io_outs_up[54] ,
    \ces_2_0_io_outs_up[53] ,
    \ces_2_0_io_outs_up[52] ,
    \ces_2_0_io_outs_up[51] ,
    \ces_2_0_io_outs_up[50] ,
    \ces_2_0_io_outs_up[49] ,
    \ces_2_0_io_outs_up[48] ,
    \ces_2_0_io_outs_up[47] ,
    \ces_2_0_io_outs_up[46] ,
    \ces_2_0_io_outs_up[45] ,
    \ces_2_0_io_outs_up[44] ,
    \ces_2_0_io_outs_up[43] ,
    \ces_2_0_io_outs_up[42] ,
    \ces_2_0_io_outs_up[41] ,
    \ces_2_0_io_outs_up[40] ,
    \ces_2_0_io_outs_up[39] ,
    \ces_2_0_io_outs_up[38] ,
    \ces_2_0_io_outs_up[37] ,
    \ces_2_0_io_outs_up[36] ,
    \ces_2_0_io_outs_up[35] ,
    \ces_2_0_io_outs_up[34] ,
    \ces_2_0_io_outs_up[33] ,
    \ces_2_0_io_outs_up[32] ,
    \ces_2_0_io_outs_up[31] ,
    \ces_2_0_io_outs_up[30] ,
    \ces_2_0_io_outs_up[29] ,
    \ces_2_0_io_outs_up[28] ,
    \ces_2_0_io_outs_up[27] ,
    \ces_2_0_io_outs_up[26] ,
    \ces_2_0_io_outs_up[25] ,
    \ces_2_0_io_outs_up[24] ,
    \ces_2_0_io_outs_up[23] ,
    \ces_2_0_io_outs_up[22] ,
    \ces_2_0_io_outs_up[21] ,
    \ces_2_0_io_outs_up[20] ,
    \ces_2_0_io_outs_up[19] ,
    \ces_2_0_io_outs_up[18] ,
    \ces_2_0_io_outs_up[17] ,
    \ces_2_0_io_outs_up[16] ,
    \ces_2_0_io_outs_up[15] ,
    \ces_2_0_io_outs_up[14] ,
    \ces_2_0_io_outs_up[13] ,
    \ces_2_0_io_outs_up[12] ,
    \ces_2_0_io_outs_up[11] ,
    \ces_2_0_io_outs_up[10] ,
    \ces_2_0_io_outs_up[9] ,
    \ces_2_0_io_outs_up[8] ,
    \ces_2_0_io_outs_up[7] ,
    \ces_2_0_io_outs_up[6] ,
    \ces_2_0_io_outs_up[5] ,
    \ces_2_0_io_outs_up[4] ,
    \ces_2_0_io_outs_up[3] ,
    \ces_2_0_io_outs_up[2] ,
    \ces_2_0_io_outs_up[1] ,
    \ces_2_0_io_outs_up[0] }));
 Element ces_2_1 (.clock(clknet_3_1_0_clock),
    .io_lsbIns_1(ces_2_0_io_lsbOuts_1),
    .io_lsbIns_2(ces_2_0_io_lsbOuts_2),
    .io_lsbIns_3(ces_2_0_io_lsbOuts_3),
    .io_lsbIns_4(ces_2_0_io_lsbOuts_4),
    .io_lsbIns_5(ces_2_0_io_lsbOuts_5),
    .io_lsbIns_6(ces_2_0_io_lsbOuts_6),
    .io_lsbIns_7(ces_2_0_io_lsbOuts_7),
    .io_lsbOuts_0(ces_2_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_1_io_lsbOuts_7),
    .io_ins_down({\ces_2_1_io_ins_down[63] ,
    \ces_2_1_io_ins_down[62] ,
    \ces_2_1_io_ins_down[61] ,
    \ces_2_1_io_ins_down[60] ,
    \ces_2_1_io_ins_down[59] ,
    \ces_2_1_io_ins_down[58] ,
    \ces_2_1_io_ins_down[57] ,
    \ces_2_1_io_ins_down[56] ,
    \ces_2_1_io_ins_down[55] ,
    \ces_2_1_io_ins_down[54] ,
    \ces_2_1_io_ins_down[53] ,
    \ces_2_1_io_ins_down[52] ,
    \ces_2_1_io_ins_down[51] ,
    \ces_2_1_io_ins_down[50] ,
    \ces_2_1_io_ins_down[49] ,
    \ces_2_1_io_ins_down[48] ,
    \ces_2_1_io_ins_down[47] ,
    \ces_2_1_io_ins_down[46] ,
    \ces_2_1_io_ins_down[45] ,
    \ces_2_1_io_ins_down[44] ,
    \ces_2_1_io_ins_down[43] ,
    \ces_2_1_io_ins_down[42] ,
    \ces_2_1_io_ins_down[41] ,
    \ces_2_1_io_ins_down[40] ,
    \ces_2_1_io_ins_down[39] ,
    \ces_2_1_io_ins_down[38] ,
    \ces_2_1_io_ins_down[37] ,
    \ces_2_1_io_ins_down[36] ,
    \ces_2_1_io_ins_down[35] ,
    \ces_2_1_io_ins_down[34] ,
    \ces_2_1_io_ins_down[33] ,
    \ces_2_1_io_ins_down[32] ,
    \ces_2_1_io_ins_down[31] ,
    \ces_2_1_io_ins_down[30] ,
    \ces_2_1_io_ins_down[29] ,
    \ces_2_1_io_ins_down[28] ,
    \ces_2_1_io_ins_down[27] ,
    \ces_2_1_io_ins_down[26] ,
    \ces_2_1_io_ins_down[25] ,
    \ces_2_1_io_ins_down[24] ,
    \ces_2_1_io_ins_down[23] ,
    \ces_2_1_io_ins_down[22] ,
    \ces_2_1_io_ins_down[21] ,
    \ces_2_1_io_ins_down[20] ,
    \ces_2_1_io_ins_down[19] ,
    \ces_2_1_io_ins_down[18] ,
    \ces_2_1_io_ins_down[17] ,
    \ces_2_1_io_ins_down[16] ,
    \ces_2_1_io_ins_down[15] ,
    \ces_2_1_io_ins_down[14] ,
    \ces_2_1_io_ins_down[13] ,
    \ces_2_1_io_ins_down[12] ,
    \ces_2_1_io_ins_down[11] ,
    \ces_2_1_io_ins_down[10] ,
    \ces_2_1_io_ins_down[9] ,
    \ces_2_1_io_ins_down[8] ,
    \ces_2_1_io_ins_down[7] ,
    \ces_2_1_io_ins_down[6] ,
    \ces_2_1_io_ins_down[5] ,
    \ces_2_1_io_ins_down[4] ,
    \ces_2_1_io_ins_down[3] ,
    \ces_2_1_io_ins_down[2] ,
    \ces_2_1_io_ins_down[1] ,
    \ces_2_1_io_ins_down[0] }),
    .io_ins_left({\ces_2_1_io_ins_left[63] ,
    \ces_2_1_io_ins_left[62] ,
    \ces_2_1_io_ins_left[61] ,
    \ces_2_1_io_ins_left[60] ,
    \ces_2_1_io_ins_left[59] ,
    \ces_2_1_io_ins_left[58] ,
    \ces_2_1_io_ins_left[57] ,
    \ces_2_1_io_ins_left[56] ,
    \ces_2_1_io_ins_left[55] ,
    \ces_2_1_io_ins_left[54] ,
    \ces_2_1_io_ins_left[53] ,
    \ces_2_1_io_ins_left[52] ,
    \ces_2_1_io_ins_left[51] ,
    \ces_2_1_io_ins_left[50] ,
    \ces_2_1_io_ins_left[49] ,
    \ces_2_1_io_ins_left[48] ,
    \ces_2_1_io_ins_left[47] ,
    \ces_2_1_io_ins_left[46] ,
    \ces_2_1_io_ins_left[45] ,
    \ces_2_1_io_ins_left[44] ,
    \ces_2_1_io_ins_left[43] ,
    \ces_2_1_io_ins_left[42] ,
    \ces_2_1_io_ins_left[41] ,
    \ces_2_1_io_ins_left[40] ,
    \ces_2_1_io_ins_left[39] ,
    \ces_2_1_io_ins_left[38] ,
    \ces_2_1_io_ins_left[37] ,
    \ces_2_1_io_ins_left[36] ,
    \ces_2_1_io_ins_left[35] ,
    \ces_2_1_io_ins_left[34] ,
    \ces_2_1_io_ins_left[33] ,
    \ces_2_1_io_ins_left[32] ,
    \ces_2_1_io_ins_left[31] ,
    \ces_2_1_io_ins_left[30] ,
    \ces_2_1_io_ins_left[29] ,
    \ces_2_1_io_ins_left[28] ,
    \ces_2_1_io_ins_left[27] ,
    \ces_2_1_io_ins_left[26] ,
    \ces_2_1_io_ins_left[25] ,
    \ces_2_1_io_ins_left[24] ,
    \ces_2_1_io_ins_left[23] ,
    \ces_2_1_io_ins_left[22] ,
    \ces_2_1_io_ins_left[21] ,
    \ces_2_1_io_ins_left[20] ,
    \ces_2_1_io_ins_left[19] ,
    \ces_2_1_io_ins_left[18] ,
    \ces_2_1_io_ins_left[17] ,
    \ces_2_1_io_ins_left[16] ,
    \ces_2_1_io_ins_left[15] ,
    \ces_2_1_io_ins_left[14] ,
    \ces_2_1_io_ins_left[13] ,
    \ces_2_1_io_ins_left[12] ,
    \ces_2_1_io_ins_left[11] ,
    \ces_2_1_io_ins_left[10] ,
    \ces_2_1_io_ins_left[9] ,
    \ces_2_1_io_ins_left[8] ,
    \ces_2_1_io_ins_left[7] ,
    \ces_2_1_io_ins_left[6] ,
    \ces_2_1_io_ins_left[5] ,
    \ces_2_1_io_ins_left[4] ,
    \ces_2_1_io_ins_left[3] ,
    \ces_2_1_io_ins_left[2] ,
    \ces_2_1_io_ins_left[1] ,
    \ces_2_1_io_ins_left[0] }),
    .io_ins_right({\ces_2_0_io_outs_right[63] ,
    \ces_2_0_io_outs_right[62] ,
    \ces_2_0_io_outs_right[61] ,
    \ces_2_0_io_outs_right[60] ,
    \ces_2_0_io_outs_right[59] ,
    \ces_2_0_io_outs_right[58] ,
    \ces_2_0_io_outs_right[57] ,
    \ces_2_0_io_outs_right[56] ,
    \ces_2_0_io_outs_right[55] ,
    \ces_2_0_io_outs_right[54] ,
    \ces_2_0_io_outs_right[53] ,
    \ces_2_0_io_outs_right[52] ,
    \ces_2_0_io_outs_right[51] ,
    \ces_2_0_io_outs_right[50] ,
    \ces_2_0_io_outs_right[49] ,
    \ces_2_0_io_outs_right[48] ,
    \ces_2_0_io_outs_right[47] ,
    \ces_2_0_io_outs_right[46] ,
    \ces_2_0_io_outs_right[45] ,
    \ces_2_0_io_outs_right[44] ,
    \ces_2_0_io_outs_right[43] ,
    \ces_2_0_io_outs_right[42] ,
    \ces_2_0_io_outs_right[41] ,
    \ces_2_0_io_outs_right[40] ,
    \ces_2_0_io_outs_right[39] ,
    \ces_2_0_io_outs_right[38] ,
    \ces_2_0_io_outs_right[37] ,
    \ces_2_0_io_outs_right[36] ,
    \ces_2_0_io_outs_right[35] ,
    \ces_2_0_io_outs_right[34] ,
    \ces_2_0_io_outs_right[33] ,
    \ces_2_0_io_outs_right[32] ,
    \ces_2_0_io_outs_right[31] ,
    \ces_2_0_io_outs_right[30] ,
    \ces_2_0_io_outs_right[29] ,
    \ces_2_0_io_outs_right[28] ,
    \ces_2_0_io_outs_right[27] ,
    \ces_2_0_io_outs_right[26] ,
    \ces_2_0_io_outs_right[25] ,
    \ces_2_0_io_outs_right[24] ,
    \ces_2_0_io_outs_right[23] ,
    \ces_2_0_io_outs_right[22] ,
    \ces_2_0_io_outs_right[21] ,
    \ces_2_0_io_outs_right[20] ,
    \ces_2_0_io_outs_right[19] ,
    \ces_2_0_io_outs_right[18] ,
    \ces_2_0_io_outs_right[17] ,
    \ces_2_0_io_outs_right[16] ,
    \ces_2_0_io_outs_right[15] ,
    \ces_2_0_io_outs_right[14] ,
    \ces_2_0_io_outs_right[13] ,
    \ces_2_0_io_outs_right[12] ,
    \ces_2_0_io_outs_right[11] ,
    \ces_2_0_io_outs_right[10] ,
    \ces_2_0_io_outs_right[9] ,
    \ces_2_0_io_outs_right[8] ,
    \ces_2_0_io_outs_right[7] ,
    \ces_2_0_io_outs_right[6] ,
    \ces_2_0_io_outs_right[5] ,
    \ces_2_0_io_outs_right[4] ,
    \ces_2_0_io_outs_right[3] ,
    \ces_2_0_io_outs_right[2] ,
    \ces_2_0_io_outs_right[1] ,
    \ces_2_0_io_outs_right[0] }),
    .io_ins_up({\ces_1_1_io_outs_up[63] ,
    \ces_1_1_io_outs_up[62] ,
    \ces_1_1_io_outs_up[61] ,
    \ces_1_1_io_outs_up[60] ,
    \ces_1_1_io_outs_up[59] ,
    \ces_1_1_io_outs_up[58] ,
    \ces_1_1_io_outs_up[57] ,
    \ces_1_1_io_outs_up[56] ,
    \ces_1_1_io_outs_up[55] ,
    \ces_1_1_io_outs_up[54] ,
    \ces_1_1_io_outs_up[53] ,
    \ces_1_1_io_outs_up[52] ,
    \ces_1_1_io_outs_up[51] ,
    \ces_1_1_io_outs_up[50] ,
    \ces_1_1_io_outs_up[49] ,
    \ces_1_1_io_outs_up[48] ,
    \ces_1_1_io_outs_up[47] ,
    \ces_1_1_io_outs_up[46] ,
    \ces_1_1_io_outs_up[45] ,
    \ces_1_1_io_outs_up[44] ,
    \ces_1_1_io_outs_up[43] ,
    \ces_1_1_io_outs_up[42] ,
    \ces_1_1_io_outs_up[41] ,
    \ces_1_1_io_outs_up[40] ,
    \ces_1_1_io_outs_up[39] ,
    \ces_1_1_io_outs_up[38] ,
    \ces_1_1_io_outs_up[37] ,
    \ces_1_1_io_outs_up[36] ,
    \ces_1_1_io_outs_up[35] ,
    \ces_1_1_io_outs_up[34] ,
    \ces_1_1_io_outs_up[33] ,
    \ces_1_1_io_outs_up[32] ,
    \ces_1_1_io_outs_up[31] ,
    \ces_1_1_io_outs_up[30] ,
    \ces_1_1_io_outs_up[29] ,
    \ces_1_1_io_outs_up[28] ,
    \ces_1_1_io_outs_up[27] ,
    \ces_1_1_io_outs_up[26] ,
    \ces_1_1_io_outs_up[25] ,
    \ces_1_1_io_outs_up[24] ,
    \ces_1_1_io_outs_up[23] ,
    \ces_1_1_io_outs_up[22] ,
    \ces_1_1_io_outs_up[21] ,
    \ces_1_1_io_outs_up[20] ,
    \ces_1_1_io_outs_up[19] ,
    \ces_1_1_io_outs_up[18] ,
    \ces_1_1_io_outs_up[17] ,
    \ces_1_1_io_outs_up[16] ,
    \ces_1_1_io_outs_up[15] ,
    \ces_1_1_io_outs_up[14] ,
    \ces_1_1_io_outs_up[13] ,
    \ces_1_1_io_outs_up[12] ,
    \ces_1_1_io_outs_up[11] ,
    \ces_1_1_io_outs_up[10] ,
    \ces_1_1_io_outs_up[9] ,
    \ces_1_1_io_outs_up[8] ,
    \ces_1_1_io_outs_up[7] ,
    \ces_1_1_io_outs_up[6] ,
    \ces_1_1_io_outs_up[5] ,
    \ces_1_1_io_outs_up[4] ,
    \ces_1_1_io_outs_up[3] ,
    \ces_1_1_io_outs_up[2] ,
    \ces_1_1_io_outs_up[1] ,
    \ces_1_1_io_outs_up[0] }),
    .io_outs_down({\ces_1_1_io_ins_down[63] ,
    \ces_1_1_io_ins_down[62] ,
    \ces_1_1_io_ins_down[61] ,
    \ces_1_1_io_ins_down[60] ,
    \ces_1_1_io_ins_down[59] ,
    \ces_1_1_io_ins_down[58] ,
    \ces_1_1_io_ins_down[57] ,
    \ces_1_1_io_ins_down[56] ,
    \ces_1_1_io_ins_down[55] ,
    \ces_1_1_io_ins_down[54] ,
    \ces_1_1_io_ins_down[53] ,
    \ces_1_1_io_ins_down[52] ,
    \ces_1_1_io_ins_down[51] ,
    \ces_1_1_io_ins_down[50] ,
    \ces_1_1_io_ins_down[49] ,
    \ces_1_1_io_ins_down[48] ,
    \ces_1_1_io_ins_down[47] ,
    \ces_1_1_io_ins_down[46] ,
    \ces_1_1_io_ins_down[45] ,
    \ces_1_1_io_ins_down[44] ,
    \ces_1_1_io_ins_down[43] ,
    \ces_1_1_io_ins_down[42] ,
    \ces_1_1_io_ins_down[41] ,
    \ces_1_1_io_ins_down[40] ,
    \ces_1_1_io_ins_down[39] ,
    \ces_1_1_io_ins_down[38] ,
    \ces_1_1_io_ins_down[37] ,
    \ces_1_1_io_ins_down[36] ,
    \ces_1_1_io_ins_down[35] ,
    \ces_1_1_io_ins_down[34] ,
    \ces_1_1_io_ins_down[33] ,
    \ces_1_1_io_ins_down[32] ,
    \ces_1_1_io_ins_down[31] ,
    \ces_1_1_io_ins_down[30] ,
    \ces_1_1_io_ins_down[29] ,
    \ces_1_1_io_ins_down[28] ,
    \ces_1_1_io_ins_down[27] ,
    \ces_1_1_io_ins_down[26] ,
    \ces_1_1_io_ins_down[25] ,
    \ces_1_1_io_ins_down[24] ,
    \ces_1_1_io_ins_down[23] ,
    \ces_1_1_io_ins_down[22] ,
    \ces_1_1_io_ins_down[21] ,
    \ces_1_1_io_ins_down[20] ,
    \ces_1_1_io_ins_down[19] ,
    \ces_1_1_io_ins_down[18] ,
    \ces_1_1_io_ins_down[17] ,
    \ces_1_1_io_ins_down[16] ,
    \ces_1_1_io_ins_down[15] ,
    \ces_1_1_io_ins_down[14] ,
    \ces_1_1_io_ins_down[13] ,
    \ces_1_1_io_ins_down[12] ,
    \ces_1_1_io_ins_down[11] ,
    \ces_1_1_io_ins_down[10] ,
    \ces_1_1_io_ins_down[9] ,
    \ces_1_1_io_ins_down[8] ,
    \ces_1_1_io_ins_down[7] ,
    \ces_1_1_io_ins_down[6] ,
    \ces_1_1_io_ins_down[5] ,
    \ces_1_1_io_ins_down[4] ,
    \ces_1_1_io_ins_down[3] ,
    \ces_1_1_io_ins_down[2] ,
    \ces_1_1_io_ins_down[1] ,
    \ces_1_1_io_ins_down[0] }),
    .io_outs_left({\ces_2_0_io_ins_left[63] ,
    \ces_2_0_io_ins_left[62] ,
    \ces_2_0_io_ins_left[61] ,
    \ces_2_0_io_ins_left[60] ,
    \ces_2_0_io_ins_left[59] ,
    \ces_2_0_io_ins_left[58] ,
    \ces_2_0_io_ins_left[57] ,
    \ces_2_0_io_ins_left[56] ,
    \ces_2_0_io_ins_left[55] ,
    \ces_2_0_io_ins_left[54] ,
    \ces_2_0_io_ins_left[53] ,
    \ces_2_0_io_ins_left[52] ,
    \ces_2_0_io_ins_left[51] ,
    \ces_2_0_io_ins_left[50] ,
    \ces_2_0_io_ins_left[49] ,
    \ces_2_0_io_ins_left[48] ,
    \ces_2_0_io_ins_left[47] ,
    \ces_2_0_io_ins_left[46] ,
    \ces_2_0_io_ins_left[45] ,
    \ces_2_0_io_ins_left[44] ,
    \ces_2_0_io_ins_left[43] ,
    \ces_2_0_io_ins_left[42] ,
    \ces_2_0_io_ins_left[41] ,
    \ces_2_0_io_ins_left[40] ,
    \ces_2_0_io_ins_left[39] ,
    \ces_2_0_io_ins_left[38] ,
    \ces_2_0_io_ins_left[37] ,
    \ces_2_0_io_ins_left[36] ,
    \ces_2_0_io_ins_left[35] ,
    \ces_2_0_io_ins_left[34] ,
    \ces_2_0_io_ins_left[33] ,
    \ces_2_0_io_ins_left[32] ,
    \ces_2_0_io_ins_left[31] ,
    \ces_2_0_io_ins_left[30] ,
    \ces_2_0_io_ins_left[29] ,
    \ces_2_0_io_ins_left[28] ,
    \ces_2_0_io_ins_left[27] ,
    \ces_2_0_io_ins_left[26] ,
    \ces_2_0_io_ins_left[25] ,
    \ces_2_0_io_ins_left[24] ,
    \ces_2_0_io_ins_left[23] ,
    \ces_2_0_io_ins_left[22] ,
    \ces_2_0_io_ins_left[21] ,
    \ces_2_0_io_ins_left[20] ,
    \ces_2_0_io_ins_left[19] ,
    \ces_2_0_io_ins_left[18] ,
    \ces_2_0_io_ins_left[17] ,
    \ces_2_0_io_ins_left[16] ,
    \ces_2_0_io_ins_left[15] ,
    \ces_2_0_io_ins_left[14] ,
    \ces_2_0_io_ins_left[13] ,
    \ces_2_0_io_ins_left[12] ,
    \ces_2_0_io_ins_left[11] ,
    \ces_2_0_io_ins_left[10] ,
    \ces_2_0_io_ins_left[9] ,
    \ces_2_0_io_ins_left[8] ,
    \ces_2_0_io_ins_left[7] ,
    \ces_2_0_io_ins_left[6] ,
    \ces_2_0_io_ins_left[5] ,
    \ces_2_0_io_ins_left[4] ,
    \ces_2_0_io_ins_left[3] ,
    \ces_2_0_io_ins_left[2] ,
    \ces_2_0_io_ins_left[1] ,
    \ces_2_0_io_ins_left[0] }),
    .io_outs_right({\ces_2_1_io_outs_right[63] ,
    \ces_2_1_io_outs_right[62] ,
    \ces_2_1_io_outs_right[61] ,
    \ces_2_1_io_outs_right[60] ,
    \ces_2_1_io_outs_right[59] ,
    \ces_2_1_io_outs_right[58] ,
    \ces_2_1_io_outs_right[57] ,
    \ces_2_1_io_outs_right[56] ,
    \ces_2_1_io_outs_right[55] ,
    \ces_2_1_io_outs_right[54] ,
    \ces_2_1_io_outs_right[53] ,
    \ces_2_1_io_outs_right[52] ,
    \ces_2_1_io_outs_right[51] ,
    \ces_2_1_io_outs_right[50] ,
    \ces_2_1_io_outs_right[49] ,
    \ces_2_1_io_outs_right[48] ,
    \ces_2_1_io_outs_right[47] ,
    \ces_2_1_io_outs_right[46] ,
    \ces_2_1_io_outs_right[45] ,
    \ces_2_1_io_outs_right[44] ,
    \ces_2_1_io_outs_right[43] ,
    \ces_2_1_io_outs_right[42] ,
    \ces_2_1_io_outs_right[41] ,
    \ces_2_1_io_outs_right[40] ,
    \ces_2_1_io_outs_right[39] ,
    \ces_2_1_io_outs_right[38] ,
    \ces_2_1_io_outs_right[37] ,
    \ces_2_1_io_outs_right[36] ,
    \ces_2_1_io_outs_right[35] ,
    \ces_2_1_io_outs_right[34] ,
    \ces_2_1_io_outs_right[33] ,
    \ces_2_1_io_outs_right[32] ,
    \ces_2_1_io_outs_right[31] ,
    \ces_2_1_io_outs_right[30] ,
    \ces_2_1_io_outs_right[29] ,
    \ces_2_1_io_outs_right[28] ,
    \ces_2_1_io_outs_right[27] ,
    \ces_2_1_io_outs_right[26] ,
    \ces_2_1_io_outs_right[25] ,
    \ces_2_1_io_outs_right[24] ,
    \ces_2_1_io_outs_right[23] ,
    \ces_2_1_io_outs_right[22] ,
    \ces_2_1_io_outs_right[21] ,
    \ces_2_1_io_outs_right[20] ,
    \ces_2_1_io_outs_right[19] ,
    \ces_2_1_io_outs_right[18] ,
    \ces_2_1_io_outs_right[17] ,
    \ces_2_1_io_outs_right[16] ,
    \ces_2_1_io_outs_right[15] ,
    \ces_2_1_io_outs_right[14] ,
    \ces_2_1_io_outs_right[13] ,
    \ces_2_1_io_outs_right[12] ,
    \ces_2_1_io_outs_right[11] ,
    \ces_2_1_io_outs_right[10] ,
    \ces_2_1_io_outs_right[9] ,
    \ces_2_1_io_outs_right[8] ,
    \ces_2_1_io_outs_right[7] ,
    \ces_2_1_io_outs_right[6] ,
    \ces_2_1_io_outs_right[5] ,
    \ces_2_1_io_outs_right[4] ,
    \ces_2_1_io_outs_right[3] ,
    \ces_2_1_io_outs_right[2] ,
    \ces_2_1_io_outs_right[1] ,
    \ces_2_1_io_outs_right[0] }),
    .io_outs_up({\ces_2_1_io_outs_up[63] ,
    \ces_2_1_io_outs_up[62] ,
    \ces_2_1_io_outs_up[61] ,
    \ces_2_1_io_outs_up[60] ,
    \ces_2_1_io_outs_up[59] ,
    \ces_2_1_io_outs_up[58] ,
    \ces_2_1_io_outs_up[57] ,
    \ces_2_1_io_outs_up[56] ,
    \ces_2_1_io_outs_up[55] ,
    \ces_2_1_io_outs_up[54] ,
    \ces_2_1_io_outs_up[53] ,
    \ces_2_1_io_outs_up[52] ,
    \ces_2_1_io_outs_up[51] ,
    \ces_2_1_io_outs_up[50] ,
    \ces_2_1_io_outs_up[49] ,
    \ces_2_1_io_outs_up[48] ,
    \ces_2_1_io_outs_up[47] ,
    \ces_2_1_io_outs_up[46] ,
    \ces_2_1_io_outs_up[45] ,
    \ces_2_1_io_outs_up[44] ,
    \ces_2_1_io_outs_up[43] ,
    \ces_2_1_io_outs_up[42] ,
    \ces_2_1_io_outs_up[41] ,
    \ces_2_1_io_outs_up[40] ,
    \ces_2_1_io_outs_up[39] ,
    \ces_2_1_io_outs_up[38] ,
    \ces_2_1_io_outs_up[37] ,
    \ces_2_1_io_outs_up[36] ,
    \ces_2_1_io_outs_up[35] ,
    \ces_2_1_io_outs_up[34] ,
    \ces_2_1_io_outs_up[33] ,
    \ces_2_1_io_outs_up[32] ,
    \ces_2_1_io_outs_up[31] ,
    \ces_2_1_io_outs_up[30] ,
    \ces_2_1_io_outs_up[29] ,
    \ces_2_1_io_outs_up[28] ,
    \ces_2_1_io_outs_up[27] ,
    \ces_2_1_io_outs_up[26] ,
    \ces_2_1_io_outs_up[25] ,
    \ces_2_1_io_outs_up[24] ,
    \ces_2_1_io_outs_up[23] ,
    \ces_2_1_io_outs_up[22] ,
    \ces_2_1_io_outs_up[21] ,
    \ces_2_1_io_outs_up[20] ,
    \ces_2_1_io_outs_up[19] ,
    \ces_2_1_io_outs_up[18] ,
    \ces_2_1_io_outs_up[17] ,
    \ces_2_1_io_outs_up[16] ,
    \ces_2_1_io_outs_up[15] ,
    \ces_2_1_io_outs_up[14] ,
    \ces_2_1_io_outs_up[13] ,
    \ces_2_1_io_outs_up[12] ,
    \ces_2_1_io_outs_up[11] ,
    \ces_2_1_io_outs_up[10] ,
    \ces_2_1_io_outs_up[9] ,
    \ces_2_1_io_outs_up[8] ,
    \ces_2_1_io_outs_up[7] ,
    \ces_2_1_io_outs_up[6] ,
    \ces_2_1_io_outs_up[5] ,
    \ces_2_1_io_outs_up[4] ,
    \ces_2_1_io_outs_up[3] ,
    \ces_2_1_io_outs_up[2] ,
    \ces_2_1_io_outs_up[1] ,
    \ces_2_1_io_outs_up[0] }));
 Element ces_2_2 (.clock(clknet_3_1_0_clock),
    .io_lsbIns_1(ces_2_1_io_lsbOuts_1),
    .io_lsbIns_2(ces_2_1_io_lsbOuts_2),
    .io_lsbIns_3(ces_2_1_io_lsbOuts_3),
    .io_lsbIns_4(ces_2_1_io_lsbOuts_4),
    .io_lsbIns_5(ces_2_1_io_lsbOuts_5),
    .io_lsbIns_6(ces_2_1_io_lsbOuts_6),
    .io_lsbIns_7(ces_2_1_io_lsbOuts_7),
    .io_lsbOuts_0(ces_2_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_2_io_lsbOuts_7),
    .io_ins_down({\ces_2_2_io_ins_down[63] ,
    \ces_2_2_io_ins_down[62] ,
    \ces_2_2_io_ins_down[61] ,
    \ces_2_2_io_ins_down[60] ,
    \ces_2_2_io_ins_down[59] ,
    \ces_2_2_io_ins_down[58] ,
    \ces_2_2_io_ins_down[57] ,
    \ces_2_2_io_ins_down[56] ,
    \ces_2_2_io_ins_down[55] ,
    \ces_2_2_io_ins_down[54] ,
    \ces_2_2_io_ins_down[53] ,
    \ces_2_2_io_ins_down[52] ,
    \ces_2_2_io_ins_down[51] ,
    \ces_2_2_io_ins_down[50] ,
    \ces_2_2_io_ins_down[49] ,
    \ces_2_2_io_ins_down[48] ,
    \ces_2_2_io_ins_down[47] ,
    \ces_2_2_io_ins_down[46] ,
    \ces_2_2_io_ins_down[45] ,
    \ces_2_2_io_ins_down[44] ,
    \ces_2_2_io_ins_down[43] ,
    \ces_2_2_io_ins_down[42] ,
    \ces_2_2_io_ins_down[41] ,
    \ces_2_2_io_ins_down[40] ,
    \ces_2_2_io_ins_down[39] ,
    \ces_2_2_io_ins_down[38] ,
    \ces_2_2_io_ins_down[37] ,
    \ces_2_2_io_ins_down[36] ,
    \ces_2_2_io_ins_down[35] ,
    \ces_2_2_io_ins_down[34] ,
    \ces_2_2_io_ins_down[33] ,
    \ces_2_2_io_ins_down[32] ,
    \ces_2_2_io_ins_down[31] ,
    \ces_2_2_io_ins_down[30] ,
    \ces_2_2_io_ins_down[29] ,
    \ces_2_2_io_ins_down[28] ,
    \ces_2_2_io_ins_down[27] ,
    \ces_2_2_io_ins_down[26] ,
    \ces_2_2_io_ins_down[25] ,
    \ces_2_2_io_ins_down[24] ,
    \ces_2_2_io_ins_down[23] ,
    \ces_2_2_io_ins_down[22] ,
    \ces_2_2_io_ins_down[21] ,
    \ces_2_2_io_ins_down[20] ,
    \ces_2_2_io_ins_down[19] ,
    \ces_2_2_io_ins_down[18] ,
    \ces_2_2_io_ins_down[17] ,
    \ces_2_2_io_ins_down[16] ,
    \ces_2_2_io_ins_down[15] ,
    \ces_2_2_io_ins_down[14] ,
    \ces_2_2_io_ins_down[13] ,
    \ces_2_2_io_ins_down[12] ,
    \ces_2_2_io_ins_down[11] ,
    \ces_2_2_io_ins_down[10] ,
    \ces_2_2_io_ins_down[9] ,
    \ces_2_2_io_ins_down[8] ,
    \ces_2_2_io_ins_down[7] ,
    \ces_2_2_io_ins_down[6] ,
    \ces_2_2_io_ins_down[5] ,
    \ces_2_2_io_ins_down[4] ,
    \ces_2_2_io_ins_down[3] ,
    \ces_2_2_io_ins_down[2] ,
    \ces_2_2_io_ins_down[1] ,
    \ces_2_2_io_ins_down[0] }),
    .io_ins_left({\ces_2_2_io_ins_left[63] ,
    \ces_2_2_io_ins_left[62] ,
    \ces_2_2_io_ins_left[61] ,
    \ces_2_2_io_ins_left[60] ,
    \ces_2_2_io_ins_left[59] ,
    \ces_2_2_io_ins_left[58] ,
    \ces_2_2_io_ins_left[57] ,
    \ces_2_2_io_ins_left[56] ,
    \ces_2_2_io_ins_left[55] ,
    \ces_2_2_io_ins_left[54] ,
    \ces_2_2_io_ins_left[53] ,
    \ces_2_2_io_ins_left[52] ,
    \ces_2_2_io_ins_left[51] ,
    \ces_2_2_io_ins_left[50] ,
    \ces_2_2_io_ins_left[49] ,
    \ces_2_2_io_ins_left[48] ,
    \ces_2_2_io_ins_left[47] ,
    \ces_2_2_io_ins_left[46] ,
    \ces_2_2_io_ins_left[45] ,
    \ces_2_2_io_ins_left[44] ,
    \ces_2_2_io_ins_left[43] ,
    \ces_2_2_io_ins_left[42] ,
    \ces_2_2_io_ins_left[41] ,
    \ces_2_2_io_ins_left[40] ,
    \ces_2_2_io_ins_left[39] ,
    \ces_2_2_io_ins_left[38] ,
    \ces_2_2_io_ins_left[37] ,
    \ces_2_2_io_ins_left[36] ,
    \ces_2_2_io_ins_left[35] ,
    \ces_2_2_io_ins_left[34] ,
    \ces_2_2_io_ins_left[33] ,
    \ces_2_2_io_ins_left[32] ,
    \ces_2_2_io_ins_left[31] ,
    \ces_2_2_io_ins_left[30] ,
    \ces_2_2_io_ins_left[29] ,
    \ces_2_2_io_ins_left[28] ,
    \ces_2_2_io_ins_left[27] ,
    \ces_2_2_io_ins_left[26] ,
    \ces_2_2_io_ins_left[25] ,
    \ces_2_2_io_ins_left[24] ,
    \ces_2_2_io_ins_left[23] ,
    \ces_2_2_io_ins_left[22] ,
    \ces_2_2_io_ins_left[21] ,
    \ces_2_2_io_ins_left[20] ,
    \ces_2_2_io_ins_left[19] ,
    \ces_2_2_io_ins_left[18] ,
    \ces_2_2_io_ins_left[17] ,
    \ces_2_2_io_ins_left[16] ,
    \ces_2_2_io_ins_left[15] ,
    \ces_2_2_io_ins_left[14] ,
    \ces_2_2_io_ins_left[13] ,
    \ces_2_2_io_ins_left[12] ,
    \ces_2_2_io_ins_left[11] ,
    \ces_2_2_io_ins_left[10] ,
    \ces_2_2_io_ins_left[9] ,
    \ces_2_2_io_ins_left[8] ,
    \ces_2_2_io_ins_left[7] ,
    \ces_2_2_io_ins_left[6] ,
    \ces_2_2_io_ins_left[5] ,
    \ces_2_2_io_ins_left[4] ,
    \ces_2_2_io_ins_left[3] ,
    \ces_2_2_io_ins_left[2] ,
    \ces_2_2_io_ins_left[1] ,
    \ces_2_2_io_ins_left[0] }),
    .io_ins_right({\ces_2_1_io_outs_right[63] ,
    \ces_2_1_io_outs_right[62] ,
    \ces_2_1_io_outs_right[61] ,
    \ces_2_1_io_outs_right[60] ,
    \ces_2_1_io_outs_right[59] ,
    \ces_2_1_io_outs_right[58] ,
    \ces_2_1_io_outs_right[57] ,
    \ces_2_1_io_outs_right[56] ,
    \ces_2_1_io_outs_right[55] ,
    \ces_2_1_io_outs_right[54] ,
    \ces_2_1_io_outs_right[53] ,
    \ces_2_1_io_outs_right[52] ,
    \ces_2_1_io_outs_right[51] ,
    \ces_2_1_io_outs_right[50] ,
    \ces_2_1_io_outs_right[49] ,
    \ces_2_1_io_outs_right[48] ,
    \ces_2_1_io_outs_right[47] ,
    \ces_2_1_io_outs_right[46] ,
    \ces_2_1_io_outs_right[45] ,
    \ces_2_1_io_outs_right[44] ,
    \ces_2_1_io_outs_right[43] ,
    \ces_2_1_io_outs_right[42] ,
    \ces_2_1_io_outs_right[41] ,
    \ces_2_1_io_outs_right[40] ,
    \ces_2_1_io_outs_right[39] ,
    \ces_2_1_io_outs_right[38] ,
    \ces_2_1_io_outs_right[37] ,
    \ces_2_1_io_outs_right[36] ,
    \ces_2_1_io_outs_right[35] ,
    \ces_2_1_io_outs_right[34] ,
    \ces_2_1_io_outs_right[33] ,
    \ces_2_1_io_outs_right[32] ,
    \ces_2_1_io_outs_right[31] ,
    \ces_2_1_io_outs_right[30] ,
    \ces_2_1_io_outs_right[29] ,
    \ces_2_1_io_outs_right[28] ,
    \ces_2_1_io_outs_right[27] ,
    \ces_2_1_io_outs_right[26] ,
    \ces_2_1_io_outs_right[25] ,
    \ces_2_1_io_outs_right[24] ,
    \ces_2_1_io_outs_right[23] ,
    \ces_2_1_io_outs_right[22] ,
    \ces_2_1_io_outs_right[21] ,
    \ces_2_1_io_outs_right[20] ,
    \ces_2_1_io_outs_right[19] ,
    \ces_2_1_io_outs_right[18] ,
    \ces_2_1_io_outs_right[17] ,
    \ces_2_1_io_outs_right[16] ,
    \ces_2_1_io_outs_right[15] ,
    \ces_2_1_io_outs_right[14] ,
    \ces_2_1_io_outs_right[13] ,
    \ces_2_1_io_outs_right[12] ,
    \ces_2_1_io_outs_right[11] ,
    \ces_2_1_io_outs_right[10] ,
    \ces_2_1_io_outs_right[9] ,
    \ces_2_1_io_outs_right[8] ,
    \ces_2_1_io_outs_right[7] ,
    \ces_2_1_io_outs_right[6] ,
    \ces_2_1_io_outs_right[5] ,
    \ces_2_1_io_outs_right[4] ,
    \ces_2_1_io_outs_right[3] ,
    \ces_2_1_io_outs_right[2] ,
    \ces_2_1_io_outs_right[1] ,
    \ces_2_1_io_outs_right[0] }),
    .io_ins_up({\ces_1_2_io_outs_up[63] ,
    \ces_1_2_io_outs_up[62] ,
    \ces_1_2_io_outs_up[61] ,
    \ces_1_2_io_outs_up[60] ,
    \ces_1_2_io_outs_up[59] ,
    \ces_1_2_io_outs_up[58] ,
    \ces_1_2_io_outs_up[57] ,
    \ces_1_2_io_outs_up[56] ,
    \ces_1_2_io_outs_up[55] ,
    \ces_1_2_io_outs_up[54] ,
    \ces_1_2_io_outs_up[53] ,
    \ces_1_2_io_outs_up[52] ,
    \ces_1_2_io_outs_up[51] ,
    \ces_1_2_io_outs_up[50] ,
    \ces_1_2_io_outs_up[49] ,
    \ces_1_2_io_outs_up[48] ,
    \ces_1_2_io_outs_up[47] ,
    \ces_1_2_io_outs_up[46] ,
    \ces_1_2_io_outs_up[45] ,
    \ces_1_2_io_outs_up[44] ,
    \ces_1_2_io_outs_up[43] ,
    \ces_1_2_io_outs_up[42] ,
    \ces_1_2_io_outs_up[41] ,
    \ces_1_2_io_outs_up[40] ,
    \ces_1_2_io_outs_up[39] ,
    \ces_1_2_io_outs_up[38] ,
    \ces_1_2_io_outs_up[37] ,
    \ces_1_2_io_outs_up[36] ,
    \ces_1_2_io_outs_up[35] ,
    \ces_1_2_io_outs_up[34] ,
    \ces_1_2_io_outs_up[33] ,
    \ces_1_2_io_outs_up[32] ,
    \ces_1_2_io_outs_up[31] ,
    \ces_1_2_io_outs_up[30] ,
    \ces_1_2_io_outs_up[29] ,
    \ces_1_2_io_outs_up[28] ,
    \ces_1_2_io_outs_up[27] ,
    \ces_1_2_io_outs_up[26] ,
    \ces_1_2_io_outs_up[25] ,
    \ces_1_2_io_outs_up[24] ,
    \ces_1_2_io_outs_up[23] ,
    \ces_1_2_io_outs_up[22] ,
    \ces_1_2_io_outs_up[21] ,
    \ces_1_2_io_outs_up[20] ,
    \ces_1_2_io_outs_up[19] ,
    \ces_1_2_io_outs_up[18] ,
    \ces_1_2_io_outs_up[17] ,
    \ces_1_2_io_outs_up[16] ,
    \ces_1_2_io_outs_up[15] ,
    \ces_1_2_io_outs_up[14] ,
    \ces_1_2_io_outs_up[13] ,
    \ces_1_2_io_outs_up[12] ,
    \ces_1_2_io_outs_up[11] ,
    \ces_1_2_io_outs_up[10] ,
    \ces_1_2_io_outs_up[9] ,
    \ces_1_2_io_outs_up[8] ,
    \ces_1_2_io_outs_up[7] ,
    \ces_1_2_io_outs_up[6] ,
    \ces_1_2_io_outs_up[5] ,
    \ces_1_2_io_outs_up[4] ,
    \ces_1_2_io_outs_up[3] ,
    \ces_1_2_io_outs_up[2] ,
    \ces_1_2_io_outs_up[1] ,
    \ces_1_2_io_outs_up[0] }),
    .io_outs_down({\ces_1_2_io_ins_down[63] ,
    \ces_1_2_io_ins_down[62] ,
    \ces_1_2_io_ins_down[61] ,
    \ces_1_2_io_ins_down[60] ,
    \ces_1_2_io_ins_down[59] ,
    \ces_1_2_io_ins_down[58] ,
    \ces_1_2_io_ins_down[57] ,
    \ces_1_2_io_ins_down[56] ,
    \ces_1_2_io_ins_down[55] ,
    \ces_1_2_io_ins_down[54] ,
    \ces_1_2_io_ins_down[53] ,
    \ces_1_2_io_ins_down[52] ,
    \ces_1_2_io_ins_down[51] ,
    \ces_1_2_io_ins_down[50] ,
    \ces_1_2_io_ins_down[49] ,
    \ces_1_2_io_ins_down[48] ,
    \ces_1_2_io_ins_down[47] ,
    \ces_1_2_io_ins_down[46] ,
    \ces_1_2_io_ins_down[45] ,
    \ces_1_2_io_ins_down[44] ,
    \ces_1_2_io_ins_down[43] ,
    \ces_1_2_io_ins_down[42] ,
    \ces_1_2_io_ins_down[41] ,
    \ces_1_2_io_ins_down[40] ,
    \ces_1_2_io_ins_down[39] ,
    \ces_1_2_io_ins_down[38] ,
    \ces_1_2_io_ins_down[37] ,
    \ces_1_2_io_ins_down[36] ,
    \ces_1_2_io_ins_down[35] ,
    \ces_1_2_io_ins_down[34] ,
    \ces_1_2_io_ins_down[33] ,
    \ces_1_2_io_ins_down[32] ,
    \ces_1_2_io_ins_down[31] ,
    \ces_1_2_io_ins_down[30] ,
    \ces_1_2_io_ins_down[29] ,
    \ces_1_2_io_ins_down[28] ,
    \ces_1_2_io_ins_down[27] ,
    \ces_1_2_io_ins_down[26] ,
    \ces_1_2_io_ins_down[25] ,
    \ces_1_2_io_ins_down[24] ,
    \ces_1_2_io_ins_down[23] ,
    \ces_1_2_io_ins_down[22] ,
    \ces_1_2_io_ins_down[21] ,
    \ces_1_2_io_ins_down[20] ,
    \ces_1_2_io_ins_down[19] ,
    \ces_1_2_io_ins_down[18] ,
    \ces_1_2_io_ins_down[17] ,
    \ces_1_2_io_ins_down[16] ,
    \ces_1_2_io_ins_down[15] ,
    \ces_1_2_io_ins_down[14] ,
    \ces_1_2_io_ins_down[13] ,
    \ces_1_2_io_ins_down[12] ,
    \ces_1_2_io_ins_down[11] ,
    \ces_1_2_io_ins_down[10] ,
    \ces_1_2_io_ins_down[9] ,
    \ces_1_2_io_ins_down[8] ,
    \ces_1_2_io_ins_down[7] ,
    \ces_1_2_io_ins_down[6] ,
    \ces_1_2_io_ins_down[5] ,
    \ces_1_2_io_ins_down[4] ,
    \ces_1_2_io_ins_down[3] ,
    \ces_1_2_io_ins_down[2] ,
    \ces_1_2_io_ins_down[1] ,
    \ces_1_2_io_ins_down[0] }),
    .io_outs_left({\ces_2_1_io_ins_left[63] ,
    \ces_2_1_io_ins_left[62] ,
    \ces_2_1_io_ins_left[61] ,
    \ces_2_1_io_ins_left[60] ,
    \ces_2_1_io_ins_left[59] ,
    \ces_2_1_io_ins_left[58] ,
    \ces_2_1_io_ins_left[57] ,
    \ces_2_1_io_ins_left[56] ,
    \ces_2_1_io_ins_left[55] ,
    \ces_2_1_io_ins_left[54] ,
    \ces_2_1_io_ins_left[53] ,
    \ces_2_1_io_ins_left[52] ,
    \ces_2_1_io_ins_left[51] ,
    \ces_2_1_io_ins_left[50] ,
    \ces_2_1_io_ins_left[49] ,
    \ces_2_1_io_ins_left[48] ,
    \ces_2_1_io_ins_left[47] ,
    \ces_2_1_io_ins_left[46] ,
    \ces_2_1_io_ins_left[45] ,
    \ces_2_1_io_ins_left[44] ,
    \ces_2_1_io_ins_left[43] ,
    \ces_2_1_io_ins_left[42] ,
    \ces_2_1_io_ins_left[41] ,
    \ces_2_1_io_ins_left[40] ,
    \ces_2_1_io_ins_left[39] ,
    \ces_2_1_io_ins_left[38] ,
    \ces_2_1_io_ins_left[37] ,
    \ces_2_1_io_ins_left[36] ,
    \ces_2_1_io_ins_left[35] ,
    \ces_2_1_io_ins_left[34] ,
    \ces_2_1_io_ins_left[33] ,
    \ces_2_1_io_ins_left[32] ,
    \ces_2_1_io_ins_left[31] ,
    \ces_2_1_io_ins_left[30] ,
    \ces_2_1_io_ins_left[29] ,
    \ces_2_1_io_ins_left[28] ,
    \ces_2_1_io_ins_left[27] ,
    \ces_2_1_io_ins_left[26] ,
    \ces_2_1_io_ins_left[25] ,
    \ces_2_1_io_ins_left[24] ,
    \ces_2_1_io_ins_left[23] ,
    \ces_2_1_io_ins_left[22] ,
    \ces_2_1_io_ins_left[21] ,
    \ces_2_1_io_ins_left[20] ,
    \ces_2_1_io_ins_left[19] ,
    \ces_2_1_io_ins_left[18] ,
    \ces_2_1_io_ins_left[17] ,
    \ces_2_1_io_ins_left[16] ,
    \ces_2_1_io_ins_left[15] ,
    \ces_2_1_io_ins_left[14] ,
    \ces_2_1_io_ins_left[13] ,
    \ces_2_1_io_ins_left[12] ,
    \ces_2_1_io_ins_left[11] ,
    \ces_2_1_io_ins_left[10] ,
    \ces_2_1_io_ins_left[9] ,
    \ces_2_1_io_ins_left[8] ,
    \ces_2_1_io_ins_left[7] ,
    \ces_2_1_io_ins_left[6] ,
    \ces_2_1_io_ins_left[5] ,
    \ces_2_1_io_ins_left[4] ,
    \ces_2_1_io_ins_left[3] ,
    \ces_2_1_io_ins_left[2] ,
    \ces_2_1_io_ins_left[1] ,
    \ces_2_1_io_ins_left[0] }),
    .io_outs_right({\ces_2_2_io_outs_right[63] ,
    \ces_2_2_io_outs_right[62] ,
    \ces_2_2_io_outs_right[61] ,
    \ces_2_2_io_outs_right[60] ,
    \ces_2_2_io_outs_right[59] ,
    \ces_2_2_io_outs_right[58] ,
    \ces_2_2_io_outs_right[57] ,
    \ces_2_2_io_outs_right[56] ,
    \ces_2_2_io_outs_right[55] ,
    \ces_2_2_io_outs_right[54] ,
    \ces_2_2_io_outs_right[53] ,
    \ces_2_2_io_outs_right[52] ,
    \ces_2_2_io_outs_right[51] ,
    \ces_2_2_io_outs_right[50] ,
    \ces_2_2_io_outs_right[49] ,
    \ces_2_2_io_outs_right[48] ,
    \ces_2_2_io_outs_right[47] ,
    \ces_2_2_io_outs_right[46] ,
    \ces_2_2_io_outs_right[45] ,
    \ces_2_2_io_outs_right[44] ,
    \ces_2_2_io_outs_right[43] ,
    \ces_2_2_io_outs_right[42] ,
    \ces_2_2_io_outs_right[41] ,
    \ces_2_2_io_outs_right[40] ,
    \ces_2_2_io_outs_right[39] ,
    \ces_2_2_io_outs_right[38] ,
    \ces_2_2_io_outs_right[37] ,
    \ces_2_2_io_outs_right[36] ,
    \ces_2_2_io_outs_right[35] ,
    \ces_2_2_io_outs_right[34] ,
    \ces_2_2_io_outs_right[33] ,
    \ces_2_2_io_outs_right[32] ,
    \ces_2_2_io_outs_right[31] ,
    \ces_2_2_io_outs_right[30] ,
    \ces_2_2_io_outs_right[29] ,
    \ces_2_2_io_outs_right[28] ,
    \ces_2_2_io_outs_right[27] ,
    \ces_2_2_io_outs_right[26] ,
    \ces_2_2_io_outs_right[25] ,
    \ces_2_2_io_outs_right[24] ,
    \ces_2_2_io_outs_right[23] ,
    \ces_2_2_io_outs_right[22] ,
    \ces_2_2_io_outs_right[21] ,
    \ces_2_2_io_outs_right[20] ,
    \ces_2_2_io_outs_right[19] ,
    \ces_2_2_io_outs_right[18] ,
    \ces_2_2_io_outs_right[17] ,
    \ces_2_2_io_outs_right[16] ,
    \ces_2_2_io_outs_right[15] ,
    \ces_2_2_io_outs_right[14] ,
    \ces_2_2_io_outs_right[13] ,
    \ces_2_2_io_outs_right[12] ,
    \ces_2_2_io_outs_right[11] ,
    \ces_2_2_io_outs_right[10] ,
    \ces_2_2_io_outs_right[9] ,
    \ces_2_2_io_outs_right[8] ,
    \ces_2_2_io_outs_right[7] ,
    \ces_2_2_io_outs_right[6] ,
    \ces_2_2_io_outs_right[5] ,
    \ces_2_2_io_outs_right[4] ,
    \ces_2_2_io_outs_right[3] ,
    \ces_2_2_io_outs_right[2] ,
    \ces_2_2_io_outs_right[1] ,
    \ces_2_2_io_outs_right[0] }),
    .io_outs_up({\ces_2_2_io_outs_up[63] ,
    \ces_2_2_io_outs_up[62] ,
    \ces_2_2_io_outs_up[61] ,
    \ces_2_2_io_outs_up[60] ,
    \ces_2_2_io_outs_up[59] ,
    \ces_2_2_io_outs_up[58] ,
    \ces_2_2_io_outs_up[57] ,
    \ces_2_2_io_outs_up[56] ,
    \ces_2_2_io_outs_up[55] ,
    \ces_2_2_io_outs_up[54] ,
    \ces_2_2_io_outs_up[53] ,
    \ces_2_2_io_outs_up[52] ,
    \ces_2_2_io_outs_up[51] ,
    \ces_2_2_io_outs_up[50] ,
    \ces_2_2_io_outs_up[49] ,
    \ces_2_2_io_outs_up[48] ,
    \ces_2_2_io_outs_up[47] ,
    \ces_2_2_io_outs_up[46] ,
    \ces_2_2_io_outs_up[45] ,
    \ces_2_2_io_outs_up[44] ,
    \ces_2_2_io_outs_up[43] ,
    \ces_2_2_io_outs_up[42] ,
    \ces_2_2_io_outs_up[41] ,
    \ces_2_2_io_outs_up[40] ,
    \ces_2_2_io_outs_up[39] ,
    \ces_2_2_io_outs_up[38] ,
    \ces_2_2_io_outs_up[37] ,
    \ces_2_2_io_outs_up[36] ,
    \ces_2_2_io_outs_up[35] ,
    \ces_2_2_io_outs_up[34] ,
    \ces_2_2_io_outs_up[33] ,
    \ces_2_2_io_outs_up[32] ,
    \ces_2_2_io_outs_up[31] ,
    \ces_2_2_io_outs_up[30] ,
    \ces_2_2_io_outs_up[29] ,
    \ces_2_2_io_outs_up[28] ,
    \ces_2_2_io_outs_up[27] ,
    \ces_2_2_io_outs_up[26] ,
    \ces_2_2_io_outs_up[25] ,
    \ces_2_2_io_outs_up[24] ,
    \ces_2_2_io_outs_up[23] ,
    \ces_2_2_io_outs_up[22] ,
    \ces_2_2_io_outs_up[21] ,
    \ces_2_2_io_outs_up[20] ,
    \ces_2_2_io_outs_up[19] ,
    \ces_2_2_io_outs_up[18] ,
    \ces_2_2_io_outs_up[17] ,
    \ces_2_2_io_outs_up[16] ,
    \ces_2_2_io_outs_up[15] ,
    \ces_2_2_io_outs_up[14] ,
    \ces_2_2_io_outs_up[13] ,
    \ces_2_2_io_outs_up[12] ,
    \ces_2_2_io_outs_up[11] ,
    \ces_2_2_io_outs_up[10] ,
    \ces_2_2_io_outs_up[9] ,
    \ces_2_2_io_outs_up[8] ,
    \ces_2_2_io_outs_up[7] ,
    \ces_2_2_io_outs_up[6] ,
    \ces_2_2_io_outs_up[5] ,
    \ces_2_2_io_outs_up[4] ,
    \ces_2_2_io_outs_up[3] ,
    \ces_2_2_io_outs_up[2] ,
    \ces_2_2_io_outs_up[1] ,
    \ces_2_2_io_outs_up[0] }));
 Element ces_2_3 (.clock(clknet_3_1_0_clock),
    .io_lsbIns_1(ces_2_2_io_lsbOuts_1),
    .io_lsbIns_2(ces_2_2_io_lsbOuts_2),
    .io_lsbIns_3(ces_2_2_io_lsbOuts_3),
    .io_lsbIns_4(ces_2_2_io_lsbOuts_4),
    .io_lsbIns_5(ces_2_2_io_lsbOuts_5),
    .io_lsbIns_6(ces_2_2_io_lsbOuts_6),
    .io_lsbIns_7(ces_2_2_io_lsbOuts_7),
    .io_lsbOuts_0(ces_2_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_3_io_lsbOuts_7),
    .io_ins_down({\ces_2_3_io_ins_down[63] ,
    \ces_2_3_io_ins_down[62] ,
    \ces_2_3_io_ins_down[61] ,
    \ces_2_3_io_ins_down[60] ,
    \ces_2_3_io_ins_down[59] ,
    \ces_2_3_io_ins_down[58] ,
    \ces_2_3_io_ins_down[57] ,
    \ces_2_3_io_ins_down[56] ,
    \ces_2_3_io_ins_down[55] ,
    \ces_2_3_io_ins_down[54] ,
    \ces_2_3_io_ins_down[53] ,
    \ces_2_3_io_ins_down[52] ,
    \ces_2_3_io_ins_down[51] ,
    \ces_2_3_io_ins_down[50] ,
    \ces_2_3_io_ins_down[49] ,
    \ces_2_3_io_ins_down[48] ,
    \ces_2_3_io_ins_down[47] ,
    \ces_2_3_io_ins_down[46] ,
    \ces_2_3_io_ins_down[45] ,
    \ces_2_3_io_ins_down[44] ,
    \ces_2_3_io_ins_down[43] ,
    \ces_2_3_io_ins_down[42] ,
    \ces_2_3_io_ins_down[41] ,
    \ces_2_3_io_ins_down[40] ,
    \ces_2_3_io_ins_down[39] ,
    \ces_2_3_io_ins_down[38] ,
    \ces_2_3_io_ins_down[37] ,
    \ces_2_3_io_ins_down[36] ,
    \ces_2_3_io_ins_down[35] ,
    \ces_2_3_io_ins_down[34] ,
    \ces_2_3_io_ins_down[33] ,
    \ces_2_3_io_ins_down[32] ,
    \ces_2_3_io_ins_down[31] ,
    \ces_2_3_io_ins_down[30] ,
    \ces_2_3_io_ins_down[29] ,
    \ces_2_3_io_ins_down[28] ,
    \ces_2_3_io_ins_down[27] ,
    \ces_2_3_io_ins_down[26] ,
    \ces_2_3_io_ins_down[25] ,
    \ces_2_3_io_ins_down[24] ,
    \ces_2_3_io_ins_down[23] ,
    \ces_2_3_io_ins_down[22] ,
    \ces_2_3_io_ins_down[21] ,
    \ces_2_3_io_ins_down[20] ,
    \ces_2_3_io_ins_down[19] ,
    \ces_2_3_io_ins_down[18] ,
    \ces_2_3_io_ins_down[17] ,
    \ces_2_3_io_ins_down[16] ,
    \ces_2_3_io_ins_down[15] ,
    \ces_2_3_io_ins_down[14] ,
    \ces_2_3_io_ins_down[13] ,
    \ces_2_3_io_ins_down[12] ,
    \ces_2_3_io_ins_down[11] ,
    \ces_2_3_io_ins_down[10] ,
    \ces_2_3_io_ins_down[9] ,
    \ces_2_3_io_ins_down[8] ,
    \ces_2_3_io_ins_down[7] ,
    \ces_2_3_io_ins_down[6] ,
    \ces_2_3_io_ins_down[5] ,
    \ces_2_3_io_ins_down[4] ,
    \ces_2_3_io_ins_down[3] ,
    \ces_2_3_io_ins_down[2] ,
    \ces_2_3_io_ins_down[1] ,
    \ces_2_3_io_ins_down[0] }),
    .io_ins_left({\ces_2_3_io_ins_left[63] ,
    \ces_2_3_io_ins_left[62] ,
    \ces_2_3_io_ins_left[61] ,
    \ces_2_3_io_ins_left[60] ,
    \ces_2_3_io_ins_left[59] ,
    \ces_2_3_io_ins_left[58] ,
    \ces_2_3_io_ins_left[57] ,
    \ces_2_3_io_ins_left[56] ,
    \ces_2_3_io_ins_left[55] ,
    \ces_2_3_io_ins_left[54] ,
    \ces_2_3_io_ins_left[53] ,
    \ces_2_3_io_ins_left[52] ,
    \ces_2_3_io_ins_left[51] ,
    \ces_2_3_io_ins_left[50] ,
    \ces_2_3_io_ins_left[49] ,
    \ces_2_3_io_ins_left[48] ,
    \ces_2_3_io_ins_left[47] ,
    \ces_2_3_io_ins_left[46] ,
    \ces_2_3_io_ins_left[45] ,
    \ces_2_3_io_ins_left[44] ,
    \ces_2_3_io_ins_left[43] ,
    \ces_2_3_io_ins_left[42] ,
    \ces_2_3_io_ins_left[41] ,
    \ces_2_3_io_ins_left[40] ,
    \ces_2_3_io_ins_left[39] ,
    \ces_2_3_io_ins_left[38] ,
    \ces_2_3_io_ins_left[37] ,
    \ces_2_3_io_ins_left[36] ,
    \ces_2_3_io_ins_left[35] ,
    \ces_2_3_io_ins_left[34] ,
    \ces_2_3_io_ins_left[33] ,
    \ces_2_3_io_ins_left[32] ,
    \ces_2_3_io_ins_left[31] ,
    \ces_2_3_io_ins_left[30] ,
    \ces_2_3_io_ins_left[29] ,
    \ces_2_3_io_ins_left[28] ,
    \ces_2_3_io_ins_left[27] ,
    \ces_2_3_io_ins_left[26] ,
    \ces_2_3_io_ins_left[25] ,
    \ces_2_3_io_ins_left[24] ,
    \ces_2_3_io_ins_left[23] ,
    \ces_2_3_io_ins_left[22] ,
    \ces_2_3_io_ins_left[21] ,
    \ces_2_3_io_ins_left[20] ,
    \ces_2_3_io_ins_left[19] ,
    \ces_2_3_io_ins_left[18] ,
    \ces_2_3_io_ins_left[17] ,
    \ces_2_3_io_ins_left[16] ,
    \ces_2_3_io_ins_left[15] ,
    \ces_2_3_io_ins_left[14] ,
    \ces_2_3_io_ins_left[13] ,
    \ces_2_3_io_ins_left[12] ,
    \ces_2_3_io_ins_left[11] ,
    \ces_2_3_io_ins_left[10] ,
    \ces_2_3_io_ins_left[9] ,
    \ces_2_3_io_ins_left[8] ,
    \ces_2_3_io_ins_left[7] ,
    \ces_2_3_io_ins_left[6] ,
    \ces_2_3_io_ins_left[5] ,
    \ces_2_3_io_ins_left[4] ,
    \ces_2_3_io_ins_left[3] ,
    \ces_2_3_io_ins_left[2] ,
    \ces_2_3_io_ins_left[1] ,
    \ces_2_3_io_ins_left[0] }),
    .io_ins_right({\ces_2_2_io_outs_right[63] ,
    \ces_2_2_io_outs_right[62] ,
    \ces_2_2_io_outs_right[61] ,
    \ces_2_2_io_outs_right[60] ,
    \ces_2_2_io_outs_right[59] ,
    \ces_2_2_io_outs_right[58] ,
    \ces_2_2_io_outs_right[57] ,
    \ces_2_2_io_outs_right[56] ,
    \ces_2_2_io_outs_right[55] ,
    \ces_2_2_io_outs_right[54] ,
    \ces_2_2_io_outs_right[53] ,
    \ces_2_2_io_outs_right[52] ,
    \ces_2_2_io_outs_right[51] ,
    \ces_2_2_io_outs_right[50] ,
    \ces_2_2_io_outs_right[49] ,
    \ces_2_2_io_outs_right[48] ,
    \ces_2_2_io_outs_right[47] ,
    \ces_2_2_io_outs_right[46] ,
    \ces_2_2_io_outs_right[45] ,
    \ces_2_2_io_outs_right[44] ,
    \ces_2_2_io_outs_right[43] ,
    \ces_2_2_io_outs_right[42] ,
    \ces_2_2_io_outs_right[41] ,
    \ces_2_2_io_outs_right[40] ,
    \ces_2_2_io_outs_right[39] ,
    \ces_2_2_io_outs_right[38] ,
    \ces_2_2_io_outs_right[37] ,
    \ces_2_2_io_outs_right[36] ,
    \ces_2_2_io_outs_right[35] ,
    \ces_2_2_io_outs_right[34] ,
    \ces_2_2_io_outs_right[33] ,
    \ces_2_2_io_outs_right[32] ,
    \ces_2_2_io_outs_right[31] ,
    \ces_2_2_io_outs_right[30] ,
    \ces_2_2_io_outs_right[29] ,
    \ces_2_2_io_outs_right[28] ,
    \ces_2_2_io_outs_right[27] ,
    \ces_2_2_io_outs_right[26] ,
    \ces_2_2_io_outs_right[25] ,
    \ces_2_2_io_outs_right[24] ,
    \ces_2_2_io_outs_right[23] ,
    \ces_2_2_io_outs_right[22] ,
    \ces_2_2_io_outs_right[21] ,
    \ces_2_2_io_outs_right[20] ,
    \ces_2_2_io_outs_right[19] ,
    \ces_2_2_io_outs_right[18] ,
    \ces_2_2_io_outs_right[17] ,
    \ces_2_2_io_outs_right[16] ,
    \ces_2_2_io_outs_right[15] ,
    \ces_2_2_io_outs_right[14] ,
    \ces_2_2_io_outs_right[13] ,
    \ces_2_2_io_outs_right[12] ,
    \ces_2_2_io_outs_right[11] ,
    \ces_2_2_io_outs_right[10] ,
    \ces_2_2_io_outs_right[9] ,
    \ces_2_2_io_outs_right[8] ,
    \ces_2_2_io_outs_right[7] ,
    \ces_2_2_io_outs_right[6] ,
    \ces_2_2_io_outs_right[5] ,
    \ces_2_2_io_outs_right[4] ,
    \ces_2_2_io_outs_right[3] ,
    \ces_2_2_io_outs_right[2] ,
    \ces_2_2_io_outs_right[1] ,
    \ces_2_2_io_outs_right[0] }),
    .io_ins_up({\ces_1_3_io_outs_up[63] ,
    \ces_1_3_io_outs_up[62] ,
    \ces_1_3_io_outs_up[61] ,
    \ces_1_3_io_outs_up[60] ,
    \ces_1_3_io_outs_up[59] ,
    \ces_1_3_io_outs_up[58] ,
    \ces_1_3_io_outs_up[57] ,
    \ces_1_3_io_outs_up[56] ,
    \ces_1_3_io_outs_up[55] ,
    \ces_1_3_io_outs_up[54] ,
    \ces_1_3_io_outs_up[53] ,
    \ces_1_3_io_outs_up[52] ,
    \ces_1_3_io_outs_up[51] ,
    \ces_1_3_io_outs_up[50] ,
    \ces_1_3_io_outs_up[49] ,
    \ces_1_3_io_outs_up[48] ,
    \ces_1_3_io_outs_up[47] ,
    \ces_1_3_io_outs_up[46] ,
    \ces_1_3_io_outs_up[45] ,
    \ces_1_3_io_outs_up[44] ,
    \ces_1_3_io_outs_up[43] ,
    \ces_1_3_io_outs_up[42] ,
    \ces_1_3_io_outs_up[41] ,
    \ces_1_3_io_outs_up[40] ,
    \ces_1_3_io_outs_up[39] ,
    \ces_1_3_io_outs_up[38] ,
    \ces_1_3_io_outs_up[37] ,
    \ces_1_3_io_outs_up[36] ,
    \ces_1_3_io_outs_up[35] ,
    \ces_1_3_io_outs_up[34] ,
    \ces_1_3_io_outs_up[33] ,
    \ces_1_3_io_outs_up[32] ,
    \ces_1_3_io_outs_up[31] ,
    \ces_1_3_io_outs_up[30] ,
    \ces_1_3_io_outs_up[29] ,
    \ces_1_3_io_outs_up[28] ,
    \ces_1_3_io_outs_up[27] ,
    \ces_1_3_io_outs_up[26] ,
    \ces_1_3_io_outs_up[25] ,
    \ces_1_3_io_outs_up[24] ,
    \ces_1_3_io_outs_up[23] ,
    \ces_1_3_io_outs_up[22] ,
    \ces_1_3_io_outs_up[21] ,
    \ces_1_3_io_outs_up[20] ,
    \ces_1_3_io_outs_up[19] ,
    \ces_1_3_io_outs_up[18] ,
    \ces_1_3_io_outs_up[17] ,
    \ces_1_3_io_outs_up[16] ,
    \ces_1_3_io_outs_up[15] ,
    \ces_1_3_io_outs_up[14] ,
    \ces_1_3_io_outs_up[13] ,
    \ces_1_3_io_outs_up[12] ,
    \ces_1_3_io_outs_up[11] ,
    \ces_1_3_io_outs_up[10] ,
    \ces_1_3_io_outs_up[9] ,
    \ces_1_3_io_outs_up[8] ,
    \ces_1_3_io_outs_up[7] ,
    \ces_1_3_io_outs_up[6] ,
    \ces_1_3_io_outs_up[5] ,
    \ces_1_3_io_outs_up[4] ,
    \ces_1_3_io_outs_up[3] ,
    \ces_1_3_io_outs_up[2] ,
    \ces_1_3_io_outs_up[1] ,
    \ces_1_3_io_outs_up[0] }),
    .io_outs_down({\ces_1_3_io_ins_down[63] ,
    \ces_1_3_io_ins_down[62] ,
    \ces_1_3_io_ins_down[61] ,
    \ces_1_3_io_ins_down[60] ,
    \ces_1_3_io_ins_down[59] ,
    \ces_1_3_io_ins_down[58] ,
    \ces_1_3_io_ins_down[57] ,
    \ces_1_3_io_ins_down[56] ,
    \ces_1_3_io_ins_down[55] ,
    \ces_1_3_io_ins_down[54] ,
    \ces_1_3_io_ins_down[53] ,
    \ces_1_3_io_ins_down[52] ,
    \ces_1_3_io_ins_down[51] ,
    \ces_1_3_io_ins_down[50] ,
    \ces_1_3_io_ins_down[49] ,
    \ces_1_3_io_ins_down[48] ,
    \ces_1_3_io_ins_down[47] ,
    \ces_1_3_io_ins_down[46] ,
    \ces_1_3_io_ins_down[45] ,
    \ces_1_3_io_ins_down[44] ,
    \ces_1_3_io_ins_down[43] ,
    \ces_1_3_io_ins_down[42] ,
    \ces_1_3_io_ins_down[41] ,
    \ces_1_3_io_ins_down[40] ,
    \ces_1_3_io_ins_down[39] ,
    \ces_1_3_io_ins_down[38] ,
    \ces_1_3_io_ins_down[37] ,
    \ces_1_3_io_ins_down[36] ,
    \ces_1_3_io_ins_down[35] ,
    \ces_1_3_io_ins_down[34] ,
    \ces_1_3_io_ins_down[33] ,
    \ces_1_3_io_ins_down[32] ,
    \ces_1_3_io_ins_down[31] ,
    \ces_1_3_io_ins_down[30] ,
    \ces_1_3_io_ins_down[29] ,
    \ces_1_3_io_ins_down[28] ,
    \ces_1_3_io_ins_down[27] ,
    \ces_1_3_io_ins_down[26] ,
    \ces_1_3_io_ins_down[25] ,
    \ces_1_3_io_ins_down[24] ,
    \ces_1_3_io_ins_down[23] ,
    \ces_1_3_io_ins_down[22] ,
    \ces_1_3_io_ins_down[21] ,
    \ces_1_3_io_ins_down[20] ,
    \ces_1_3_io_ins_down[19] ,
    \ces_1_3_io_ins_down[18] ,
    \ces_1_3_io_ins_down[17] ,
    \ces_1_3_io_ins_down[16] ,
    \ces_1_3_io_ins_down[15] ,
    \ces_1_3_io_ins_down[14] ,
    \ces_1_3_io_ins_down[13] ,
    \ces_1_3_io_ins_down[12] ,
    \ces_1_3_io_ins_down[11] ,
    \ces_1_3_io_ins_down[10] ,
    \ces_1_3_io_ins_down[9] ,
    \ces_1_3_io_ins_down[8] ,
    \ces_1_3_io_ins_down[7] ,
    \ces_1_3_io_ins_down[6] ,
    \ces_1_3_io_ins_down[5] ,
    \ces_1_3_io_ins_down[4] ,
    \ces_1_3_io_ins_down[3] ,
    \ces_1_3_io_ins_down[2] ,
    \ces_1_3_io_ins_down[1] ,
    \ces_1_3_io_ins_down[0] }),
    .io_outs_left({\ces_2_2_io_ins_left[63] ,
    \ces_2_2_io_ins_left[62] ,
    \ces_2_2_io_ins_left[61] ,
    \ces_2_2_io_ins_left[60] ,
    \ces_2_2_io_ins_left[59] ,
    \ces_2_2_io_ins_left[58] ,
    \ces_2_2_io_ins_left[57] ,
    \ces_2_2_io_ins_left[56] ,
    \ces_2_2_io_ins_left[55] ,
    \ces_2_2_io_ins_left[54] ,
    \ces_2_2_io_ins_left[53] ,
    \ces_2_2_io_ins_left[52] ,
    \ces_2_2_io_ins_left[51] ,
    \ces_2_2_io_ins_left[50] ,
    \ces_2_2_io_ins_left[49] ,
    \ces_2_2_io_ins_left[48] ,
    \ces_2_2_io_ins_left[47] ,
    \ces_2_2_io_ins_left[46] ,
    \ces_2_2_io_ins_left[45] ,
    \ces_2_2_io_ins_left[44] ,
    \ces_2_2_io_ins_left[43] ,
    \ces_2_2_io_ins_left[42] ,
    \ces_2_2_io_ins_left[41] ,
    \ces_2_2_io_ins_left[40] ,
    \ces_2_2_io_ins_left[39] ,
    \ces_2_2_io_ins_left[38] ,
    \ces_2_2_io_ins_left[37] ,
    \ces_2_2_io_ins_left[36] ,
    \ces_2_2_io_ins_left[35] ,
    \ces_2_2_io_ins_left[34] ,
    \ces_2_2_io_ins_left[33] ,
    \ces_2_2_io_ins_left[32] ,
    \ces_2_2_io_ins_left[31] ,
    \ces_2_2_io_ins_left[30] ,
    \ces_2_2_io_ins_left[29] ,
    \ces_2_2_io_ins_left[28] ,
    \ces_2_2_io_ins_left[27] ,
    \ces_2_2_io_ins_left[26] ,
    \ces_2_2_io_ins_left[25] ,
    \ces_2_2_io_ins_left[24] ,
    \ces_2_2_io_ins_left[23] ,
    \ces_2_2_io_ins_left[22] ,
    \ces_2_2_io_ins_left[21] ,
    \ces_2_2_io_ins_left[20] ,
    \ces_2_2_io_ins_left[19] ,
    \ces_2_2_io_ins_left[18] ,
    \ces_2_2_io_ins_left[17] ,
    \ces_2_2_io_ins_left[16] ,
    \ces_2_2_io_ins_left[15] ,
    \ces_2_2_io_ins_left[14] ,
    \ces_2_2_io_ins_left[13] ,
    \ces_2_2_io_ins_left[12] ,
    \ces_2_2_io_ins_left[11] ,
    \ces_2_2_io_ins_left[10] ,
    \ces_2_2_io_ins_left[9] ,
    \ces_2_2_io_ins_left[8] ,
    \ces_2_2_io_ins_left[7] ,
    \ces_2_2_io_ins_left[6] ,
    \ces_2_2_io_ins_left[5] ,
    \ces_2_2_io_ins_left[4] ,
    \ces_2_2_io_ins_left[3] ,
    \ces_2_2_io_ins_left[2] ,
    \ces_2_2_io_ins_left[1] ,
    \ces_2_2_io_ins_left[0] }),
    .io_outs_right({\ces_2_3_io_outs_right[63] ,
    \ces_2_3_io_outs_right[62] ,
    \ces_2_3_io_outs_right[61] ,
    \ces_2_3_io_outs_right[60] ,
    \ces_2_3_io_outs_right[59] ,
    \ces_2_3_io_outs_right[58] ,
    \ces_2_3_io_outs_right[57] ,
    \ces_2_3_io_outs_right[56] ,
    \ces_2_3_io_outs_right[55] ,
    \ces_2_3_io_outs_right[54] ,
    \ces_2_3_io_outs_right[53] ,
    \ces_2_3_io_outs_right[52] ,
    \ces_2_3_io_outs_right[51] ,
    \ces_2_3_io_outs_right[50] ,
    \ces_2_3_io_outs_right[49] ,
    \ces_2_3_io_outs_right[48] ,
    \ces_2_3_io_outs_right[47] ,
    \ces_2_3_io_outs_right[46] ,
    \ces_2_3_io_outs_right[45] ,
    \ces_2_3_io_outs_right[44] ,
    \ces_2_3_io_outs_right[43] ,
    \ces_2_3_io_outs_right[42] ,
    \ces_2_3_io_outs_right[41] ,
    \ces_2_3_io_outs_right[40] ,
    \ces_2_3_io_outs_right[39] ,
    \ces_2_3_io_outs_right[38] ,
    \ces_2_3_io_outs_right[37] ,
    \ces_2_3_io_outs_right[36] ,
    \ces_2_3_io_outs_right[35] ,
    \ces_2_3_io_outs_right[34] ,
    \ces_2_3_io_outs_right[33] ,
    \ces_2_3_io_outs_right[32] ,
    \ces_2_3_io_outs_right[31] ,
    \ces_2_3_io_outs_right[30] ,
    \ces_2_3_io_outs_right[29] ,
    \ces_2_3_io_outs_right[28] ,
    \ces_2_3_io_outs_right[27] ,
    \ces_2_3_io_outs_right[26] ,
    \ces_2_3_io_outs_right[25] ,
    \ces_2_3_io_outs_right[24] ,
    \ces_2_3_io_outs_right[23] ,
    \ces_2_3_io_outs_right[22] ,
    \ces_2_3_io_outs_right[21] ,
    \ces_2_3_io_outs_right[20] ,
    \ces_2_3_io_outs_right[19] ,
    \ces_2_3_io_outs_right[18] ,
    \ces_2_3_io_outs_right[17] ,
    \ces_2_3_io_outs_right[16] ,
    \ces_2_3_io_outs_right[15] ,
    \ces_2_3_io_outs_right[14] ,
    \ces_2_3_io_outs_right[13] ,
    \ces_2_3_io_outs_right[12] ,
    \ces_2_3_io_outs_right[11] ,
    \ces_2_3_io_outs_right[10] ,
    \ces_2_3_io_outs_right[9] ,
    \ces_2_3_io_outs_right[8] ,
    \ces_2_3_io_outs_right[7] ,
    \ces_2_3_io_outs_right[6] ,
    \ces_2_3_io_outs_right[5] ,
    \ces_2_3_io_outs_right[4] ,
    \ces_2_3_io_outs_right[3] ,
    \ces_2_3_io_outs_right[2] ,
    \ces_2_3_io_outs_right[1] ,
    \ces_2_3_io_outs_right[0] }),
    .io_outs_up({\ces_2_3_io_outs_up[63] ,
    \ces_2_3_io_outs_up[62] ,
    \ces_2_3_io_outs_up[61] ,
    \ces_2_3_io_outs_up[60] ,
    \ces_2_3_io_outs_up[59] ,
    \ces_2_3_io_outs_up[58] ,
    \ces_2_3_io_outs_up[57] ,
    \ces_2_3_io_outs_up[56] ,
    \ces_2_3_io_outs_up[55] ,
    \ces_2_3_io_outs_up[54] ,
    \ces_2_3_io_outs_up[53] ,
    \ces_2_3_io_outs_up[52] ,
    \ces_2_3_io_outs_up[51] ,
    \ces_2_3_io_outs_up[50] ,
    \ces_2_3_io_outs_up[49] ,
    \ces_2_3_io_outs_up[48] ,
    \ces_2_3_io_outs_up[47] ,
    \ces_2_3_io_outs_up[46] ,
    \ces_2_3_io_outs_up[45] ,
    \ces_2_3_io_outs_up[44] ,
    \ces_2_3_io_outs_up[43] ,
    \ces_2_3_io_outs_up[42] ,
    \ces_2_3_io_outs_up[41] ,
    \ces_2_3_io_outs_up[40] ,
    \ces_2_3_io_outs_up[39] ,
    \ces_2_3_io_outs_up[38] ,
    \ces_2_3_io_outs_up[37] ,
    \ces_2_3_io_outs_up[36] ,
    \ces_2_3_io_outs_up[35] ,
    \ces_2_3_io_outs_up[34] ,
    \ces_2_3_io_outs_up[33] ,
    \ces_2_3_io_outs_up[32] ,
    \ces_2_3_io_outs_up[31] ,
    \ces_2_3_io_outs_up[30] ,
    \ces_2_3_io_outs_up[29] ,
    \ces_2_3_io_outs_up[28] ,
    \ces_2_3_io_outs_up[27] ,
    \ces_2_3_io_outs_up[26] ,
    \ces_2_3_io_outs_up[25] ,
    \ces_2_3_io_outs_up[24] ,
    \ces_2_3_io_outs_up[23] ,
    \ces_2_3_io_outs_up[22] ,
    \ces_2_3_io_outs_up[21] ,
    \ces_2_3_io_outs_up[20] ,
    \ces_2_3_io_outs_up[19] ,
    \ces_2_3_io_outs_up[18] ,
    \ces_2_3_io_outs_up[17] ,
    \ces_2_3_io_outs_up[16] ,
    \ces_2_3_io_outs_up[15] ,
    \ces_2_3_io_outs_up[14] ,
    \ces_2_3_io_outs_up[13] ,
    \ces_2_3_io_outs_up[12] ,
    \ces_2_3_io_outs_up[11] ,
    \ces_2_3_io_outs_up[10] ,
    \ces_2_3_io_outs_up[9] ,
    \ces_2_3_io_outs_up[8] ,
    \ces_2_3_io_outs_up[7] ,
    \ces_2_3_io_outs_up[6] ,
    \ces_2_3_io_outs_up[5] ,
    \ces_2_3_io_outs_up[4] ,
    \ces_2_3_io_outs_up[3] ,
    \ces_2_3_io_outs_up[2] ,
    \ces_2_3_io_outs_up[1] ,
    \ces_2_3_io_outs_up[0] }));
 Element ces_2_4 (.clock(clknet_3_3_0_clock),
    .io_lsbIns_1(ces_2_3_io_lsbOuts_1),
    .io_lsbIns_2(ces_2_3_io_lsbOuts_2),
    .io_lsbIns_3(ces_2_3_io_lsbOuts_3),
    .io_lsbIns_4(ces_2_3_io_lsbOuts_4),
    .io_lsbIns_5(ces_2_3_io_lsbOuts_5),
    .io_lsbIns_6(ces_2_3_io_lsbOuts_6),
    .io_lsbIns_7(ces_2_3_io_lsbOuts_7),
    .io_lsbOuts_0(ces_2_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_4_io_lsbOuts_7),
    .io_ins_down({\ces_2_4_io_ins_down[63] ,
    \ces_2_4_io_ins_down[62] ,
    \ces_2_4_io_ins_down[61] ,
    \ces_2_4_io_ins_down[60] ,
    \ces_2_4_io_ins_down[59] ,
    \ces_2_4_io_ins_down[58] ,
    \ces_2_4_io_ins_down[57] ,
    \ces_2_4_io_ins_down[56] ,
    \ces_2_4_io_ins_down[55] ,
    \ces_2_4_io_ins_down[54] ,
    \ces_2_4_io_ins_down[53] ,
    \ces_2_4_io_ins_down[52] ,
    \ces_2_4_io_ins_down[51] ,
    \ces_2_4_io_ins_down[50] ,
    \ces_2_4_io_ins_down[49] ,
    \ces_2_4_io_ins_down[48] ,
    \ces_2_4_io_ins_down[47] ,
    \ces_2_4_io_ins_down[46] ,
    \ces_2_4_io_ins_down[45] ,
    \ces_2_4_io_ins_down[44] ,
    \ces_2_4_io_ins_down[43] ,
    \ces_2_4_io_ins_down[42] ,
    \ces_2_4_io_ins_down[41] ,
    \ces_2_4_io_ins_down[40] ,
    \ces_2_4_io_ins_down[39] ,
    \ces_2_4_io_ins_down[38] ,
    \ces_2_4_io_ins_down[37] ,
    \ces_2_4_io_ins_down[36] ,
    \ces_2_4_io_ins_down[35] ,
    \ces_2_4_io_ins_down[34] ,
    \ces_2_4_io_ins_down[33] ,
    \ces_2_4_io_ins_down[32] ,
    \ces_2_4_io_ins_down[31] ,
    \ces_2_4_io_ins_down[30] ,
    \ces_2_4_io_ins_down[29] ,
    \ces_2_4_io_ins_down[28] ,
    \ces_2_4_io_ins_down[27] ,
    \ces_2_4_io_ins_down[26] ,
    \ces_2_4_io_ins_down[25] ,
    \ces_2_4_io_ins_down[24] ,
    \ces_2_4_io_ins_down[23] ,
    \ces_2_4_io_ins_down[22] ,
    \ces_2_4_io_ins_down[21] ,
    \ces_2_4_io_ins_down[20] ,
    \ces_2_4_io_ins_down[19] ,
    \ces_2_4_io_ins_down[18] ,
    \ces_2_4_io_ins_down[17] ,
    \ces_2_4_io_ins_down[16] ,
    \ces_2_4_io_ins_down[15] ,
    \ces_2_4_io_ins_down[14] ,
    \ces_2_4_io_ins_down[13] ,
    \ces_2_4_io_ins_down[12] ,
    \ces_2_4_io_ins_down[11] ,
    \ces_2_4_io_ins_down[10] ,
    \ces_2_4_io_ins_down[9] ,
    \ces_2_4_io_ins_down[8] ,
    \ces_2_4_io_ins_down[7] ,
    \ces_2_4_io_ins_down[6] ,
    \ces_2_4_io_ins_down[5] ,
    \ces_2_4_io_ins_down[4] ,
    \ces_2_4_io_ins_down[3] ,
    \ces_2_4_io_ins_down[2] ,
    \ces_2_4_io_ins_down[1] ,
    \ces_2_4_io_ins_down[0] }),
    .io_ins_left({\ces_2_4_io_ins_left[63] ,
    \ces_2_4_io_ins_left[62] ,
    \ces_2_4_io_ins_left[61] ,
    \ces_2_4_io_ins_left[60] ,
    \ces_2_4_io_ins_left[59] ,
    \ces_2_4_io_ins_left[58] ,
    \ces_2_4_io_ins_left[57] ,
    \ces_2_4_io_ins_left[56] ,
    \ces_2_4_io_ins_left[55] ,
    \ces_2_4_io_ins_left[54] ,
    \ces_2_4_io_ins_left[53] ,
    \ces_2_4_io_ins_left[52] ,
    \ces_2_4_io_ins_left[51] ,
    \ces_2_4_io_ins_left[50] ,
    \ces_2_4_io_ins_left[49] ,
    \ces_2_4_io_ins_left[48] ,
    \ces_2_4_io_ins_left[47] ,
    \ces_2_4_io_ins_left[46] ,
    \ces_2_4_io_ins_left[45] ,
    \ces_2_4_io_ins_left[44] ,
    \ces_2_4_io_ins_left[43] ,
    \ces_2_4_io_ins_left[42] ,
    \ces_2_4_io_ins_left[41] ,
    \ces_2_4_io_ins_left[40] ,
    \ces_2_4_io_ins_left[39] ,
    \ces_2_4_io_ins_left[38] ,
    \ces_2_4_io_ins_left[37] ,
    \ces_2_4_io_ins_left[36] ,
    \ces_2_4_io_ins_left[35] ,
    \ces_2_4_io_ins_left[34] ,
    \ces_2_4_io_ins_left[33] ,
    \ces_2_4_io_ins_left[32] ,
    \ces_2_4_io_ins_left[31] ,
    \ces_2_4_io_ins_left[30] ,
    \ces_2_4_io_ins_left[29] ,
    \ces_2_4_io_ins_left[28] ,
    \ces_2_4_io_ins_left[27] ,
    \ces_2_4_io_ins_left[26] ,
    \ces_2_4_io_ins_left[25] ,
    \ces_2_4_io_ins_left[24] ,
    \ces_2_4_io_ins_left[23] ,
    \ces_2_4_io_ins_left[22] ,
    \ces_2_4_io_ins_left[21] ,
    \ces_2_4_io_ins_left[20] ,
    \ces_2_4_io_ins_left[19] ,
    \ces_2_4_io_ins_left[18] ,
    \ces_2_4_io_ins_left[17] ,
    \ces_2_4_io_ins_left[16] ,
    \ces_2_4_io_ins_left[15] ,
    \ces_2_4_io_ins_left[14] ,
    \ces_2_4_io_ins_left[13] ,
    \ces_2_4_io_ins_left[12] ,
    \ces_2_4_io_ins_left[11] ,
    \ces_2_4_io_ins_left[10] ,
    \ces_2_4_io_ins_left[9] ,
    \ces_2_4_io_ins_left[8] ,
    \ces_2_4_io_ins_left[7] ,
    \ces_2_4_io_ins_left[6] ,
    \ces_2_4_io_ins_left[5] ,
    \ces_2_4_io_ins_left[4] ,
    \ces_2_4_io_ins_left[3] ,
    \ces_2_4_io_ins_left[2] ,
    \ces_2_4_io_ins_left[1] ,
    \ces_2_4_io_ins_left[0] }),
    .io_ins_right({\ces_2_3_io_outs_right[63] ,
    \ces_2_3_io_outs_right[62] ,
    \ces_2_3_io_outs_right[61] ,
    \ces_2_3_io_outs_right[60] ,
    \ces_2_3_io_outs_right[59] ,
    \ces_2_3_io_outs_right[58] ,
    \ces_2_3_io_outs_right[57] ,
    \ces_2_3_io_outs_right[56] ,
    \ces_2_3_io_outs_right[55] ,
    \ces_2_3_io_outs_right[54] ,
    \ces_2_3_io_outs_right[53] ,
    \ces_2_3_io_outs_right[52] ,
    \ces_2_3_io_outs_right[51] ,
    \ces_2_3_io_outs_right[50] ,
    \ces_2_3_io_outs_right[49] ,
    \ces_2_3_io_outs_right[48] ,
    \ces_2_3_io_outs_right[47] ,
    \ces_2_3_io_outs_right[46] ,
    \ces_2_3_io_outs_right[45] ,
    \ces_2_3_io_outs_right[44] ,
    \ces_2_3_io_outs_right[43] ,
    \ces_2_3_io_outs_right[42] ,
    \ces_2_3_io_outs_right[41] ,
    \ces_2_3_io_outs_right[40] ,
    \ces_2_3_io_outs_right[39] ,
    \ces_2_3_io_outs_right[38] ,
    \ces_2_3_io_outs_right[37] ,
    \ces_2_3_io_outs_right[36] ,
    \ces_2_3_io_outs_right[35] ,
    \ces_2_3_io_outs_right[34] ,
    \ces_2_3_io_outs_right[33] ,
    \ces_2_3_io_outs_right[32] ,
    \ces_2_3_io_outs_right[31] ,
    \ces_2_3_io_outs_right[30] ,
    \ces_2_3_io_outs_right[29] ,
    \ces_2_3_io_outs_right[28] ,
    \ces_2_3_io_outs_right[27] ,
    \ces_2_3_io_outs_right[26] ,
    \ces_2_3_io_outs_right[25] ,
    \ces_2_3_io_outs_right[24] ,
    \ces_2_3_io_outs_right[23] ,
    \ces_2_3_io_outs_right[22] ,
    \ces_2_3_io_outs_right[21] ,
    \ces_2_3_io_outs_right[20] ,
    \ces_2_3_io_outs_right[19] ,
    \ces_2_3_io_outs_right[18] ,
    \ces_2_3_io_outs_right[17] ,
    \ces_2_3_io_outs_right[16] ,
    \ces_2_3_io_outs_right[15] ,
    \ces_2_3_io_outs_right[14] ,
    \ces_2_3_io_outs_right[13] ,
    \ces_2_3_io_outs_right[12] ,
    \ces_2_3_io_outs_right[11] ,
    \ces_2_3_io_outs_right[10] ,
    \ces_2_3_io_outs_right[9] ,
    \ces_2_3_io_outs_right[8] ,
    \ces_2_3_io_outs_right[7] ,
    \ces_2_3_io_outs_right[6] ,
    \ces_2_3_io_outs_right[5] ,
    \ces_2_3_io_outs_right[4] ,
    \ces_2_3_io_outs_right[3] ,
    \ces_2_3_io_outs_right[2] ,
    \ces_2_3_io_outs_right[1] ,
    \ces_2_3_io_outs_right[0] }),
    .io_ins_up({\ces_1_4_io_outs_up[63] ,
    \ces_1_4_io_outs_up[62] ,
    \ces_1_4_io_outs_up[61] ,
    \ces_1_4_io_outs_up[60] ,
    \ces_1_4_io_outs_up[59] ,
    \ces_1_4_io_outs_up[58] ,
    \ces_1_4_io_outs_up[57] ,
    \ces_1_4_io_outs_up[56] ,
    \ces_1_4_io_outs_up[55] ,
    \ces_1_4_io_outs_up[54] ,
    \ces_1_4_io_outs_up[53] ,
    \ces_1_4_io_outs_up[52] ,
    \ces_1_4_io_outs_up[51] ,
    \ces_1_4_io_outs_up[50] ,
    \ces_1_4_io_outs_up[49] ,
    \ces_1_4_io_outs_up[48] ,
    \ces_1_4_io_outs_up[47] ,
    \ces_1_4_io_outs_up[46] ,
    \ces_1_4_io_outs_up[45] ,
    \ces_1_4_io_outs_up[44] ,
    \ces_1_4_io_outs_up[43] ,
    \ces_1_4_io_outs_up[42] ,
    \ces_1_4_io_outs_up[41] ,
    \ces_1_4_io_outs_up[40] ,
    \ces_1_4_io_outs_up[39] ,
    \ces_1_4_io_outs_up[38] ,
    \ces_1_4_io_outs_up[37] ,
    \ces_1_4_io_outs_up[36] ,
    \ces_1_4_io_outs_up[35] ,
    \ces_1_4_io_outs_up[34] ,
    \ces_1_4_io_outs_up[33] ,
    \ces_1_4_io_outs_up[32] ,
    \ces_1_4_io_outs_up[31] ,
    \ces_1_4_io_outs_up[30] ,
    \ces_1_4_io_outs_up[29] ,
    \ces_1_4_io_outs_up[28] ,
    \ces_1_4_io_outs_up[27] ,
    \ces_1_4_io_outs_up[26] ,
    \ces_1_4_io_outs_up[25] ,
    \ces_1_4_io_outs_up[24] ,
    \ces_1_4_io_outs_up[23] ,
    \ces_1_4_io_outs_up[22] ,
    \ces_1_4_io_outs_up[21] ,
    \ces_1_4_io_outs_up[20] ,
    \ces_1_4_io_outs_up[19] ,
    \ces_1_4_io_outs_up[18] ,
    \ces_1_4_io_outs_up[17] ,
    \ces_1_4_io_outs_up[16] ,
    \ces_1_4_io_outs_up[15] ,
    \ces_1_4_io_outs_up[14] ,
    \ces_1_4_io_outs_up[13] ,
    \ces_1_4_io_outs_up[12] ,
    \ces_1_4_io_outs_up[11] ,
    \ces_1_4_io_outs_up[10] ,
    \ces_1_4_io_outs_up[9] ,
    \ces_1_4_io_outs_up[8] ,
    \ces_1_4_io_outs_up[7] ,
    \ces_1_4_io_outs_up[6] ,
    \ces_1_4_io_outs_up[5] ,
    \ces_1_4_io_outs_up[4] ,
    \ces_1_4_io_outs_up[3] ,
    \ces_1_4_io_outs_up[2] ,
    \ces_1_4_io_outs_up[1] ,
    \ces_1_4_io_outs_up[0] }),
    .io_outs_down({\ces_1_4_io_ins_down[63] ,
    \ces_1_4_io_ins_down[62] ,
    \ces_1_4_io_ins_down[61] ,
    \ces_1_4_io_ins_down[60] ,
    \ces_1_4_io_ins_down[59] ,
    \ces_1_4_io_ins_down[58] ,
    \ces_1_4_io_ins_down[57] ,
    \ces_1_4_io_ins_down[56] ,
    \ces_1_4_io_ins_down[55] ,
    \ces_1_4_io_ins_down[54] ,
    \ces_1_4_io_ins_down[53] ,
    \ces_1_4_io_ins_down[52] ,
    \ces_1_4_io_ins_down[51] ,
    \ces_1_4_io_ins_down[50] ,
    \ces_1_4_io_ins_down[49] ,
    \ces_1_4_io_ins_down[48] ,
    \ces_1_4_io_ins_down[47] ,
    \ces_1_4_io_ins_down[46] ,
    \ces_1_4_io_ins_down[45] ,
    \ces_1_4_io_ins_down[44] ,
    \ces_1_4_io_ins_down[43] ,
    \ces_1_4_io_ins_down[42] ,
    \ces_1_4_io_ins_down[41] ,
    \ces_1_4_io_ins_down[40] ,
    \ces_1_4_io_ins_down[39] ,
    \ces_1_4_io_ins_down[38] ,
    \ces_1_4_io_ins_down[37] ,
    \ces_1_4_io_ins_down[36] ,
    \ces_1_4_io_ins_down[35] ,
    \ces_1_4_io_ins_down[34] ,
    \ces_1_4_io_ins_down[33] ,
    \ces_1_4_io_ins_down[32] ,
    \ces_1_4_io_ins_down[31] ,
    \ces_1_4_io_ins_down[30] ,
    \ces_1_4_io_ins_down[29] ,
    \ces_1_4_io_ins_down[28] ,
    \ces_1_4_io_ins_down[27] ,
    \ces_1_4_io_ins_down[26] ,
    \ces_1_4_io_ins_down[25] ,
    \ces_1_4_io_ins_down[24] ,
    \ces_1_4_io_ins_down[23] ,
    \ces_1_4_io_ins_down[22] ,
    \ces_1_4_io_ins_down[21] ,
    \ces_1_4_io_ins_down[20] ,
    \ces_1_4_io_ins_down[19] ,
    \ces_1_4_io_ins_down[18] ,
    \ces_1_4_io_ins_down[17] ,
    \ces_1_4_io_ins_down[16] ,
    \ces_1_4_io_ins_down[15] ,
    \ces_1_4_io_ins_down[14] ,
    \ces_1_4_io_ins_down[13] ,
    \ces_1_4_io_ins_down[12] ,
    \ces_1_4_io_ins_down[11] ,
    \ces_1_4_io_ins_down[10] ,
    \ces_1_4_io_ins_down[9] ,
    \ces_1_4_io_ins_down[8] ,
    \ces_1_4_io_ins_down[7] ,
    \ces_1_4_io_ins_down[6] ,
    \ces_1_4_io_ins_down[5] ,
    \ces_1_4_io_ins_down[4] ,
    \ces_1_4_io_ins_down[3] ,
    \ces_1_4_io_ins_down[2] ,
    \ces_1_4_io_ins_down[1] ,
    \ces_1_4_io_ins_down[0] }),
    .io_outs_left({\ces_2_3_io_ins_left[63] ,
    \ces_2_3_io_ins_left[62] ,
    \ces_2_3_io_ins_left[61] ,
    \ces_2_3_io_ins_left[60] ,
    \ces_2_3_io_ins_left[59] ,
    \ces_2_3_io_ins_left[58] ,
    \ces_2_3_io_ins_left[57] ,
    \ces_2_3_io_ins_left[56] ,
    \ces_2_3_io_ins_left[55] ,
    \ces_2_3_io_ins_left[54] ,
    \ces_2_3_io_ins_left[53] ,
    \ces_2_3_io_ins_left[52] ,
    \ces_2_3_io_ins_left[51] ,
    \ces_2_3_io_ins_left[50] ,
    \ces_2_3_io_ins_left[49] ,
    \ces_2_3_io_ins_left[48] ,
    \ces_2_3_io_ins_left[47] ,
    \ces_2_3_io_ins_left[46] ,
    \ces_2_3_io_ins_left[45] ,
    \ces_2_3_io_ins_left[44] ,
    \ces_2_3_io_ins_left[43] ,
    \ces_2_3_io_ins_left[42] ,
    \ces_2_3_io_ins_left[41] ,
    \ces_2_3_io_ins_left[40] ,
    \ces_2_3_io_ins_left[39] ,
    \ces_2_3_io_ins_left[38] ,
    \ces_2_3_io_ins_left[37] ,
    \ces_2_3_io_ins_left[36] ,
    \ces_2_3_io_ins_left[35] ,
    \ces_2_3_io_ins_left[34] ,
    \ces_2_3_io_ins_left[33] ,
    \ces_2_3_io_ins_left[32] ,
    \ces_2_3_io_ins_left[31] ,
    \ces_2_3_io_ins_left[30] ,
    \ces_2_3_io_ins_left[29] ,
    \ces_2_3_io_ins_left[28] ,
    \ces_2_3_io_ins_left[27] ,
    \ces_2_3_io_ins_left[26] ,
    \ces_2_3_io_ins_left[25] ,
    \ces_2_3_io_ins_left[24] ,
    \ces_2_3_io_ins_left[23] ,
    \ces_2_3_io_ins_left[22] ,
    \ces_2_3_io_ins_left[21] ,
    \ces_2_3_io_ins_left[20] ,
    \ces_2_3_io_ins_left[19] ,
    \ces_2_3_io_ins_left[18] ,
    \ces_2_3_io_ins_left[17] ,
    \ces_2_3_io_ins_left[16] ,
    \ces_2_3_io_ins_left[15] ,
    \ces_2_3_io_ins_left[14] ,
    \ces_2_3_io_ins_left[13] ,
    \ces_2_3_io_ins_left[12] ,
    \ces_2_3_io_ins_left[11] ,
    \ces_2_3_io_ins_left[10] ,
    \ces_2_3_io_ins_left[9] ,
    \ces_2_3_io_ins_left[8] ,
    \ces_2_3_io_ins_left[7] ,
    \ces_2_3_io_ins_left[6] ,
    \ces_2_3_io_ins_left[5] ,
    \ces_2_3_io_ins_left[4] ,
    \ces_2_3_io_ins_left[3] ,
    \ces_2_3_io_ins_left[2] ,
    \ces_2_3_io_ins_left[1] ,
    \ces_2_3_io_ins_left[0] }),
    .io_outs_right({\ces_2_4_io_outs_right[63] ,
    \ces_2_4_io_outs_right[62] ,
    \ces_2_4_io_outs_right[61] ,
    \ces_2_4_io_outs_right[60] ,
    \ces_2_4_io_outs_right[59] ,
    \ces_2_4_io_outs_right[58] ,
    \ces_2_4_io_outs_right[57] ,
    \ces_2_4_io_outs_right[56] ,
    \ces_2_4_io_outs_right[55] ,
    \ces_2_4_io_outs_right[54] ,
    \ces_2_4_io_outs_right[53] ,
    \ces_2_4_io_outs_right[52] ,
    \ces_2_4_io_outs_right[51] ,
    \ces_2_4_io_outs_right[50] ,
    \ces_2_4_io_outs_right[49] ,
    \ces_2_4_io_outs_right[48] ,
    \ces_2_4_io_outs_right[47] ,
    \ces_2_4_io_outs_right[46] ,
    \ces_2_4_io_outs_right[45] ,
    \ces_2_4_io_outs_right[44] ,
    \ces_2_4_io_outs_right[43] ,
    \ces_2_4_io_outs_right[42] ,
    \ces_2_4_io_outs_right[41] ,
    \ces_2_4_io_outs_right[40] ,
    \ces_2_4_io_outs_right[39] ,
    \ces_2_4_io_outs_right[38] ,
    \ces_2_4_io_outs_right[37] ,
    \ces_2_4_io_outs_right[36] ,
    \ces_2_4_io_outs_right[35] ,
    \ces_2_4_io_outs_right[34] ,
    \ces_2_4_io_outs_right[33] ,
    \ces_2_4_io_outs_right[32] ,
    \ces_2_4_io_outs_right[31] ,
    \ces_2_4_io_outs_right[30] ,
    \ces_2_4_io_outs_right[29] ,
    \ces_2_4_io_outs_right[28] ,
    \ces_2_4_io_outs_right[27] ,
    \ces_2_4_io_outs_right[26] ,
    \ces_2_4_io_outs_right[25] ,
    \ces_2_4_io_outs_right[24] ,
    \ces_2_4_io_outs_right[23] ,
    \ces_2_4_io_outs_right[22] ,
    \ces_2_4_io_outs_right[21] ,
    \ces_2_4_io_outs_right[20] ,
    \ces_2_4_io_outs_right[19] ,
    \ces_2_4_io_outs_right[18] ,
    \ces_2_4_io_outs_right[17] ,
    \ces_2_4_io_outs_right[16] ,
    \ces_2_4_io_outs_right[15] ,
    \ces_2_4_io_outs_right[14] ,
    \ces_2_4_io_outs_right[13] ,
    \ces_2_4_io_outs_right[12] ,
    \ces_2_4_io_outs_right[11] ,
    \ces_2_4_io_outs_right[10] ,
    \ces_2_4_io_outs_right[9] ,
    \ces_2_4_io_outs_right[8] ,
    \ces_2_4_io_outs_right[7] ,
    \ces_2_4_io_outs_right[6] ,
    \ces_2_4_io_outs_right[5] ,
    \ces_2_4_io_outs_right[4] ,
    \ces_2_4_io_outs_right[3] ,
    \ces_2_4_io_outs_right[2] ,
    \ces_2_4_io_outs_right[1] ,
    \ces_2_4_io_outs_right[0] }),
    .io_outs_up({\ces_2_4_io_outs_up[63] ,
    \ces_2_4_io_outs_up[62] ,
    \ces_2_4_io_outs_up[61] ,
    \ces_2_4_io_outs_up[60] ,
    \ces_2_4_io_outs_up[59] ,
    \ces_2_4_io_outs_up[58] ,
    \ces_2_4_io_outs_up[57] ,
    \ces_2_4_io_outs_up[56] ,
    \ces_2_4_io_outs_up[55] ,
    \ces_2_4_io_outs_up[54] ,
    \ces_2_4_io_outs_up[53] ,
    \ces_2_4_io_outs_up[52] ,
    \ces_2_4_io_outs_up[51] ,
    \ces_2_4_io_outs_up[50] ,
    \ces_2_4_io_outs_up[49] ,
    \ces_2_4_io_outs_up[48] ,
    \ces_2_4_io_outs_up[47] ,
    \ces_2_4_io_outs_up[46] ,
    \ces_2_4_io_outs_up[45] ,
    \ces_2_4_io_outs_up[44] ,
    \ces_2_4_io_outs_up[43] ,
    \ces_2_4_io_outs_up[42] ,
    \ces_2_4_io_outs_up[41] ,
    \ces_2_4_io_outs_up[40] ,
    \ces_2_4_io_outs_up[39] ,
    \ces_2_4_io_outs_up[38] ,
    \ces_2_4_io_outs_up[37] ,
    \ces_2_4_io_outs_up[36] ,
    \ces_2_4_io_outs_up[35] ,
    \ces_2_4_io_outs_up[34] ,
    \ces_2_4_io_outs_up[33] ,
    \ces_2_4_io_outs_up[32] ,
    \ces_2_4_io_outs_up[31] ,
    \ces_2_4_io_outs_up[30] ,
    \ces_2_4_io_outs_up[29] ,
    \ces_2_4_io_outs_up[28] ,
    \ces_2_4_io_outs_up[27] ,
    \ces_2_4_io_outs_up[26] ,
    \ces_2_4_io_outs_up[25] ,
    \ces_2_4_io_outs_up[24] ,
    \ces_2_4_io_outs_up[23] ,
    \ces_2_4_io_outs_up[22] ,
    \ces_2_4_io_outs_up[21] ,
    \ces_2_4_io_outs_up[20] ,
    \ces_2_4_io_outs_up[19] ,
    \ces_2_4_io_outs_up[18] ,
    \ces_2_4_io_outs_up[17] ,
    \ces_2_4_io_outs_up[16] ,
    \ces_2_4_io_outs_up[15] ,
    \ces_2_4_io_outs_up[14] ,
    \ces_2_4_io_outs_up[13] ,
    \ces_2_4_io_outs_up[12] ,
    \ces_2_4_io_outs_up[11] ,
    \ces_2_4_io_outs_up[10] ,
    \ces_2_4_io_outs_up[9] ,
    \ces_2_4_io_outs_up[8] ,
    \ces_2_4_io_outs_up[7] ,
    \ces_2_4_io_outs_up[6] ,
    \ces_2_4_io_outs_up[5] ,
    \ces_2_4_io_outs_up[4] ,
    \ces_2_4_io_outs_up[3] ,
    \ces_2_4_io_outs_up[2] ,
    \ces_2_4_io_outs_up[1] ,
    \ces_2_4_io_outs_up[0] }));
 Element ces_2_5 (.clock(clknet_3_3_0_clock),
    .io_lsbIns_1(ces_2_4_io_lsbOuts_1),
    .io_lsbIns_2(ces_2_4_io_lsbOuts_2),
    .io_lsbIns_3(ces_2_4_io_lsbOuts_3),
    .io_lsbIns_4(ces_2_4_io_lsbOuts_4),
    .io_lsbIns_5(ces_2_4_io_lsbOuts_5),
    .io_lsbIns_6(ces_2_4_io_lsbOuts_6),
    .io_lsbIns_7(ces_2_4_io_lsbOuts_7),
    .io_lsbOuts_0(ces_2_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_5_io_lsbOuts_7),
    .io_ins_down({\ces_2_5_io_ins_down[63] ,
    \ces_2_5_io_ins_down[62] ,
    \ces_2_5_io_ins_down[61] ,
    \ces_2_5_io_ins_down[60] ,
    \ces_2_5_io_ins_down[59] ,
    \ces_2_5_io_ins_down[58] ,
    \ces_2_5_io_ins_down[57] ,
    \ces_2_5_io_ins_down[56] ,
    \ces_2_5_io_ins_down[55] ,
    \ces_2_5_io_ins_down[54] ,
    \ces_2_5_io_ins_down[53] ,
    \ces_2_5_io_ins_down[52] ,
    \ces_2_5_io_ins_down[51] ,
    \ces_2_5_io_ins_down[50] ,
    \ces_2_5_io_ins_down[49] ,
    \ces_2_5_io_ins_down[48] ,
    \ces_2_5_io_ins_down[47] ,
    \ces_2_5_io_ins_down[46] ,
    \ces_2_5_io_ins_down[45] ,
    \ces_2_5_io_ins_down[44] ,
    \ces_2_5_io_ins_down[43] ,
    \ces_2_5_io_ins_down[42] ,
    \ces_2_5_io_ins_down[41] ,
    \ces_2_5_io_ins_down[40] ,
    \ces_2_5_io_ins_down[39] ,
    \ces_2_5_io_ins_down[38] ,
    \ces_2_5_io_ins_down[37] ,
    \ces_2_5_io_ins_down[36] ,
    \ces_2_5_io_ins_down[35] ,
    \ces_2_5_io_ins_down[34] ,
    \ces_2_5_io_ins_down[33] ,
    \ces_2_5_io_ins_down[32] ,
    \ces_2_5_io_ins_down[31] ,
    \ces_2_5_io_ins_down[30] ,
    \ces_2_5_io_ins_down[29] ,
    \ces_2_5_io_ins_down[28] ,
    \ces_2_5_io_ins_down[27] ,
    \ces_2_5_io_ins_down[26] ,
    \ces_2_5_io_ins_down[25] ,
    \ces_2_5_io_ins_down[24] ,
    \ces_2_5_io_ins_down[23] ,
    \ces_2_5_io_ins_down[22] ,
    \ces_2_5_io_ins_down[21] ,
    \ces_2_5_io_ins_down[20] ,
    \ces_2_5_io_ins_down[19] ,
    \ces_2_5_io_ins_down[18] ,
    \ces_2_5_io_ins_down[17] ,
    \ces_2_5_io_ins_down[16] ,
    \ces_2_5_io_ins_down[15] ,
    \ces_2_5_io_ins_down[14] ,
    \ces_2_5_io_ins_down[13] ,
    \ces_2_5_io_ins_down[12] ,
    \ces_2_5_io_ins_down[11] ,
    \ces_2_5_io_ins_down[10] ,
    \ces_2_5_io_ins_down[9] ,
    \ces_2_5_io_ins_down[8] ,
    \ces_2_5_io_ins_down[7] ,
    \ces_2_5_io_ins_down[6] ,
    \ces_2_5_io_ins_down[5] ,
    \ces_2_5_io_ins_down[4] ,
    \ces_2_5_io_ins_down[3] ,
    \ces_2_5_io_ins_down[2] ,
    \ces_2_5_io_ins_down[1] ,
    \ces_2_5_io_ins_down[0] }),
    .io_ins_left({\ces_2_5_io_ins_left[63] ,
    \ces_2_5_io_ins_left[62] ,
    \ces_2_5_io_ins_left[61] ,
    \ces_2_5_io_ins_left[60] ,
    \ces_2_5_io_ins_left[59] ,
    \ces_2_5_io_ins_left[58] ,
    \ces_2_5_io_ins_left[57] ,
    \ces_2_5_io_ins_left[56] ,
    \ces_2_5_io_ins_left[55] ,
    \ces_2_5_io_ins_left[54] ,
    \ces_2_5_io_ins_left[53] ,
    \ces_2_5_io_ins_left[52] ,
    \ces_2_5_io_ins_left[51] ,
    \ces_2_5_io_ins_left[50] ,
    \ces_2_5_io_ins_left[49] ,
    \ces_2_5_io_ins_left[48] ,
    \ces_2_5_io_ins_left[47] ,
    \ces_2_5_io_ins_left[46] ,
    \ces_2_5_io_ins_left[45] ,
    \ces_2_5_io_ins_left[44] ,
    \ces_2_5_io_ins_left[43] ,
    \ces_2_5_io_ins_left[42] ,
    \ces_2_5_io_ins_left[41] ,
    \ces_2_5_io_ins_left[40] ,
    \ces_2_5_io_ins_left[39] ,
    \ces_2_5_io_ins_left[38] ,
    \ces_2_5_io_ins_left[37] ,
    \ces_2_5_io_ins_left[36] ,
    \ces_2_5_io_ins_left[35] ,
    \ces_2_5_io_ins_left[34] ,
    \ces_2_5_io_ins_left[33] ,
    \ces_2_5_io_ins_left[32] ,
    \ces_2_5_io_ins_left[31] ,
    \ces_2_5_io_ins_left[30] ,
    \ces_2_5_io_ins_left[29] ,
    \ces_2_5_io_ins_left[28] ,
    \ces_2_5_io_ins_left[27] ,
    \ces_2_5_io_ins_left[26] ,
    \ces_2_5_io_ins_left[25] ,
    \ces_2_5_io_ins_left[24] ,
    \ces_2_5_io_ins_left[23] ,
    \ces_2_5_io_ins_left[22] ,
    \ces_2_5_io_ins_left[21] ,
    \ces_2_5_io_ins_left[20] ,
    \ces_2_5_io_ins_left[19] ,
    \ces_2_5_io_ins_left[18] ,
    \ces_2_5_io_ins_left[17] ,
    \ces_2_5_io_ins_left[16] ,
    \ces_2_5_io_ins_left[15] ,
    \ces_2_5_io_ins_left[14] ,
    \ces_2_5_io_ins_left[13] ,
    \ces_2_5_io_ins_left[12] ,
    \ces_2_5_io_ins_left[11] ,
    \ces_2_5_io_ins_left[10] ,
    \ces_2_5_io_ins_left[9] ,
    \ces_2_5_io_ins_left[8] ,
    \ces_2_5_io_ins_left[7] ,
    \ces_2_5_io_ins_left[6] ,
    \ces_2_5_io_ins_left[5] ,
    \ces_2_5_io_ins_left[4] ,
    \ces_2_5_io_ins_left[3] ,
    \ces_2_5_io_ins_left[2] ,
    \ces_2_5_io_ins_left[1] ,
    \ces_2_5_io_ins_left[0] }),
    .io_ins_right({\ces_2_4_io_outs_right[63] ,
    \ces_2_4_io_outs_right[62] ,
    \ces_2_4_io_outs_right[61] ,
    \ces_2_4_io_outs_right[60] ,
    \ces_2_4_io_outs_right[59] ,
    \ces_2_4_io_outs_right[58] ,
    \ces_2_4_io_outs_right[57] ,
    \ces_2_4_io_outs_right[56] ,
    \ces_2_4_io_outs_right[55] ,
    \ces_2_4_io_outs_right[54] ,
    \ces_2_4_io_outs_right[53] ,
    \ces_2_4_io_outs_right[52] ,
    \ces_2_4_io_outs_right[51] ,
    \ces_2_4_io_outs_right[50] ,
    \ces_2_4_io_outs_right[49] ,
    \ces_2_4_io_outs_right[48] ,
    \ces_2_4_io_outs_right[47] ,
    \ces_2_4_io_outs_right[46] ,
    \ces_2_4_io_outs_right[45] ,
    \ces_2_4_io_outs_right[44] ,
    \ces_2_4_io_outs_right[43] ,
    \ces_2_4_io_outs_right[42] ,
    \ces_2_4_io_outs_right[41] ,
    \ces_2_4_io_outs_right[40] ,
    \ces_2_4_io_outs_right[39] ,
    \ces_2_4_io_outs_right[38] ,
    \ces_2_4_io_outs_right[37] ,
    \ces_2_4_io_outs_right[36] ,
    \ces_2_4_io_outs_right[35] ,
    \ces_2_4_io_outs_right[34] ,
    \ces_2_4_io_outs_right[33] ,
    \ces_2_4_io_outs_right[32] ,
    \ces_2_4_io_outs_right[31] ,
    \ces_2_4_io_outs_right[30] ,
    \ces_2_4_io_outs_right[29] ,
    \ces_2_4_io_outs_right[28] ,
    \ces_2_4_io_outs_right[27] ,
    \ces_2_4_io_outs_right[26] ,
    \ces_2_4_io_outs_right[25] ,
    \ces_2_4_io_outs_right[24] ,
    \ces_2_4_io_outs_right[23] ,
    \ces_2_4_io_outs_right[22] ,
    \ces_2_4_io_outs_right[21] ,
    \ces_2_4_io_outs_right[20] ,
    \ces_2_4_io_outs_right[19] ,
    \ces_2_4_io_outs_right[18] ,
    \ces_2_4_io_outs_right[17] ,
    \ces_2_4_io_outs_right[16] ,
    \ces_2_4_io_outs_right[15] ,
    \ces_2_4_io_outs_right[14] ,
    \ces_2_4_io_outs_right[13] ,
    \ces_2_4_io_outs_right[12] ,
    \ces_2_4_io_outs_right[11] ,
    \ces_2_4_io_outs_right[10] ,
    \ces_2_4_io_outs_right[9] ,
    \ces_2_4_io_outs_right[8] ,
    \ces_2_4_io_outs_right[7] ,
    \ces_2_4_io_outs_right[6] ,
    \ces_2_4_io_outs_right[5] ,
    \ces_2_4_io_outs_right[4] ,
    \ces_2_4_io_outs_right[3] ,
    \ces_2_4_io_outs_right[2] ,
    \ces_2_4_io_outs_right[1] ,
    \ces_2_4_io_outs_right[0] }),
    .io_ins_up({\ces_1_5_io_outs_up[63] ,
    \ces_1_5_io_outs_up[62] ,
    \ces_1_5_io_outs_up[61] ,
    \ces_1_5_io_outs_up[60] ,
    \ces_1_5_io_outs_up[59] ,
    \ces_1_5_io_outs_up[58] ,
    \ces_1_5_io_outs_up[57] ,
    \ces_1_5_io_outs_up[56] ,
    \ces_1_5_io_outs_up[55] ,
    \ces_1_5_io_outs_up[54] ,
    \ces_1_5_io_outs_up[53] ,
    \ces_1_5_io_outs_up[52] ,
    \ces_1_5_io_outs_up[51] ,
    \ces_1_5_io_outs_up[50] ,
    \ces_1_5_io_outs_up[49] ,
    \ces_1_5_io_outs_up[48] ,
    \ces_1_5_io_outs_up[47] ,
    \ces_1_5_io_outs_up[46] ,
    \ces_1_5_io_outs_up[45] ,
    \ces_1_5_io_outs_up[44] ,
    \ces_1_5_io_outs_up[43] ,
    \ces_1_5_io_outs_up[42] ,
    \ces_1_5_io_outs_up[41] ,
    \ces_1_5_io_outs_up[40] ,
    \ces_1_5_io_outs_up[39] ,
    \ces_1_5_io_outs_up[38] ,
    \ces_1_5_io_outs_up[37] ,
    \ces_1_5_io_outs_up[36] ,
    \ces_1_5_io_outs_up[35] ,
    \ces_1_5_io_outs_up[34] ,
    \ces_1_5_io_outs_up[33] ,
    \ces_1_5_io_outs_up[32] ,
    \ces_1_5_io_outs_up[31] ,
    \ces_1_5_io_outs_up[30] ,
    \ces_1_5_io_outs_up[29] ,
    \ces_1_5_io_outs_up[28] ,
    \ces_1_5_io_outs_up[27] ,
    \ces_1_5_io_outs_up[26] ,
    \ces_1_5_io_outs_up[25] ,
    \ces_1_5_io_outs_up[24] ,
    \ces_1_5_io_outs_up[23] ,
    \ces_1_5_io_outs_up[22] ,
    \ces_1_5_io_outs_up[21] ,
    \ces_1_5_io_outs_up[20] ,
    \ces_1_5_io_outs_up[19] ,
    \ces_1_5_io_outs_up[18] ,
    \ces_1_5_io_outs_up[17] ,
    \ces_1_5_io_outs_up[16] ,
    \ces_1_5_io_outs_up[15] ,
    \ces_1_5_io_outs_up[14] ,
    \ces_1_5_io_outs_up[13] ,
    \ces_1_5_io_outs_up[12] ,
    \ces_1_5_io_outs_up[11] ,
    \ces_1_5_io_outs_up[10] ,
    \ces_1_5_io_outs_up[9] ,
    \ces_1_5_io_outs_up[8] ,
    \ces_1_5_io_outs_up[7] ,
    \ces_1_5_io_outs_up[6] ,
    \ces_1_5_io_outs_up[5] ,
    \ces_1_5_io_outs_up[4] ,
    \ces_1_5_io_outs_up[3] ,
    \ces_1_5_io_outs_up[2] ,
    \ces_1_5_io_outs_up[1] ,
    \ces_1_5_io_outs_up[0] }),
    .io_outs_down({\ces_1_5_io_ins_down[63] ,
    \ces_1_5_io_ins_down[62] ,
    \ces_1_5_io_ins_down[61] ,
    \ces_1_5_io_ins_down[60] ,
    \ces_1_5_io_ins_down[59] ,
    \ces_1_5_io_ins_down[58] ,
    \ces_1_5_io_ins_down[57] ,
    \ces_1_5_io_ins_down[56] ,
    \ces_1_5_io_ins_down[55] ,
    \ces_1_5_io_ins_down[54] ,
    \ces_1_5_io_ins_down[53] ,
    \ces_1_5_io_ins_down[52] ,
    \ces_1_5_io_ins_down[51] ,
    \ces_1_5_io_ins_down[50] ,
    \ces_1_5_io_ins_down[49] ,
    \ces_1_5_io_ins_down[48] ,
    \ces_1_5_io_ins_down[47] ,
    \ces_1_5_io_ins_down[46] ,
    \ces_1_5_io_ins_down[45] ,
    \ces_1_5_io_ins_down[44] ,
    \ces_1_5_io_ins_down[43] ,
    \ces_1_5_io_ins_down[42] ,
    \ces_1_5_io_ins_down[41] ,
    \ces_1_5_io_ins_down[40] ,
    \ces_1_5_io_ins_down[39] ,
    \ces_1_5_io_ins_down[38] ,
    \ces_1_5_io_ins_down[37] ,
    \ces_1_5_io_ins_down[36] ,
    \ces_1_5_io_ins_down[35] ,
    \ces_1_5_io_ins_down[34] ,
    \ces_1_5_io_ins_down[33] ,
    \ces_1_5_io_ins_down[32] ,
    \ces_1_5_io_ins_down[31] ,
    \ces_1_5_io_ins_down[30] ,
    \ces_1_5_io_ins_down[29] ,
    \ces_1_5_io_ins_down[28] ,
    \ces_1_5_io_ins_down[27] ,
    \ces_1_5_io_ins_down[26] ,
    \ces_1_5_io_ins_down[25] ,
    \ces_1_5_io_ins_down[24] ,
    \ces_1_5_io_ins_down[23] ,
    \ces_1_5_io_ins_down[22] ,
    \ces_1_5_io_ins_down[21] ,
    \ces_1_5_io_ins_down[20] ,
    \ces_1_5_io_ins_down[19] ,
    \ces_1_5_io_ins_down[18] ,
    \ces_1_5_io_ins_down[17] ,
    \ces_1_5_io_ins_down[16] ,
    \ces_1_5_io_ins_down[15] ,
    \ces_1_5_io_ins_down[14] ,
    \ces_1_5_io_ins_down[13] ,
    \ces_1_5_io_ins_down[12] ,
    \ces_1_5_io_ins_down[11] ,
    \ces_1_5_io_ins_down[10] ,
    \ces_1_5_io_ins_down[9] ,
    \ces_1_5_io_ins_down[8] ,
    \ces_1_5_io_ins_down[7] ,
    \ces_1_5_io_ins_down[6] ,
    \ces_1_5_io_ins_down[5] ,
    \ces_1_5_io_ins_down[4] ,
    \ces_1_5_io_ins_down[3] ,
    \ces_1_5_io_ins_down[2] ,
    \ces_1_5_io_ins_down[1] ,
    \ces_1_5_io_ins_down[0] }),
    .io_outs_left({\ces_2_4_io_ins_left[63] ,
    \ces_2_4_io_ins_left[62] ,
    \ces_2_4_io_ins_left[61] ,
    \ces_2_4_io_ins_left[60] ,
    \ces_2_4_io_ins_left[59] ,
    \ces_2_4_io_ins_left[58] ,
    \ces_2_4_io_ins_left[57] ,
    \ces_2_4_io_ins_left[56] ,
    \ces_2_4_io_ins_left[55] ,
    \ces_2_4_io_ins_left[54] ,
    \ces_2_4_io_ins_left[53] ,
    \ces_2_4_io_ins_left[52] ,
    \ces_2_4_io_ins_left[51] ,
    \ces_2_4_io_ins_left[50] ,
    \ces_2_4_io_ins_left[49] ,
    \ces_2_4_io_ins_left[48] ,
    \ces_2_4_io_ins_left[47] ,
    \ces_2_4_io_ins_left[46] ,
    \ces_2_4_io_ins_left[45] ,
    \ces_2_4_io_ins_left[44] ,
    \ces_2_4_io_ins_left[43] ,
    \ces_2_4_io_ins_left[42] ,
    \ces_2_4_io_ins_left[41] ,
    \ces_2_4_io_ins_left[40] ,
    \ces_2_4_io_ins_left[39] ,
    \ces_2_4_io_ins_left[38] ,
    \ces_2_4_io_ins_left[37] ,
    \ces_2_4_io_ins_left[36] ,
    \ces_2_4_io_ins_left[35] ,
    \ces_2_4_io_ins_left[34] ,
    \ces_2_4_io_ins_left[33] ,
    \ces_2_4_io_ins_left[32] ,
    \ces_2_4_io_ins_left[31] ,
    \ces_2_4_io_ins_left[30] ,
    \ces_2_4_io_ins_left[29] ,
    \ces_2_4_io_ins_left[28] ,
    \ces_2_4_io_ins_left[27] ,
    \ces_2_4_io_ins_left[26] ,
    \ces_2_4_io_ins_left[25] ,
    \ces_2_4_io_ins_left[24] ,
    \ces_2_4_io_ins_left[23] ,
    \ces_2_4_io_ins_left[22] ,
    \ces_2_4_io_ins_left[21] ,
    \ces_2_4_io_ins_left[20] ,
    \ces_2_4_io_ins_left[19] ,
    \ces_2_4_io_ins_left[18] ,
    \ces_2_4_io_ins_left[17] ,
    \ces_2_4_io_ins_left[16] ,
    \ces_2_4_io_ins_left[15] ,
    \ces_2_4_io_ins_left[14] ,
    \ces_2_4_io_ins_left[13] ,
    \ces_2_4_io_ins_left[12] ,
    \ces_2_4_io_ins_left[11] ,
    \ces_2_4_io_ins_left[10] ,
    \ces_2_4_io_ins_left[9] ,
    \ces_2_4_io_ins_left[8] ,
    \ces_2_4_io_ins_left[7] ,
    \ces_2_4_io_ins_left[6] ,
    \ces_2_4_io_ins_left[5] ,
    \ces_2_4_io_ins_left[4] ,
    \ces_2_4_io_ins_left[3] ,
    \ces_2_4_io_ins_left[2] ,
    \ces_2_4_io_ins_left[1] ,
    \ces_2_4_io_ins_left[0] }),
    .io_outs_right({\ces_2_5_io_outs_right[63] ,
    \ces_2_5_io_outs_right[62] ,
    \ces_2_5_io_outs_right[61] ,
    \ces_2_5_io_outs_right[60] ,
    \ces_2_5_io_outs_right[59] ,
    \ces_2_5_io_outs_right[58] ,
    \ces_2_5_io_outs_right[57] ,
    \ces_2_5_io_outs_right[56] ,
    \ces_2_5_io_outs_right[55] ,
    \ces_2_5_io_outs_right[54] ,
    \ces_2_5_io_outs_right[53] ,
    \ces_2_5_io_outs_right[52] ,
    \ces_2_5_io_outs_right[51] ,
    \ces_2_5_io_outs_right[50] ,
    \ces_2_5_io_outs_right[49] ,
    \ces_2_5_io_outs_right[48] ,
    \ces_2_5_io_outs_right[47] ,
    \ces_2_5_io_outs_right[46] ,
    \ces_2_5_io_outs_right[45] ,
    \ces_2_5_io_outs_right[44] ,
    \ces_2_5_io_outs_right[43] ,
    \ces_2_5_io_outs_right[42] ,
    \ces_2_5_io_outs_right[41] ,
    \ces_2_5_io_outs_right[40] ,
    \ces_2_5_io_outs_right[39] ,
    \ces_2_5_io_outs_right[38] ,
    \ces_2_5_io_outs_right[37] ,
    \ces_2_5_io_outs_right[36] ,
    \ces_2_5_io_outs_right[35] ,
    \ces_2_5_io_outs_right[34] ,
    \ces_2_5_io_outs_right[33] ,
    \ces_2_5_io_outs_right[32] ,
    \ces_2_5_io_outs_right[31] ,
    \ces_2_5_io_outs_right[30] ,
    \ces_2_5_io_outs_right[29] ,
    \ces_2_5_io_outs_right[28] ,
    \ces_2_5_io_outs_right[27] ,
    \ces_2_5_io_outs_right[26] ,
    \ces_2_5_io_outs_right[25] ,
    \ces_2_5_io_outs_right[24] ,
    \ces_2_5_io_outs_right[23] ,
    \ces_2_5_io_outs_right[22] ,
    \ces_2_5_io_outs_right[21] ,
    \ces_2_5_io_outs_right[20] ,
    \ces_2_5_io_outs_right[19] ,
    \ces_2_5_io_outs_right[18] ,
    \ces_2_5_io_outs_right[17] ,
    \ces_2_5_io_outs_right[16] ,
    \ces_2_5_io_outs_right[15] ,
    \ces_2_5_io_outs_right[14] ,
    \ces_2_5_io_outs_right[13] ,
    \ces_2_5_io_outs_right[12] ,
    \ces_2_5_io_outs_right[11] ,
    \ces_2_5_io_outs_right[10] ,
    \ces_2_5_io_outs_right[9] ,
    \ces_2_5_io_outs_right[8] ,
    \ces_2_5_io_outs_right[7] ,
    \ces_2_5_io_outs_right[6] ,
    \ces_2_5_io_outs_right[5] ,
    \ces_2_5_io_outs_right[4] ,
    \ces_2_5_io_outs_right[3] ,
    \ces_2_5_io_outs_right[2] ,
    \ces_2_5_io_outs_right[1] ,
    \ces_2_5_io_outs_right[0] }),
    .io_outs_up({\ces_2_5_io_outs_up[63] ,
    \ces_2_5_io_outs_up[62] ,
    \ces_2_5_io_outs_up[61] ,
    \ces_2_5_io_outs_up[60] ,
    \ces_2_5_io_outs_up[59] ,
    \ces_2_5_io_outs_up[58] ,
    \ces_2_5_io_outs_up[57] ,
    \ces_2_5_io_outs_up[56] ,
    \ces_2_5_io_outs_up[55] ,
    \ces_2_5_io_outs_up[54] ,
    \ces_2_5_io_outs_up[53] ,
    \ces_2_5_io_outs_up[52] ,
    \ces_2_5_io_outs_up[51] ,
    \ces_2_5_io_outs_up[50] ,
    \ces_2_5_io_outs_up[49] ,
    \ces_2_5_io_outs_up[48] ,
    \ces_2_5_io_outs_up[47] ,
    \ces_2_5_io_outs_up[46] ,
    \ces_2_5_io_outs_up[45] ,
    \ces_2_5_io_outs_up[44] ,
    \ces_2_5_io_outs_up[43] ,
    \ces_2_5_io_outs_up[42] ,
    \ces_2_5_io_outs_up[41] ,
    \ces_2_5_io_outs_up[40] ,
    \ces_2_5_io_outs_up[39] ,
    \ces_2_5_io_outs_up[38] ,
    \ces_2_5_io_outs_up[37] ,
    \ces_2_5_io_outs_up[36] ,
    \ces_2_5_io_outs_up[35] ,
    \ces_2_5_io_outs_up[34] ,
    \ces_2_5_io_outs_up[33] ,
    \ces_2_5_io_outs_up[32] ,
    \ces_2_5_io_outs_up[31] ,
    \ces_2_5_io_outs_up[30] ,
    \ces_2_5_io_outs_up[29] ,
    \ces_2_5_io_outs_up[28] ,
    \ces_2_5_io_outs_up[27] ,
    \ces_2_5_io_outs_up[26] ,
    \ces_2_5_io_outs_up[25] ,
    \ces_2_5_io_outs_up[24] ,
    \ces_2_5_io_outs_up[23] ,
    \ces_2_5_io_outs_up[22] ,
    \ces_2_5_io_outs_up[21] ,
    \ces_2_5_io_outs_up[20] ,
    \ces_2_5_io_outs_up[19] ,
    \ces_2_5_io_outs_up[18] ,
    \ces_2_5_io_outs_up[17] ,
    \ces_2_5_io_outs_up[16] ,
    \ces_2_5_io_outs_up[15] ,
    \ces_2_5_io_outs_up[14] ,
    \ces_2_5_io_outs_up[13] ,
    \ces_2_5_io_outs_up[12] ,
    \ces_2_5_io_outs_up[11] ,
    \ces_2_5_io_outs_up[10] ,
    \ces_2_5_io_outs_up[9] ,
    \ces_2_5_io_outs_up[8] ,
    \ces_2_5_io_outs_up[7] ,
    \ces_2_5_io_outs_up[6] ,
    \ces_2_5_io_outs_up[5] ,
    \ces_2_5_io_outs_up[4] ,
    \ces_2_5_io_outs_up[3] ,
    \ces_2_5_io_outs_up[2] ,
    \ces_2_5_io_outs_up[1] ,
    \ces_2_5_io_outs_up[0] }));
 Element ces_2_6 (.clock(clknet_3_3_0_clock),
    .io_lsbIns_1(ces_2_5_io_lsbOuts_1),
    .io_lsbIns_2(ces_2_5_io_lsbOuts_2),
    .io_lsbIns_3(ces_2_5_io_lsbOuts_3),
    .io_lsbIns_4(ces_2_5_io_lsbOuts_4),
    .io_lsbIns_5(ces_2_5_io_lsbOuts_5),
    .io_lsbIns_6(ces_2_5_io_lsbOuts_6),
    .io_lsbIns_7(ces_2_5_io_lsbOuts_7),
    .io_lsbOuts_0(ces_2_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_6_io_lsbOuts_7),
    .io_ins_down({\ces_2_6_io_ins_down[63] ,
    \ces_2_6_io_ins_down[62] ,
    \ces_2_6_io_ins_down[61] ,
    \ces_2_6_io_ins_down[60] ,
    \ces_2_6_io_ins_down[59] ,
    \ces_2_6_io_ins_down[58] ,
    \ces_2_6_io_ins_down[57] ,
    \ces_2_6_io_ins_down[56] ,
    \ces_2_6_io_ins_down[55] ,
    \ces_2_6_io_ins_down[54] ,
    \ces_2_6_io_ins_down[53] ,
    \ces_2_6_io_ins_down[52] ,
    \ces_2_6_io_ins_down[51] ,
    \ces_2_6_io_ins_down[50] ,
    \ces_2_6_io_ins_down[49] ,
    \ces_2_6_io_ins_down[48] ,
    \ces_2_6_io_ins_down[47] ,
    \ces_2_6_io_ins_down[46] ,
    \ces_2_6_io_ins_down[45] ,
    \ces_2_6_io_ins_down[44] ,
    \ces_2_6_io_ins_down[43] ,
    \ces_2_6_io_ins_down[42] ,
    \ces_2_6_io_ins_down[41] ,
    \ces_2_6_io_ins_down[40] ,
    \ces_2_6_io_ins_down[39] ,
    \ces_2_6_io_ins_down[38] ,
    \ces_2_6_io_ins_down[37] ,
    \ces_2_6_io_ins_down[36] ,
    \ces_2_6_io_ins_down[35] ,
    \ces_2_6_io_ins_down[34] ,
    \ces_2_6_io_ins_down[33] ,
    \ces_2_6_io_ins_down[32] ,
    \ces_2_6_io_ins_down[31] ,
    \ces_2_6_io_ins_down[30] ,
    \ces_2_6_io_ins_down[29] ,
    \ces_2_6_io_ins_down[28] ,
    \ces_2_6_io_ins_down[27] ,
    \ces_2_6_io_ins_down[26] ,
    \ces_2_6_io_ins_down[25] ,
    \ces_2_6_io_ins_down[24] ,
    \ces_2_6_io_ins_down[23] ,
    \ces_2_6_io_ins_down[22] ,
    \ces_2_6_io_ins_down[21] ,
    \ces_2_6_io_ins_down[20] ,
    \ces_2_6_io_ins_down[19] ,
    \ces_2_6_io_ins_down[18] ,
    \ces_2_6_io_ins_down[17] ,
    \ces_2_6_io_ins_down[16] ,
    \ces_2_6_io_ins_down[15] ,
    \ces_2_6_io_ins_down[14] ,
    \ces_2_6_io_ins_down[13] ,
    \ces_2_6_io_ins_down[12] ,
    \ces_2_6_io_ins_down[11] ,
    \ces_2_6_io_ins_down[10] ,
    \ces_2_6_io_ins_down[9] ,
    \ces_2_6_io_ins_down[8] ,
    \ces_2_6_io_ins_down[7] ,
    \ces_2_6_io_ins_down[6] ,
    \ces_2_6_io_ins_down[5] ,
    \ces_2_6_io_ins_down[4] ,
    \ces_2_6_io_ins_down[3] ,
    \ces_2_6_io_ins_down[2] ,
    \ces_2_6_io_ins_down[1] ,
    \ces_2_6_io_ins_down[0] }),
    .io_ins_left({\ces_2_6_io_ins_left[63] ,
    \ces_2_6_io_ins_left[62] ,
    \ces_2_6_io_ins_left[61] ,
    \ces_2_6_io_ins_left[60] ,
    \ces_2_6_io_ins_left[59] ,
    \ces_2_6_io_ins_left[58] ,
    \ces_2_6_io_ins_left[57] ,
    \ces_2_6_io_ins_left[56] ,
    \ces_2_6_io_ins_left[55] ,
    \ces_2_6_io_ins_left[54] ,
    \ces_2_6_io_ins_left[53] ,
    \ces_2_6_io_ins_left[52] ,
    \ces_2_6_io_ins_left[51] ,
    \ces_2_6_io_ins_left[50] ,
    \ces_2_6_io_ins_left[49] ,
    \ces_2_6_io_ins_left[48] ,
    \ces_2_6_io_ins_left[47] ,
    \ces_2_6_io_ins_left[46] ,
    \ces_2_6_io_ins_left[45] ,
    \ces_2_6_io_ins_left[44] ,
    \ces_2_6_io_ins_left[43] ,
    \ces_2_6_io_ins_left[42] ,
    \ces_2_6_io_ins_left[41] ,
    \ces_2_6_io_ins_left[40] ,
    \ces_2_6_io_ins_left[39] ,
    \ces_2_6_io_ins_left[38] ,
    \ces_2_6_io_ins_left[37] ,
    \ces_2_6_io_ins_left[36] ,
    \ces_2_6_io_ins_left[35] ,
    \ces_2_6_io_ins_left[34] ,
    \ces_2_6_io_ins_left[33] ,
    \ces_2_6_io_ins_left[32] ,
    \ces_2_6_io_ins_left[31] ,
    \ces_2_6_io_ins_left[30] ,
    \ces_2_6_io_ins_left[29] ,
    \ces_2_6_io_ins_left[28] ,
    \ces_2_6_io_ins_left[27] ,
    \ces_2_6_io_ins_left[26] ,
    \ces_2_6_io_ins_left[25] ,
    \ces_2_6_io_ins_left[24] ,
    \ces_2_6_io_ins_left[23] ,
    \ces_2_6_io_ins_left[22] ,
    \ces_2_6_io_ins_left[21] ,
    \ces_2_6_io_ins_left[20] ,
    \ces_2_6_io_ins_left[19] ,
    \ces_2_6_io_ins_left[18] ,
    \ces_2_6_io_ins_left[17] ,
    \ces_2_6_io_ins_left[16] ,
    \ces_2_6_io_ins_left[15] ,
    \ces_2_6_io_ins_left[14] ,
    \ces_2_6_io_ins_left[13] ,
    \ces_2_6_io_ins_left[12] ,
    \ces_2_6_io_ins_left[11] ,
    \ces_2_6_io_ins_left[10] ,
    \ces_2_6_io_ins_left[9] ,
    \ces_2_6_io_ins_left[8] ,
    \ces_2_6_io_ins_left[7] ,
    \ces_2_6_io_ins_left[6] ,
    \ces_2_6_io_ins_left[5] ,
    \ces_2_6_io_ins_left[4] ,
    \ces_2_6_io_ins_left[3] ,
    \ces_2_6_io_ins_left[2] ,
    \ces_2_6_io_ins_left[1] ,
    \ces_2_6_io_ins_left[0] }),
    .io_ins_right({\ces_2_5_io_outs_right[63] ,
    \ces_2_5_io_outs_right[62] ,
    \ces_2_5_io_outs_right[61] ,
    \ces_2_5_io_outs_right[60] ,
    \ces_2_5_io_outs_right[59] ,
    \ces_2_5_io_outs_right[58] ,
    \ces_2_5_io_outs_right[57] ,
    \ces_2_5_io_outs_right[56] ,
    \ces_2_5_io_outs_right[55] ,
    \ces_2_5_io_outs_right[54] ,
    \ces_2_5_io_outs_right[53] ,
    \ces_2_5_io_outs_right[52] ,
    \ces_2_5_io_outs_right[51] ,
    \ces_2_5_io_outs_right[50] ,
    \ces_2_5_io_outs_right[49] ,
    \ces_2_5_io_outs_right[48] ,
    \ces_2_5_io_outs_right[47] ,
    \ces_2_5_io_outs_right[46] ,
    \ces_2_5_io_outs_right[45] ,
    \ces_2_5_io_outs_right[44] ,
    \ces_2_5_io_outs_right[43] ,
    \ces_2_5_io_outs_right[42] ,
    \ces_2_5_io_outs_right[41] ,
    \ces_2_5_io_outs_right[40] ,
    \ces_2_5_io_outs_right[39] ,
    \ces_2_5_io_outs_right[38] ,
    \ces_2_5_io_outs_right[37] ,
    \ces_2_5_io_outs_right[36] ,
    \ces_2_5_io_outs_right[35] ,
    \ces_2_5_io_outs_right[34] ,
    \ces_2_5_io_outs_right[33] ,
    \ces_2_5_io_outs_right[32] ,
    \ces_2_5_io_outs_right[31] ,
    \ces_2_5_io_outs_right[30] ,
    \ces_2_5_io_outs_right[29] ,
    \ces_2_5_io_outs_right[28] ,
    \ces_2_5_io_outs_right[27] ,
    \ces_2_5_io_outs_right[26] ,
    \ces_2_5_io_outs_right[25] ,
    \ces_2_5_io_outs_right[24] ,
    \ces_2_5_io_outs_right[23] ,
    \ces_2_5_io_outs_right[22] ,
    \ces_2_5_io_outs_right[21] ,
    \ces_2_5_io_outs_right[20] ,
    \ces_2_5_io_outs_right[19] ,
    \ces_2_5_io_outs_right[18] ,
    \ces_2_5_io_outs_right[17] ,
    \ces_2_5_io_outs_right[16] ,
    \ces_2_5_io_outs_right[15] ,
    \ces_2_5_io_outs_right[14] ,
    \ces_2_5_io_outs_right[13] ,
    \ces_2_5_io_outs_right[12] ,
    \ces_2_5_io_outs_right[11] ,
    \ces_2_5_io_outs_right[10] ,
    \ces_2_5_io_outs_right[9] ,
    \ces_2_5_io_outs_right[8] ,
    \ces_2_5_io_outs_right[7] ,
    \ces_2_5_io_outs_right[6] ,
    \ces_2_5_io_outs_right[5] ,
    \ces_2_5_io_outs_right[4] ,
    \ces_2_5_io_outs_right[3] ,
    \ces_2_5_io_outs_right[2] ,
    \ces_2_5_io_outs_right[1] ,
    \ces_2_5_io_outs_right[0] }),
    .io_ins_up({\ces_1_6_io_outs_up[63] ,
    \ces_1_6_io_outs_up[62] ,
    \ces_1_6_io_outs_up[61] ,
    \ces_1_6_io_outs_up[60] ,
    \ces_1_6_io_outs_up[59] ,
    \ces_1_6_io_outs_up[58] ,
    \ces_1_6_io_outs_up[57] ,
    \ces_1_6_io_outs_up[56] ,
    \ces_1_6_io_outs_up[55] ,
    \ces_1_6_io_outs_up[54] ,
    \ces_1_6_io_outs_up[53] ,
    \ces_1_6_io_outs_up[52] ,
    \ces_1_6_io_outs_up[51] ,
    \ces_1_6_io_outs_up[50] ,
    \ces_1_6_io_outs_up[49] ,
    \ces_1_6_io_outs_up[48] ,
    \ces_1_6_io_outs_up[47] ,
    \ces_1_6_io_outs_up[46] ,
    \ces_1_6_io_outs_up[45] ,
    \ces_1_6_io_outs_up[44] ,
    \ces_1_6_io_outs_up[43] ,
    \ces_1_6_io_outs_up[42] ,
    \ces_1_6_io_outs_up[41] ,
    \ces_1_6_io_outs_up[40] ,
    \ces_1_6_io_outs_up[39] ,
    \ces_1_6_io_outs_up[38] ,
    \ces_1_6_io_outs_up[37] ,
    \ces_1_6_io_outs_up[36] ,
    \ces_1_6_io_outs_up[35] ,
    \ces_1_6_io_outs_up[34] ,
    \ces_1_6_io_outs_up[33] ,
    \ces_1_6_io_outs_up[32] ,
    \ces_1_6_io_outs_up[31] ,
    \ces_1_6_io_outs_up[30] ,
    \ces_1_6_io_outs_up[29] ,
    \ces_1_6_io_outs_up[28] ,
    \ces_1_6_io_outs_up[27] ,
    \ces_1_6_io_outs_up[26] ,
    \ces_1_6_io_outs_up[25] ,
    \ces_1_6_io_outs_up[24] ,
    \ces_1_6_io_outs_up[23] ,
    \ces_1_6_io_outs_up[22] ,
    \ces_1_6_io_outs_up[21] ,
    \ces_1_6_io_outs_up[20] ,
    \ces_1_6_io_outs_up[19] ,
    \ces_1_6_io_outs_up[18] ,
    \ces_1_6_io_outs_up[17] ,
    \ces_1_6_io_outs_up[16] ,
    \ces_1_6_io_outs_up[15] ,
    \ces_1_6_io_outs_up[14] ,
    \ces_1_6_io_outs_up[13] ,
    \ces_1_6_io_outs_up[12] ,
    \ces_1_6_io_outs_up[11] ,
    \ces_1_6_io_outs_up[10] ,
    \ces_1_6_io_outs_up[9] ,
    \ces_1_6_io_outs_up[8] ,
    \ces_1_6_io_outs_up[7] ,
    \ces_1_6_io_outs_up[6] ,
    \ces_1_6_io_outs_up[5] ,
    \ces_1_6_io_outs_up[4] ,
    \ces_1_6_io_outs_up[3] ,
    \ces_1_6_io_outs_up[2] ,
    \ces_1_6_io_outs_up[1] ,
    \ces_1_6_io_outs_up[0] }),
    .io_outs_down({\ces_1_6_io_ins_down[63] ,
    \ces_1_6_io_ins_down[62] ,
    \ces_1_6_io_ins_down[61] ,
    \ces_1_6_io_ins_down[60] ,
    \ces_1_6_io_ins_down[59] ,
    \ces_1_6_io_ins_down[58] ,
    \ces_1_6_io_ins_down[57] ,
    \ces_1_6_io_ins_down[56] ,
    \ces_1_6_io_ins_down[55] ,
    \ces_1_6_io_ins_down[54] ,
    \ces_1_6_io_ins_down[53] ,
    \ces_1_6_io_ins_down[52] ,
    \ces_1_6_io_ins_down[51] ,
    \ces_1_6_io_ins_down[50] ,
    \ces_1_6_io_ins_down[49] ,
    \ces_1_6_io_ins_down[48] ,
    \ces_1_6_io_ins_down[47] ,
    \ces_1_6_io_ins_down[46] ,
    \ces_1_6_io_ins_down[45] ,
    \ces_1_6_io_ins_down[44] ,
    \ces_1_6_io_ins_down[43] ,
    \ces_1_6_io_ins_down[42] ,
    \ces_1_6_io_ins_down[41] ,
    \ces_1_6_io_ins_down[40] ,
    \ces_1_6_io_ins_down[39] ,
    \ces_1_6_io_ins_down[38] ,
    \ces_1_6_io_ins_down[37] ,
    \ces_1_6_io_ins_down[36] ,
    \ces_1_6_io_ins_down[35] ,
    \ces_1_6_io_ins_down[34] ,
    \ces_1_6_io_ins_down[33] ,
    \ces_1_6_io_ins_down[32] ,
    \ces_1_6_io_ins_down[31] ,
    \ces_1_6_io_ins_down[30] ,
    \ces_1_6_io_ins_down[29] ,
    \ces_1_6_io_ins_down[28] ,
    \ces_1_6_io_ins_down[27] ,
    \ces_1_6_io_ins_down[26] ,
    \ces_1_6_io_ins_down[25] ,
    \ces_1_6_io_ins_down[24] ,
    \ces_1_6_io_ins_down[23] ,
    \ces_1_6_io_ins_down[22] ,
    \ces_1_6_io_ins_down[21] ,
    \ces_1_6_io_ins_down[20] ,
    \ces_1_6_io_ins_down[19] ,
    \ces_1_6_io_ins_down[18] ,
    \ces_1_6_io_ins_down[17] ,
    \ces_1_6_io_ins_down[16] ,
    \ces_1_6_io_ins_down[15] ,
    \ces_1_6_io_ins_down[14] ,
    \ces_1_6_io_ins_down[13] ,
    \ces_1_6_io_ins_down[12] ,
    \ces_1_6_io_ins_down[11] ,
    \ces_1_6_io_ins_down[10] ,
    \ces_1_6_io_ins_down[9] ,
    \ces_1_6_io_ins_down[8] ,
    \ces_1_6_io_ins_down[7] ,
    \ces_1_6_io_ins_down[6] ,
    \ces_1_6_io_ins_down[5] ,
    \ces_1_6_io_ins_down[4] ,
    \ces_1_6_io_ins_down[3] ,
    \ces_1_6_io_ins_down[2] ,
    \ces_1_6_io_ins_down[1] ,
    \ces_1_6_io_ins_down[0] }),
    .io_outs_left({\ces_2_5_io_ins_left[63] ,
    \ces_2_5_io_ins_left[62] ,
    \ces_2_5_io_ins_left[61] ,
    \ces_2_5_io_ins_left[60] ,
    \ces_2_5_io_ins_left[59] ,
    \ces_2_5_io_ins_left[58] ,
    \ces_2_5_io_ins_left[57] ,
    \ces_2_5_io_ins_left[56] ,
    \ces_2_5_io_ins_left[55] ,
    \ces_2_5_io_ins_left[54] ,
    \ces_2_5_io_ins_left[53] ,
    \ces_2_5_io_ins_left[52] ,
    \ces_2_5_io_ins_left[51] ,
    \ces_2_5_io_ins_left[50] ,
    \ces_2_5_io_ins_left[49] ,
    \ces_2_5_io_ins_left[48] ,
    \ces_2_5_io_ins_left[47] ,
    \ces_2_5_io_ins_left[46] ,
    \ces_2_5_io_ins_left[45] ,
    \ces_2_5_io_ins_left[44] ,
    \ces_2_5_io_ins_left[43] ,
    \ces_2_5_io_ins_left[42] ,
    \ces_2_5_io_ins_left[41] ,
    \ces_2_5_io_ins_left[40] ,
    \ces_2_5_io_ins_left[39] ,
    \ces_2_5_io_ins_left[38] ,
    \ces_2_5_io_ins_left[37] ,
    \ces_2_5_io_ins_left[36] ,
    \ces_2_5_io_ins_left[35] ,
    \ces_2_5_io_ins_left[34] ,
    \ces_2_5_io_ins_left[33] ,
    \ces_2_5_io_ins_left[32] ,
    \ces_2_5_io_ins_left[31] ,
    \ces_2_5_io_ins_left[30] ,
    \ces_2_5_io_ins_left[29] ,
    \ces_2_5_io_ins_left[28] ,
    \ces_2_5_io_ins_left[27] ,
    \ces_2_5_io_ins_left[26] ,
    \ces_2_5_io_ins_left[25] ,
    \ces_2_5_io_ins_left[24] ,
    \ces_2_5_io_ins_left[23] ,
    \ces_2_5_io_ins_left[22] ,
    \ces_2_5_io_ins_left[21] ,
    \ces_2_5_io_ins_left[20] ,
    \ces_2_5_io_ins_left[19] ,
    \ces_2_5_io_ins_left[18] ,
    \ces_2_5_io_ins_left[17] ,
    \ces_2_5_io_ins_left[16] ,
    \ces_2_5_io_ins_left[15] ,
    \ces_2_5_io_ins_left[14] ,
    \ces_2_5_io_ins_left[13] ,
    \ces_2_5_io_ins_left[12] ,
    \ces_2_5_io_ins_left[11] ,
    \ces_2_5_io_ins_left[10] ,
    \ces_2_5_io_ins_left[9] ,
    \ces_2_5_io_ins_left[8] ,
    \ces_2_5_io_ins_left[7] ,
    \ces_2_5_io_ins_left[6] ,
    \ces_2_5_io_ins_left[5] ,
    \ces_2_5_io_ins_left[4] ,
    \ces_2_5_io_ins_left[3] ,
    \ces_2_5_io_ins_left[2] ,
    \ces_2_5_io_ins_left[1] ,
    \ces_2_5_io_ins_left[0] }),
    .io_outs_right({\ces_2_6_io_outs_right[63] ,
    \ces_2_6_io_outs_right[62] ,
    \ces_2_6_io_outs_right[61] ,
    \ces_2_6_io_outs_right[60] ,
    \ces_2_6_io_outs_right[59] ,
    \ces_2_6_io_outs_right[58] ,
    \ces_2_6_io_outs_right[57] ,
    \ces_2_6_io_outs_right[56] ,
    \ces_2_6_io_outs_right[55] ,
    \ces_2_6_io_outs_right[54] ,
    \ces_2_6_io_outs_right[53] ,
    \ces_2_6_io_outs_right[52] ,
    \ces_2_6_io_outs_right[51] ,
    \ces_2_6_io_outs_right[50] ,
    \ces_2_6_io_outs_right[49] ,
    \ces_2_6_io_outs_right[48] ,
    \ces_2_6_io_outs_right[47] ,
    \ces_2_6_io_outs_right[46] ,
    \ces_2_6_io_outs_right[45] ,
    \ces_2_6_io_outs_right[44] ,
    \ces_2_6_io_outs_right[43] ,
    \ces_2_6_io_outs_right[42] ,
    \ces_2_6_io_outs_right[41] ,
    \ces_2_6_io_outs_right[40] ,
    \ces_2_6_io_outs_right[39] ,
    \ces_2_6_io_outs_right[38] ,
    \ces_2_6_io_outs_right[37] ,
    \ces_2_6_io_outs_right[36] ,
    \ces_2_6_io_outs_right[35] ,
    \ces_2_6_io_outs_right[34] ,
    \ces_2_6_io_outs_right[33] ,
    \ces_2_6_io_outs_right[32] ,
    \ces_2_6_io_outs_right[31] ,
    \ces_2_6_io_outs_right[30] ,
    \ces_2_6_io_outs_right[29] ,
    \ces_2_6_io_outs_right[28] ,
    \ces_2_6_io_outs_right[27] ,
    \ces_2_6_io_outs_right[26] ,
    \ces_2_6_io_outs_right[25] ,
    \ces_2_6_io_outs_right[24] ,
    \ces_2_6_io_outs_right[23] ,
    \ces_2_6_io_outs_right[22] ,
    \ces_2_6_io_outs_right[21] ,
    \ces_2_6_io_outs_right[20] ,
    \ces_2_6_io_outs_right[19] ,
    \ces_2_6_io_outs_right[18] ,
    \ces_2_6_io_outs_right[17] ,
    \ces_2_6_io_outs_right[16] ,
    \ces_2_6_io_outs_right[15] ,
    \ces_2_6_io_outs_right[14] ,
    \ces_2_6_io_outs_right[13] ,
    \ces_2_6_io_outs_right[12] ,
    \ces_2_6_io_outs_right[11] ,
    \ces_2_6_io_outs_right[10] ,
    \ces_2_6_io_outs_right[9] ,
    \ces_2_6_io_outs_right[8] ,
    \ces_2_6_io_outs_right[7] ,
    \ces_2_6_io_outs_right[6] ,
    \ces_2_6_io_outs_right[5] ,
    \ces_2_6_io_outs_right[4] ,
    \ces_2_6_io_outs_right[3] ,
    \ces_2_6_io_outs_right[2] ,
    \ces_2_6_io_outs_right[1] ,
    \ces_2_6_io_outs_right[0] }),
    .io_outs_up({\ces_2_6_io_outs_up[63] ,
    \ces_2_6_io_outs_up[62] ,
    \ces_2_6_io_outs_up[61] ,
    \ces_2_6_io_outs_up[60] ,
    \ces_2_6_io_outs_up[59] ,
    \ces_2_6_io_outs_up[58] ,
    \ces_2_6_io_outs_up[57] ,
    \ces_2_6_io_outs_up[56] ,
    \ces_2_6_io_outs_up[55] ,
    \ces_2_6_io_outs_up[54] ,
    \ces_2_6_io_outs_up[53] ,
    \ces_2_6_io_outs_up[52] ,
    \ces_2_6_io_outs_up[51] ,
    \ces_2_6_io_outs_up[50] ,
    \ces_2_6_io_outs_up[49] ,
    \ces_2_6_io_outs_up[48] ,
    \ces_2_6_io_outs_up[47] ,
    \ces_2_6_io_outs_up[46] ,
    \ces_2_6_io_outs_up[45] ,
    \ces_2_6_io_outs_up[44] ,
    \ces_2_6_io_outs_up[43] ,
    \ces_2_6_io_outs_up[42] ,
    \ces_2_6_io_outs_up[41] ,
    \ces_2_6_io_outs_up[40] ,
    \ces_2_6_io_outs_up[39] ,
    \ces_2_6_io_outs_up[38] ,
    \ces_2_6_io_outs_up[37] ,
    \ces_2_6_io_outs_up[36] ,
    \ces_2_6_io_outs_up[35] ,
    \ces_2_6_io_outs_up[34] ,
    \ces_2_6_io_outs_up[33] ,
    \ces_2_6_io_outs_up[32] ,
    \ces_2_6_io_outs_up[31] ,
    \ces_2_6_io_outs_up[30] ,
    \ces_2_6_io_outs_up[29] ,
    \ces_2_6_io_outs_up[28] ,
    \ces_2_6_io_outs_up[27] ,
    \ces_2_6_io_outs_up[26] ,
    \ces_2_6_io_outs_up[25] ,
    \ces_2_6_io_outs_up[24] ,
    \ces_2_6_io_outs_up[23] ,
    \ces_2_6_io_outs_up[22] ,
    \ces_2_6_io_outs_up[21] ,
    \ces_2_6_io_outs_up[20] ,
    \ces_2_6_io_outs_up[19] ,
    \ces_2_6_io_outs_up[18] ,
    \ces_2_6_io_outs_up[17] ,
    \ces_2_6_io_outs_up[16] ,
    \ces_2_6_io_outs_up[15] ,
    \ces_2_6_io_outs_up[14] ,
    \ces_2_6_io_outs_up[13] ,
    \ces_2_6_io_outs_up[12] ,
    \ces_2_6_io_outs_up[11] ,
    \ces_2_6_io_outs_up[10] ,
    \ces_2_6_io_outs_up[9] ,
    \ces_2_6_io_outs_up[8] ,
    \ces_2_6_io_outs_up[7] ,
    \ces_2_6_io_outs_up[6] ,
    \ces_2_6_io_outs_up[5] ,
    \ces_2_6_io_outs_up[4] ,
    \ces_2_6_io_outs_up[3] ,
    \ces_2_6_io_outs_up[2] ,
    \ces_2_6_io_outs_up[1] ,
    \ces_2_6_io_outs_up[0] }));
 Element ces_2_7 (.clock(clknet_3_3_0_clock),
    .io_lsbIns_1(ces_2_6_io_lsbOuts_1),
    .io_lsbIns_2(ces_2_6_io_lsbOuts_2),
    .io_lsbIns_3(ces_2_6_io_lsbOuts_3),
    .io_lsbIns_4(ces_2_6_io_lsbOuts_4),
    .io_lsbIns_5(ces_2_6_io_lsbOuts_5),
    .io_lsbIns_6(ces_2_6_io_lsbOuts_6),
    .io_lsbIns_7(ces_2_6_io_lsbOuts_7),
    .io_lsbOuts_0(ces_2_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_2_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_2_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_2_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_2_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_2_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_2_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_2_7_io_lsbOuts_7),
    .io_ins_down({\ces_2_7_io_ins_down[63] ,
    \ces_2_7_io_ins_down[62] ,
    \ces_2_7_io_ins_down[61] ,
    \ces_2_7_io_ins_down[60] ,
    \ces_2_7_io_ins_down[59] ,
    \ces_2_7_io_ins_down[58] ,
    \ces_2_7_io_ins_down[57] ,
    \ces_2_7_io_ins_down[56] ,
    \ces_2_7_io_ins_down[55] ,
    \ces_2_7_io_ins_down[54] ,
    \ces_2_7_io_ins_down[53] ,
    \ces_2_7_io_ins_down[52] ,
    \ces_2_7_io_ins_down[51] ,
    \ces_2_7_io_ins_down[50] ,
    \ces_2_7_io_ins_down[49] ,
    \ces_2_7_io_ins_down[48] ,
    \ces_2_7_io_ins_down[47] ,
    \ces_2_7_io_ins_down[46] ,
    \ces_2_7_io_ins_down[45] ,
    \ces_2_7_io_ins_down[44] ,
    \ces_2_7_io_ins_down[43] ,
    \ces_2_7_io_ins_down[42] ,
    \ces_2_7_io_ins_down[41] ,
    \ces_2_7_io_ins_down[40] ,
    \ces_2_7_io_ins_down[39] ,
    \ces_2_7_io_ins_down[38] ,
    \ces_2_7_io_ins_down[37] ,
    \ces_2_7_io_ins_down[36] ,
    \ces_2_7_io_ins_down[35] ,
    \ces_2_7_io_ins_down[34] ,
    \ces_2_7_io_ins_down[33] ,
    \ces_2_7_io_ins_down[32] ,
    \ces_2_7_io_ins_down[31] ,
    \ces_2_7_io_ins_down[30] ,
    \ces_2_7_io_ins_down[29] ,
    \ces_2_7_io_ins_down[28] ,
    \ces_2_7_io_ins_down[27] ,
    \ces_2_7_io_ins_down[26] ,
    \ces_2_7_io_ins_down[25] ,
    \ces_2_7_io_ins_down[24] ,
    \ces_2_7_io_ins_down[23] ,
    \ces_2_7_io_ins_down[22] ,
    \ces_2_7_io_ins_down[21] ,
    \ces_2_7_io_ins_down[20] ,
    \ces_2_7_io_ins_down[19] ,
    \ces_2_7_io_ins_down[18] ,
    \ces_2_7_io_ins_down[17] ,
    \ces_2_7_io_ins_down[16] ,
    \ces_2_7_io_ins_down[15] ,
    \ces_2_7_io_ins_down[14] ,
    \ces_2_7_io_ins_down[13] ,
    \ces_2_7_io_ins_down[12] ,
    \ces_2_7_io_ins_down[11] ,
    \ces_2_7_io_ins_down[10] ,
    \ces_2_7_io_ins_down[9] ,
    \ces_2_7_io_ins_down[8] ,
    \ces_2_7_io_ins_down[7] ,
    \ces_2_7_io_ins_down[6] ,
    \ces_2_7_io_ins_down[5] ,
    \ces_2_7_io_ins_down[4] ,
    \ces_2_7_io_ins_down[3] ,
    \ces_2_7_io_ins_down[2] ,
    \ces_2_7_io_ins_down[1] ,
    \ces_2_7_io_ins_down[0] }),
    .io_ins_left({net700,
    net699,
    net698,
    net697,
    net695,
    net694,
    net693,
    net692,
    net691,
    net690,
    net689,
    net688,
    net687,
    net686,
    net684,
    net683,
    net682,
    net681,
    net680,
    net679,
    net678,
    net677,
    net676,
    net675,
    net673,
    net672,
    net671,
    net670,
    net669,
    net668,
    net667,
    net666,
    net665,
    net664,
    net662,
    net661,
    net660,
    net659,
    net658,
    net657,
    net656,
    net655,
    net654,
    net653,
    net651,
    net650,
    net649,
    net648,
    net647,
    net646,
    net645,
    net644,
    net643,
    net642,
    net704,
    net703,
    net702,
    net701,
    net696,
    net685,
    net674,
    net663,
    net652,
    net641}),
    .io_ins_right({\ces_2_6_io_outs_right[63] ,
    \ces_2_6_io_outs_right[62] ,
    \ces_2_6_io_outs_right[61] ,
    \ces_2_6_io_outs_right[60] ,
    \ces_2_6_io_outs_right[59] ,
    \ces_2_6_io_outs_right[58] ,
    \ces_2_6_io_outs_right[57] ,
    \ces_2_6_io_outs_right[56] ,
    \ces_2_6_io_outs_right[55] ,
    \ces_2_6_io_outs_right[54] ,
    \ces_2_6_io_outs_right[53] ,
    \ces_2_6_io_outs_right[52] ,
    \ces_2_6_io_outs_right[51] ,
    \ces_2_6_io_outs_right[50] ,
    \ces_2_6_io_outs_right[49] ,
    \ces_2_6_io_outs_right[48] ,
    \ces_2_6_io_outs_right[47] ,
    \ces_2_6_io_outs_right[46] ,
    \ces_2_6_io_outs_right[45] ,
    \ces_2_6_io_outs_right[44] ,
    \ces_2_6_io_outs_right[43] ,
    \ces_2_6_io_outs_right[42] ,
    \ces_2_6_io_outs_right[41] ,
    \ces_2_6_io_outs_right[40] ,
    \ces_2_6_io_outs_right[39] ,
    \ces_2_6_io_outs_right[38] ,
    \ces_2_6_io_outs_right[37] ,
    \ces_2_6_io_outs_right[36] ,
    \ces_2_6_io_outs_right[35] ,
    \ces_2_6_io_outs_right[34] ,
    \ces_2_6_io_outs_right[33] ,
    \ces_2_6_io_outs_right[32] ,
    \ces_2_6_io_outs_right[31] ,
    \ces_2_6_io_outs_right[30] ,
    \ces_2_6_io_outs_right[29] ,
    \ces_2_6_io_outs_right[28] ,
    \ces_2_6_io_outs_right[27] ,
    \ces_2_6_io_outs_right[26] ,
    \ces_2_6_io_outs_right[25] ,
    \ces_2_6_io_outs_right[24] ,
    \ces_2_6_io_outs_right[23] ,
    \ces_2_6_io_outs_right[22] ,
    \ces_2_6_io_outs_right[21] ,
    \ces_2_6_io_outs_right[20] ,
    \ces_2_6_io_outs_right[19] ,
    \ces_2_6_io_outs_right[18] ,
    \ces_2_6_io_outs_right[17] ,
    \ces_2_6_io_outs_right[16] ,
    \ces_2_6_io_outs_right[15] ,
    \ces_2_6_io_outs_right[14] ,
    \ces_2_6_io_outs_right[13] ,
    \ces_2_6_io_outs_right[12] ,
    \ces_2_6_io_outs_right[11] ,
    \ces_2_6_io_outs_right[10] ,
    \ces_2_6_io_outs_right[9] ,
    \ces_2_6_io_outs_right[8] ,
    \ces_2_6_io_outs_right[7] ,
    \ces_2_6_io_outs_right[6] ,
    \ces_2_6_io_outs_right[5] ,
    \ces_2_6_io_outs_right[4] ,
    \ces_2_6_io_outs_right[3] ,
    \ces_2_6_io_outs_right[2] ,
    \ces_2_6_io_outs_right[1] ,
    \ces_2_6_io_outs_right[0] }),
    .io_ins_up({\ces_1_7_io_outs_up[63] ,
    \ces_1_7_io_outs_up[62] ,
    \ces_1_7_io_outs_up[61] ,
    \ces_1_7_io_outs_up[60] ,
    \ces_1_7_io_outs_up[59] ,
    \ces_1_7_io_outs_up[58] ,
    \ces_1_7_io_outs_up[57] ,
    \ces_1_7_io_outs_up[56] ,
    \ces_1_7_io_outs_up[55] ,
    \ces_1_7_io_outs_up[54] ,
    \ces_1_7_io_outs_up[53] ,
    \ces_1_7_io_outs_up[52] ,
    \ces_1_7_io_outs_up[51] ,
    \ces_1_7_io_outs_up[50] ,
    \ces_1_7_io_outs_up[49] ,
    \ces_1_7_io_outs_up[48] ,
    \ces_1_7_io_outs_up[47] ,
    \ces_1_7_io_outs_up[46] ,
    \ces_1_7_io_outs_up[45] ,
    \ces_1_7_io_outs_up[44] ,
    \ces_1_7_io_outs_up[43] ,
    \ces_1_7_io_outs_up[42] ,
    \ces_1_7_io_outs_up[41] ,
    \ces_1_7_io_outs_up[40] ,
    \ces_1_7_io_outs_up[39] ,
    \ces_1_7_io_outs_up[38] ,
    \ces_1_7_io_outs_up[37] ,
    \ces_1_7_io_outs_up[36] ,
    \ces_1_7_io_outs_up[35] ,
    \ces_1_7_io_outs_up[34] ,
    \ces_1_7_io_outs_up[33] ,
    \ces_1_7_io_outs_up[32] ,
    \ces_1_7_io_outs_up[31] ,
    \ces_1_7_io_outs_up[30] ,
    \ces_1_7_io_outs_up[29] ,
    \ces_1_7_io_outs_up[28] ,
    \ces_1_7_io_outs_up[27] ,
    \ces_1_7_io_outs_up[26] ,
    \ces_1_7_io_outs_up[25] ,
    \ces_1_7_io_outs_up[24] ,
    \ces_1_7_io_outs_up[23] ,
    \ces_1_7_io_outs_up[22] ,
    \ces_1_7_io_outs_up[21] ,
    \ces_1_7_io_outs_up[20] ,
    \ces_1_7_io_outs_up[19] ,
    \ces_1_7_io_outs_up[18] ,
    \ces_1_7_io_outs_up[17] ,
    \ces_1_7_io_outs_up[16] ,
    \ces_1_7_io_outs_up[15] ,
    \ces_1_7_io_outs_up[14] ,
    \ces_1_7_io_outs_up[13] ,
    \ces_1_7_io_outs_up[12] ,
    \ces_1_7_io_outs_up[11] ,
    \ces_1_7_io_outs_up[10] ,
    \ces_1_7_io_outs_up[9] ,
    \ces_1_7_io_outs_up[8] ,
    \ces_1_7_io_outs_up[7] ,
    \ces_1_7_io_outs_up[6] ,
    \ces_1_7_io_outs_up[5] ,
    \ces_1_7_io_outs_up[4] ,
    \ces_1_7_io_outs_up[3] ,
    \ces_1_7_io_outs_up[2] ,
    \ces_1_7_io_outs_up[1] ,
    \ces_1_7_io_outs_up[0] }),
    .io_outs_down({\ces_1_7_io_ins_down[63] ,
    \ces_1_7_io_ins_down[62] ,
    \ces_1_7_io_ins_down[61] ,
    \ces_1_7_io_ins_down[60] ,
    \ces_1_7_io_ins_down[59] ,
    \ces_1_7_io_ins_down[58] ,
    \ces_1_7_io_ins_down[57] ,
    \ces_1_7_io_ins_down[56] ,
    \ces_1_7_io_ins_down[55] ,
    \ces_1_7_io_ins_down[54] ,
    \ces_1_7_io_ins_down[53] ,
    \ces_1_7_io_ins_down[52] ,
    \ces_1_7_io_ins_down[51] ,
    \ces_1_7_io_ins_down[50] ,
    \ces_1_7_io_ins_down[49] ,
    \ces_1_7_io_ins_down[48] ,
    \ces_1_7_io_ins_down[47] ,
    \ces_1_7_io_ins_down[46] ,
    \ces_1_7_io_ins_down[45] ,
    \ces_1_7_io_ins_down[44] ,
    \ces_1_7_io_ins_down[43] ,
    \ces_1_7_io_ins_down[42] ,
    \ces_1_7_io_ins_down[41] ,
    \ces_1_7_io_ins_down[40] ,
    \ces_1_7_io_ins_down[39] ,
    \ces_1_7_io_ins_down[38] ,
    \ces_1_7_io_ins_down[37] ,
    \ces_1_7_io_ins_down[36] ,
    \ces_1_7_io_ins_down[35] ,
    \ces_1_7_io_ins_down[34] ,
    \ces_1_7_io_ins_down[33] ,
    \ces_1_7_io_ins_down[32] ,
    \ces_1_7_io_ins_down[31] ,
    \ces_1_7_io_ins_down[30] ,
    \ces_1_7_io_ins_down[29] ,
    \ces_1_7_io_ins_down[28] ,
    \ces_1_7_io_ins_down[27] ,
    \ces_1_7_io_ins_down[26] ,
    \ces_1_7_io_ins_down[25] ,
    \ces_1_7_io_ins_down[24] ,
    \ces_1_7_io_ins_down[23] ,
    \ces_1_7_io_ins_down[22] ,
    \ces_1_7_io_ins_down[21] ,
    \ces_1_7_io_ins_down[20] ,
    \ces_1_7_io_ins_down[19] ,
    \ces_1_7_io_ins_down[18] ,
    \ces_1_7_io_ins_down[17] ,
    \ces_1_7_io_ins_down[16] ,
    \ces_1_7_io_ins_down[15] ,
    \ces_1_7_io_ins_down[14] ,
    \ces_1_7_io_ins_down[13] ,
    \ces_1_7_io_ins_down[12] ,
    \ces_1_7_io_ins_down[11] ,
    \ces_1_7_io_ins_down[10] ,
    \ces_1_7_io_ins_down[9] ,
    \ces_1_7_io_ins_down[8] ,
    \ces_1_7_io_ins_down[7] ,
    \ces_1_7_io_ins_down[6] ,
    \ces_1_7_io_ins_down[5] ,
    \ces_1_7_io_ins_down[4] ,
    \ces_1_7_io_ins_down[3] ,
    \ces_1_7_io_ins_down[2] ,
    \ces_1_7_io_ins_down[1] ,
    \ces_1_7_io_ins_down[0] }),
    .io_outs_left({\ces_2_6_io_ins_left[63] ,
    \ces_2_6_io_ins_left[62] ,
    \ces_2_6_io_ins_left[61] ,
    \ces_2_6_io_ins_left[60] ,
    \ces_2_6_io_ins_left[59] ,
    \ces_2_6_io_ins_left[58] ,
    \ces_2_6_io_ins_left[57] ,
    \ces_2_6_io_ins_left[56] ,
    \ces_2_6_io_ins_left[55] ,
    \ces_2_6_io_ins_left[54] ,
    \ces_2_6_io_ins_left[53] ,
    \ces_2_6_io_ins_left[52] ,
    \ces_2_6_io_ins_left[51] ,
    \ces_2_6_io_ins_left[50] ,
    \ces_2_6_io_ins_left[49] ,
    \ces_2_6_io_ins_left[48] ,
    \ces_2_6_io_ins_left[47] ,
    \ces_2_6_io_ins_left[46] ,
    \ces_2_6_io_ins_left[45] ,
    \ces_2_6_io_ins_left[44] ,
    \ces_2_6_io_ins_left[43] ,
    \ces_2_6_io_ins_left[42] ,
    \ces_2_6_io_ins_left[41] ,
    \ces_2_6_io_ins_left[40] ,
    \ces_2_6_io_ins_left[39] ,
    \ces_2_6_io_ins_left[38] ,
    \ces_2_6_io_ins_left[37] ,
    \ces_2_6_io_ins_left[36] ,
    \ces_2_6_io_ins_left[35] ,
    \ces_2_6_io_ins_left[34] ,
    \ces_2_6_io_ins_left[33] ,
    \ces_2_6_io_ins_left[32] ,
    \ces_2_6_io_ins_left[31] ,
    \ces_2_6_io_ins_left[30] ,
    \ces_2_6_io_ins_left[29] ,
    \ces_2_6_io_ins_left[28] ,
    \ces_2_6_io_ins_left[27] ,
    \ces_2_6_io_ins_left[26] ,
    \ces_2_6_io_ins_left[25] ,
    \ces_2_6_io_ins_left[24] ,
    \ces_2_6_io_ins_left[23] ,
    \ces_2_6_io_ins_left[22] ,
    \ces_2_6_io_ins_left[21] ,
    \ces_2_6_io_ins_left[20] ,
    \ces_2_6_io_ins_left[19] ,
    \ces_2_6_io_ins_left[18] ,
    \ces_2_6_io_ins_left[17] ,
    \ces_2_6_io_ins_left[16] ,
    \ces_2_6_io_ins_left[15] ,
    \ces_2_6_io_ins_left[14] ,
    \ces_2_6_io_ins_left[13] ,
    \ces_2_6_io_ins_left[12] ,
    \ces_2_6_io_ins_left[11] ,
    \ces_2_6_io_ins_left[10] ,
    \ces_2_6_io_ins_left[9] ,
    \ces_2_6_io_ins_left[8] ,
    \ces_2_6_io_ins_left[7] ,
    \ces_2_6_io_ins_left[6] ,
    \ces_2_6_io_ins_left[5] ,
    \ces_2_6_io_ins_left[4] ,
    \ces_2_6_io_ins_left[3] ,
    \ces_2_6_io_ins_left[2] ,
    \ces_2_6_io_ins_left[1] ,
    \ces_2_6_io_ins_left[0] }),
    .io_outs_right({net3324,
    net3323,
    net3322,
    net3321,
    net3319,
    net3318,
    net3317,
    net3316,
    net3315,
    net3314,
    net3313,
    net3312,
    net3311,
    net3310,
    net3308,
    net3307,
    net3306,
    net3305,
    net3304,
    net3303,
    net3302,
    net3301,
    net3300,
    net3299,
    net3297,
    net3296,
    net3295,
    net3294,
    net3293,
    net3292,
    net3291,
    net3290,
    net3289,
    net3288,
    net3286,
    net3285,
    net3284,
    net3283,
    net3282,
    net3281,
    net3280,
    net3279,
    net3278,
    net3277,
    net3275,
    net3274,
    net3273,
    net3272,
    net3271,
    net3270,
    net3269,
    net3268,
    net3267,
    net3266,
    net3328,
    net3327,
    net3326,
    net3325,
    net3320,
    net3309,
    net3298,
    net3287,
    net3276,
    net3265}),
    .io_outs_up({\ces_2_7_io_outs_up[63] ,
    \ces_2_7_io_outs_up[62] ,
    \ces_2_7_io_outs_up[61] ,
    \ces_2_7_io_outs_up[60] ,
    \ces_2_7_io_outs_up[59] ,
    \ces_2_7_io_outs_up[58] ,
    \ces_2_7_io_outs_up[57] ,
    \ces_2_7_io_outs_up[56] ,
    \ces_2_7_io_outs_up[55] ,
    \ces_2_7_io_outs_up[54] ,
    \ces_2_7_io_outs_up[53] ,
    \ces_2_7_io_outs_up[52] ,
    \ces_2_7_io_outs_up[51] ,
    \ces_2_7_io_outs_up[50] ,
    \ces_2_7_io_outs_up[49] ,
    \ces_2_7_io_outs_up[48] ,
    \ces_2_7_io_outs_up[47] ,
    \ces_2_7_io_outs_up[46] ,
    \ces_2_7_io_outs_up[45] ,
    \ces_2_7_io_outs_up[44] ,
    \ces_2_7_io_outs_up[43] ,
    \ces_2_7_io_outs_up[42] ,
    \ces_2_7_io_outs_up[41] ,
    \ces_2_7_io_outs_up[40] ,
    \ces_2_7_io_outs_up[39] ,
    \ces_2_7_io_outs_up[38] ,
    \ces_2_7_io_outs_up[37] ,
    \ces_2_7_io_outs_up[36] ,
    \ces_2_7_io_outs_up[35] ,
    \ces_2_7_io_outs_up[34] ,
    \ces_2_7_io_outs_up[33] ,
    \ces_2_7_io_outs_up[32] ,
    \ces_2_7_io_outs_up[31] ,
    \ces_2_7_io_outs_up[30] ,
    \ces_2_7_io_outs_up[29] ,
    \ces_2_7_io_outs_up[28] ,
    \ces_2_7_io_outs_up[27] ,
    \ces_2_7_io_outs_up[26] ,
    \ces_2_7_io_outs_up[25] ,
    \ces_2_7_io_outs_up[24] ,
    \ces_2_7_io_outs_up[23] ,
    \ces_2_7_io_outs_up[22] ,
    \ces_2_7_io_outs_up[21] ,
    \ces_2_7_io_outs_up[20] ,
    \ces_2_7_io_outs_up[19] ,
    \ces_2_7_io_outs_up[18] ,
    \ces_2_7_io_outs_up[17] ,
    \ces_2_7_io_outs_up[16] ,
    \ces_2_7_io_outs_up[15] ,
    \ces_2_7_io_outs_up[14] ,
    \ces_2_7_io_outs_up[13] ,
    \ces_2_7_io_outs_up[12] ,
    \ces_2_7_io_outs_up[11] ,
    \ces_2_7_io_outs_up[10] ,
    \ces_2_7_io_outs_up[9] ,
    \ces_2_7_io_outs_up[8] ,
    \ces_2_7_io_outs_up[7] ,
    \ces_2_7_io_outs_up[6] ,
    \ces_2_7_io_outs_up[5] ,
    \ces_2_7_io_outs_up[4] ,
    \ces_2_7_io_outs_up[3] ,
    \ces_2_7_io_outs_up[2] ,
    \ces_2_7_io_outs_up[1] ,
    \ces_2_7_io_outs_up[0] }));
 Element ces_3_0 (.clock(clknet_3_1_0_clock),
    .io_lsbIns_1(net4182),
    .io_lsbIns_2(net4183),
    .io_lsbIns_3(net4184),
    .io_lsbIns_4(net4185),
    .io_lsbIns_5(net4186),
    .io_lsbIns_6(net4187),
    .io_lsbIns_7(net4188),
    .io_lsbOuts_0(ces_3_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_0_io_lsbOuts_7),
    .io_ins_down({\ces_3_0_io_ins_down[63] ,
    \ces_3_0_io_ins_down[62] ,
    \ces_3_0_io_ins_down[61] ,
    \ces_3_0_io_ins_down[60] ,
    \ces_3_0_io_ins_down[59] ,
    \ces_3_0_io_ins_down[58] ,
    \ces_3_0_io_ins_down[57] ,
    \ces_3_0_io_ins_down[56] ,
    \ces_3_0_io_ins_down[55] ,
    \ces_3_0_io_ins_down[54] ,
    \ces_3_0_io_ins_down[53] ,
    \ces_3_0_io_ins_down[52] ,
    \ces_3_0_io_ins_down[51] ,
    \ces_3_0_io_ins_down[50] ,
    \ces_3_0_io_ins_down[49] ,
    \ces_3_0_io_ins_down[48] ,
    \ces_3_0_io_ins_down[47] ,
    \ces_3_0_io_ins_down[46] ,
    \ces_3_0_io_ins_down[45] ,
    \ces_3_0_io_ins_down[44] ,
    \ces_3_0_io_ins_down[43] ,
    \ces_3_0_io_ins_down[42] ,
    \ces_3_0_io_ins_down[41] ,
    \ces_3_0_io_ins_down[40] ,
    \ces_3_0_io_ins_down[39] ,
    \ces_3_0_io_ins_down[38] ,
    \ces_3_0_io_ins_down[37] ,
    \ces_3_0_io_ins_down[36] ,
    \ces_3_0_io_ins_down[35] ,
    \ces_3_0_io_ins_down[34] ,
    \ces_3_0_io_ins_down[33] ,
    \ces_3_0_io_ins_down[32] ,
    \ces_3_0_io_ins_down[31] ,
    \ces_3_0_io_ins_down[30] ,
    \ces_3_0_io_ins_down[29] ,
    \ces_3_0_io_ins_down[28] ,
    \ces_3_0_io_ins_down[27] ,
    \ces_3_0_io_ins_down[26] ,
    \ces_3_0_io_ins_down[25] ,
    \ces_3_0_io_ins_down[24] ,
    \ces_3_0_io_ins_down[23] ,
    \ces_3_0_io_ins_down[22] ,
    \ces_3_0_io_ins_down[21] ,
    \ces_3_0_io_ins_down[20] ,
    \ces_3_0_io_ins_down[19] ,
    \ces_3_0_io_ins_down[18] ,
    \ces_3_0_io_ins_down[17] ,
    \ces_3_0_io_ins_down[16] ,
    \ces_3_0_io_ins_down[15] ,
    \ces_3_0_io_ins_down[14] ,
    \ces_3_0_io_ins_down[13] ,
    \ces_3_0_io_ins_down[12] ,
    \ces_3_0_io_ins_down[11] ,
    \ces_3_0_io_ins_down[10] ,
    \ces_3_0_io_ins_down[9] ,
    \ces_3_0_io_ins_down[8] ,
    \ces_3_0_io_ins_down[7] ,
    \ces_3_0_io_ins_down[6] ,
    \ces_3_0_io_ins_down[5] ,
    \ces_3_0_io_ins_down[4] ,
    \ces_3_0_io_ins_down[3] ,
    \ces_3_0_io_ins_down[2] ,
    \ces_3_0_io_ins_down[1] ,
    \ces_3_0_io_ins_down[0] }),
    .io_ins_left({\ces_3_0_io_ins_left[63] ,
    \ces_3_0_io_ins_left[62] ,
    \ces_3_0_io_ins_left[61] ,
    \ces_3_0_io_ins_left[60] ,
    \ces_3_0_io_ins_left[59] ,
    \ces_3_0_io_ins_left[58] ,
    \ces_3_0_io_ins_left[57] ,
    \ces_3_0_io_ins_left[56] ,
    \ces_3_0_io_ins_left[55] ,
    \ces_3_0_io_ins_left[54] ,
    \ces_3_0_io_ins_left[53] ,
    \ces_3_0_io_ins_left[52] ,
    \ces_3_0_io_ins_left[51] ,
    \ces_3_0_io_ins_left[50] ,
    \ces_3_0_io_ins_left[49] ,
    \ces_3_0_io_ins_left[48] ,
    \ces_3_0_io_ins_left[47] ,
    \ces_3_0_io_ins_left[46] ,
    \ces_3_0_io_ins_left[45] ,
    \ces_3_0_io_ins_left[44] ,
    \ces_3_0_io_ins_left[43] ,
    \ces_3_0_io_ins_left[42] ,
    \ces_3_0_io_ins_left[41] ,
    \ces_3_0_io_ins_left[40] ,
    \ces_3_0_io_ins_left[39] ,
    \ces_3_0_io_ins_left[38] ,
    \ces_3_0_io_ins_left[37] ,
    \ces_3_0_io_ins_left[36] ,
    \ces_3_0_io_ins_left[35] ,
    \ces_3_0_io_ins_left[34] ,
    \ces_3_0_io_ins_left[33] ,
    \ces_3_0_io_ins_left[32] ,
    \ces_3_0_io_ins_left[31] ,
    \ces_3_0_io_ins_left[30] ,
    \ces_3_0_io_ins_left[29] ,
    \ces_3_0_io_ins_left[28] ,
    \ces_3_0_io_ins_left[27] ,
    \ces_3_0_io_ins_left[26] ,
    \ces_3_0_io_ins_left[25] ,
    \ces_3_0_io_ins_left[24] ,
    \ces_3_0_io_ins_left[23] ,
    \ces_3_0_io_ins_left[22] ,
    \ces_3_0_io_ins_left[21] ,
    \ces_3_0_io_ins_left[20] ,
    \ces_3_0_io_ins_left[19] ,
    \ces_3_0_io_ins_left[18] ,
    \ces_3_0_io_ins_left[17] ,
    \ces_3_0_io_ins_left[16] ,
    \ces_3_0_io_ins_left[15] ,
    \ces_3_0_io_ins_left[14] ,
    \ces_3_0_io_ins_left[13] ,
    \ces_3_0_io_ins_left[12] ,
    \ces_3_0_io_ins_left[11] ,
    \ces_3_0_io_ins_left[10] ,
    \ces_3_0_io_ins_left[9] ,
    \ces_3_0_io_ins_left[8] ,
    \ces_3_0_io_ins_left[7] ,
    \ces_3_0_io_ins_left[6] ,
    \ces_3_0_io_ins_left[5] ,
    \ces_3_0_io_ins_left[4] ,
    \ces_3_0_io_ins_left[3] ,
    \ces_3_0_io_ins_left[2] ,
    \ces_3_0_io_ins_left[1] ,
    \ces_3_0_io_ins_left[0] }),
    .io_ins_right({net1276,
    net1275,
    net1274,
    net1273,
    net1271,
    net1270,
    net1269,
    net1268,
    net1267,
    net1266,
    net1265,
    net1264,
    net1263,
    net1262,
    net1260,
    net1259,
    net1258,
    net1257,
    net1256,
    net1255,
    net1254,
    net1253,
    net1252,
    net1251,
    net1249,
    net1248,
    net1247,
    net1246,
    net1245,
    net1244,
    net1243,
    net1242,
    net1241,
    net1240,
    net1238,
    net1237,
    net1236,
    net1235,
    net1234,
    net1233,
    net1232,
    net1231,
    net1230,
    net1229,
    net1227,
    net1226,
    net1225,
    net1224,
    net1223,
    net1222,
    net1221,
    net1220,
    net1219,
    net1218,
    net1280,
    net1279,
    net1278,
    net1277,
    net1272,
    net1261,
    net1250,
    net1239,
    net1228,
    net1217}),
    .io_ins_up({\ces_2_0_io_outs_up[63] ,
    \ces_2_0_io_outs_up[62] ,
    \ces_2_0_io_outs_up[61] ,
    \ces_2_0_io_outs_up[60] ,
    \ces_2_0_io_outs_up[59] ,
    \ces_2_0_io_outs_up[58] ,
    \ces_2_0_io_outs_up[57] ,
    \ces_2_0_io_outs_up[56] ,
    \ces_2_0_io_outs_up[55] ,
    \ces_2_0_io_outs_up[54] ,
    \ces_2_0_io_outs_up[53] ,
    \ces_2_0_io_outs_up[52] ,
    \ces_2_0_io_outs_up[51] ,
    \ces_2_0_io_outs_up[50] ,
    \ces_2_0_io_outs_up[49] ,
    \ces_2_0_io_outs_up[48] ,
    \ces_2_0_io_outs_up[47] ,
    \ces_2_0_io_outs_up[46] ,
    \ces_2_0_io_outs_up[45] ,
    \ces_2_0_io_outs_up[44] ,
    \ces_2_0_io_outs_up[43] ,
    \ces_2_0_io_outs_up[42] ,
    \ces_2_0_io_outs_up[41] ,
    \ces_2_0_io_outs_up[40] ,
    \ces_2_0_io_outs_up[39] ,
    \ces_2_0_io_outs_up[38] ,
    \ces_2_0_io_outs_up[37] ,
    \ces_2_0_io_outs_up[36] ,
    \ces_2_0_io_outs_up[35] ,
    \ces_2_0_io_outs_up[34] ,
    \ces_2_0_io_outs_up[33] ,
    \ces_2_0_io_outs_up[32] ,
    \ces_2_0_io_outs_up[31] ,
    \ces_2_0_io_outs_up[30] ,
    \ces_2_0_io_outs_up[29] ,
    \ces_2_0_io_outs_up[28] ,
    \ces_2_0_io_outs_up[27] ,
    \ces_2_0_io_outs_up[26] ,
    \ces_2_0_io_outs_up[25] ,
    \ces_2_0_io_outs_up[24] ,
    \ces_2_0_io_outs_up[23] ,
    \ces_2_0_io_outs_up[22] ,
    \ces_2_0_io_outs_up[21] ,
    \ces_2_0_io_outs_up[20] ,
    \ces_2_0_io_outs_up[19] ,
    \ces_2_0_io_outs_up[18] ,
    \ces_2_0_io_outs_up[17] ,
    \ces_2_0_io_outs_up[16] ,
    \ces_2_0_io_outs_up[15] ,
    \ces_2_0_io_outs_up[14] ,
    \ces_2_0_io_outs_up[13] ,
    \ces_2_0_io_outs_up[12] ,
    \ces_2_0_io_outs_up[11] ,
    \ces_2_0_io_outs_up[10] ,
    \ces_2_0_io_outs_up[9] ,
    \ces_2_0_io_outs_up[8] ,
    \ces_2_0_io_outs_up[7] ,
    \ces_2_0_io_outs_up[6] ,
    \ces_2_0_io_outs_up[5] ,
    \ces_2_0_io_outs_up[4] ,
    \ces_2_0_io_outs_up[3] ,
    \ces_2_0_io_outs_up[2] ,
    \ces_2_0_io_outs_up[1] ,
    \ces_2_0_io_outs_up[0] }),
    .io_outs_down({\ces_2_0_io_ins_down[63] ,
    \ces_2_0_io_ins_down[62] ,
    \ces_2_0_io_ins_down[61] ,
    \ces_2_0_io_ins_down[60] ,
    \ces_2_0_io_ins_down[59] ,
    \ces_2_0_io_ins_down[58] ,
    \ces_2_0_io_ins_down[57] ,
    \ces_2_0_io_ins_down[56] ,
    \ces_2_0_io_ins_down[55] ,
    \ces_2_0_io_ins_down[54] ,
    \ces_2_0_io_ins_down[53] ,
    \ces_2_0_io_ins_down[52] ,
    \ces_2_0_io_ins_down[51] ,
    \ces_2_0_io_ins_down[50] ,
    \ces_2_0_io_ins_down[49] ,
    \ces_2_0_io_ins_down[48] ,
    \ces_2_0_io_ins_down[47] ,
    \ces_2_0_io_ins_down[46] ,
    \ces_2_0_io_ins_down[45] ,
    \ces_2_0_io_ins_down[44] ,
    \ces_2_0_io_ins_down[43] ,
    \ces_2_0_io_ins_down[42] ,
    \ces_2_0_io_ins_down[41] ,
    \ces_2_0_io_ins_down[40] ,
    \ces_2_0_io_ins_down[39] ,
    \ces_2_0_io_ins_down[38] ,
    \ces_2_0_io_ins_down[37] ,
    \ces_2_0_io_ins_down[36] ,
    \ces_2_0_io_ins_down[35] ,
    \ces_2_0_io_ins_down[34] ,
    \ces_2_0_io_ins_down[33] ,
    \ces_2_0_io_ins_down[32] ,
    \ces_2_0_io_ins_down[31] ,
    \ces_2_0_io_ins_down[30] ,
    \ces_2_0_io_ins_down[29] ,
    \ces_2_0_io_ins_down[28] ,
    \ces_2_0_io_ins_down[27] ,
    \ces_2_0_io_ins_down[26] ,
    \ces_2_0_io_ins_down[25] ,
    \ces_2_0_io_ins_down[24] ,
    \ces_2_0_io_ins_down[23] ,
    \ces_2_0_io_ins_down[22] ,
    \ces_2_0_io_ins_down[21] ,
    \ces_2_0_io_ins_down[20] ,
    \ces_2_0_io_ins_down[19] ,
    \ces_2_0_io_ins_down[18] ,
    \ces_2_0_io_ins_down[17] ,
    \ces_2_0_io_ins_down[16] ,
    \ces_2_0_io_ins_down[15] ,
    \ces_2_0_io_ins_down[14] ,
    \ces_2_0_io_ins_down[13] ,
    \ces_2_0_io_ins_down[12] ,
    \ces_2_0_io_ins_down[11] ,
    \ces_2_0_io_ins_down[10] ,
    \ces_2_0_io_ins_down[9] ,
    \ces_2_0_io_ins_down[8] ,
    \ces_2_0_io_ins_down[7] ,
    \ces_2_0_io_ins_down[6] ,
    \ces_2_0_io_ins_down[5] ,
    \ces_2_0_io_ins_down[4] ,
    \ces_2_0_io_ins_down[3] ,
    \ces_2_0_io_ins_down[2] ,
    \ces_2_0_io_ins_down[1] ,
    \ces_2_0_io_ins_down[0] }),
    .io_outs_left({net2876,
    net2875,
    net2874,
    net2873,
    net2871,
    net2870,
    net2869,
    net2868,
    net2867,
    net2866,
    net2865,
    net2864,
    net2863,
    net2862,
    net2860,
    net2859,
    net2858,
    net2857,
    net2856,
    net2855,
    net2854,
    net2853,
    net2852,
    net2851,
    net2849,
    net2848,
    net2847,
    net2846,
    net2845,
    net2844,
    net2843,
    net2842,
    net2841,
    net2840,
    net2838,
    net2837,
    net2836,
    net2835,
    net2834,
    net2833,
    net2832,
    net2831,
    net2830,
    net2829,
    net2827,
    net2826,
    net2825,
    net2824,
    net2823,
    net2822,
    net2821,
    net2820,
    net2819,
    net2818,
    net2880,
    net2879,
    net2878,
    net2877,
    net2872,
    net2861,
    net2850,
    net2839,
    net2828,
    net2817}),
    .io_outs_right({\ces_3_0_io_outs_right[63] ,
    \ces_3_0_io_outs_right[62] ,
    \ces_3_0_io_outs_right[61] ,
    \ces_3_0_io_outs_right[60] ,
    \ces_3_0_io_outs_right[59] ,
    \ces_3_0_io_outs_right[58] ,
    \ces_3_0_io_outs_right[57] ,
    \ces_3_0_io_outs_right[56] ,
    \ces_3_0_io_outs_right[55] ,
    \ces_3_0_io_outs_right[54] ,
    \ces_3_0_io_outs_right[53] ,
    \ces_3_0_io_outs_right[52] ,
    \ces_3_0_io_outs_right[51] ,
    \ces_3_0_io_outs_right[50] ,
    \ces_3_0_io_outs_right[49] ,
    \ces_3_0_io_outs_right[48] ,
    \ces_3_0_io_outs_right[47] ,
    \ces_3_0_io_outs_right[46] ,
    \ces_3_0_io_outs_right[45] ,
    \ces_3_0_io_outs_right[44] ,
    \ces_3_0_io_outs_right[43] ,
    \ces_3_0_io_outs_right[42] ,
    \ces_3_0_io_outs_right[41] ,
    \ces_3_0_io_outs_right[40] ,
    \ces_3_0_io_outs_right[39] ,
    \ces_3_0_io_outs_right[38] ,
    \ces_3_0_io_outs_right[37] ,
    \ces_3_0_io_outs_right[36] ,
    \ces_3_0_io_outs_right[35] ,
    \ces_3_0_io_outs_right[34] ,
    \ces_3_0_io_outs_right[33] ,
    \ces_3_0_io_outs_right[32] ,
    \ces_3_0_io_outs_right[31] ,
    \ces_3_0_io_outs_right[30] ,
    \ces_3_0_io_outs_right[29] ,
    \ces_3_0_io_outs_right[28] ,
    \ces_3_0_io_outs_right[27] ,
    \ces_3_0_io_outs_right[26] ,
    \ces_3_0_io_outs_right[25] ,
    \ces_3_0_io_outs_right[24] ,
    \ces_3_0_io_outs_right[23] ,
    \ces_3_0_io_outs_right[22] ,
    \ces_3_0_io_outs_right[21] ,
    \ces_3_0_io_outs_right[20] ,
    \ces_3_0_io_outs_right[19] ,
    \ces_3_0_io_outs_right[18] ,
    \ces_3_0_io_outs_right[17] ,
    \ces_3_0_io_outs_right[16] ,
    \ces_3_0_io_outs_right[15] ,
    \ces_3_0_io_outs_right[14] ,
    \ces_3_0_io_outs_right[13] ,
    \ces_3_0_io_outs_right[12] ,
    \ces_3_0_io_outs_right[11] ,
    \ces_3_0_io_outs_right[10] ,
    \ces_3_0_io_outs_right[9] ,
    \ces_3_0_io_outs_right[8] ,
    \ces_3_0_io_outs_right[7] ,
    \ces_3_0_io_outs_right[6] ,
    \ces_3_0_io_outs_right[5] ,
    \ces_3_0_io_outs_right[4] ,
    \ces_3_0_io_outs_right[3] ,
    \ces_3_0_io_outs_right[2] ,
    \ces_3_0_io_outs_right[1] ,
    \ces_3_0_io_outs_right[0] }),
    .io_outs_up({\ces_3_0_io_outs_up[63] ,
    \ces_3_0_io_outs_up[62] ,
    \ces_3_0_io_outs_up[61] ,
    \ces_3_0_io_outs_up[60] ,
    \ces_3_0_io_outs_up[59] ,
    \ces_3_0_io_outs_up[58] ,
    \ces_3_0_io_outs_up[57] ,
    \ces_3_0_io_outs_up[56] ,
    \ces_3_0_io_outs_up[55] ,
    \ces_3_0_io_outs_up[54] ,
    \ces_3_0_io_outs_up[53] ,
    \ces_3_0_io_outs_up[52] ,
    \ces_3_0_io_outs_up[51] ,
    \ces_3_0_io_outs_up[50] ,
    \ces_3_0_io_outs_up[49] ,
    \ces_3_0_io_outs_up[48] ,
    \ces_3_0_io_outs_up[47] ,
    \ces_3_0_io_outs_up[46] ,
    \ces_3_0_io_outs_up[45] ,
    \ces_3_0_io_outs_up[44] ,
    \ces_3_0_io_outs_up[43] ,
    \ces_3_0_io_outs_up[42] ,
    \ces_3_0_io_outs_up[41] ,
    \ces_3_0_io_outs_up[40] ,
    \ces_3_0_io_outs_up[39] ,
    \ces_3_0_io_outs_up[38] ,
    \ces_3_0_io_outs_up[37] ,
    \ces_3_0_io_outs_up[36] ,
    \ces_3_0_io_outs_up[35] ,
    \ces_3_0_io_outs_up[34] ,
    \ces_3_0_io_outs_up[33] ,
    \ces_3_0_io_outs_up[32] ,
    \ces_3_0_io_outs_up[31] ,
    \ces_3_0_io_outs_up[30] ,
    \ces_3_0_io_outs_up[29] ,
    \ces_3_0_io_outs_up[28] ,
    \ces_3_0_io_outs_up[27] ,
    \ces_3_0_io_outs_up[26] ,
    \ces_3_0_io_outs_up[25] ,
    \ces_3_0_io_outs_up[24] ,
    \ces_3_0_io_outs_up[23] ,
    \ces_3_0_io_outs_up[22] ,
    \ces_3_0_io_outs_up[21] ,
    \ces_3_0_io_outs_up[20] ,
    \ces_3_0_io_outs_up[19] ,
    \ces_3_0_io_outs_up[18] ,
    \ces_3_0_io_outs_up[17] ,
    \ces_3_0_io_outs_up[16] ,
    \ces_3_0_io_outs_up[15] ,
    \ces_3_0_io_outs_up[14] ,
    \ces_3_0_io_outs_up[13] ,
    \ces_3_0_io_outs_up[12] ,
    \ces_3_0_io_outs_up[11] ,
    \ces_3_0_io_outs_up[10] ,
    \ces_3_0_io_outs_up[9] ,
    \ces_3_0_io_outs_up[8] ,
    \ces_3_0_io_outs_up[7] ,
    \ces_3_0_io_outs_up[6] ,
    \ces_3_0_io_outs_up[5] ,
    \ces_3_0_io_outs_up[4] ,
    \ces_3_0_io_outs_up[3] ,
    \ces_3_0_io_outs_up[2] ,
    \ces_3_0_io_outs_up[1] ,
    \ces_3_0_io_outs_up[0] }));
 Element ces_3_1 (.clock(clknet_3_1_0_clock),
    .io_lsbIns_1(ces_3_0_io_lsbOuts_1),
    .io_lsbIns_2(ces_3_0_io_lsbOuts_2),
    .io_lsbIns_3(ces_3_0_io_lsbOuts_3),
    .io_lsbIns_4(ces_3_0_io_lsbOuts_4),
    .io_lsbIns_5(ces_3_0_io_lsbOuts_5),
    .io_lsbIns_6(ces_3_0_io_lsbOuts_6),
    .io_lsbIns_7(ces_3_0_io_lsbOuts_7),
    .io_lsbOuts_0(ces_3_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_1_io_lsbOuts_7),
    .io_ins_down({\ces_3_1_io_ins_down[63] ,
    \ces_3_1_io_ins_down[62] ,
    \ces_3_1_io_ins_down[61] ,
    \ces_3_1_io_ins_down[60] ,
    \ces_3_1_io_ins_down[59] ,
    \ces_3_1_io_ins_down[58] ,
    \ces_3_1_io_ins_down[57] ,
    \ces_3_1_io_ins_down[56] ,
    \ces_3_1_io_ins_down[55] ,
    \ces_3_1_io_ins_down[54] ,
    \ces_3_1_io_ins_down[53] ,
    \ces_3_1_io_ins_down[52] ,
    \ces_3_1_io_ins_down[51] ,
    \ces_3_1_io_ins_down[50] ,
    \ces_3_1_io_ins_down[49] ,
    \ces_3_1_io_ins_down[48] ,
    \ces_3_1_io_ins_down[47] ,
    \ces_3_1_io_ins_down[46] ,
    \ces_3_1_io_ins_down[45] ,
    \ces_3_1_io_ins_down[44] ,
    \ces_3_1_io_ins_down[43] ,
    \ces_3_1_io_ins_down[42] ,
    \ces_3_1_io_ins_down[41] ,
    \ces_3_1_io_ins_down[40] ,
    \ces_3_1_io_ins_down[39] ,
    \ces_3_1_io_ins_down[38] ,
    \ces_3_1_io_ins_down[37] ,
    \ces_3_1_io_ins_down[36] ,
    \ces_3_1_io_ins_down[35] ,
    \ces_3_1_io_ins_down[34] ,
    \ces_3_1_io_ins_down[33] ,
    \ces_3_1_io_ins_down[32] ,
    \ces_3_1_io_ins_down[31] ,
    \ces_3_1_io_ins_down[30] ,
    \ces_3_1_io_ins_down[29] ,
    \ces_3_1_io_ins_down[28] ,
    \ces_3_1_io_ins_down[27] ,
    \ces_3_1_io_ins_down[26] ,
    \ces_3_1_io_ins_down[25] ,
    \ces_3_1_io_ins_down[24] ,
    \ces_3_1_io_ins_down[23] ,
    \ces_3_1_io_ins_down[22] ,
    \ces_3_1_io_ins_down[21] ,
    \ces_3_1_io_ins_down[20] ,
    \ces_3_1_io_ins_down[19] ,
    \ces_3_1_io_ins_down[18] ,
    \ces_3_1_io_ins_down[17] ,
    \ces_3_1_io_ins_down[16] ,
    \ces_3_1_io_ins_down[15] ,
    \ces_3_1_io_ins_down[14] ,
    \ces_3_1_io_ins_down[13] ,
    \ces_3_1_io_ins_down[12] ,
    \ces_3_1_io_ins_down[11] ,
    \ces_3_1_io_ins_down[10] ,
    \ces_3_1_io_ins_down[9] ,
    \ces_3_1_io_ins_down[8] ,
    \ces_3_1_io_ins_down[7] ,
    \ces_3_1_io_ins_down[6] ,
    \ces_3_1_io_ins_down[5] ,
    \ces_3_1_io_ins_down[4] ,
    \ces_3_1_io_ins_down[3] ,
    \ces_3_1_io_ins_down[2] ,
    \ces_3_1_io_ins_down[1] ,
    \ces_3_1_io_ins_down[0] }),
    .io_ins_left({\ces_3_1_io_ins_left[63] ,
    \ces_3_1_io_ins_left[62] ,
    \ces_3_1_io_ins_left[61] ,
    \ces_3_1_io_ins_left[60] ,
    \ces_3_1_io_ins_left[59] ,
    \ces_3_1_io_ins_left[58] ,
    \ces_3_1_io_ins_left[57] ,
    \ces_3_1_io_ins_left[56] ,
    \ces_3_1_io_ins_left[55] ,
    \ces_3_1_io_ins_left[54] ,
    \ces_3_1_io_ins_left[53] ,
    \ces_3_1_io_ins_left[52] ,
    \ces_3_1_io_ins_left[51] ,
    \ces_3_1_io_ins_left[50] ,
    \ces_3_1_io_ins_left[49] ,
    \ces_3_1_io_ins_left[48] ,
    \ces_3_1_io_ins_left[47] ,
    \ces_3_1_io_ins_left[46] ,
    \ces_3_1_io_ins_left[45] ,
    \ces_3_1_io_ins_left[44] ,
    \ces_3_1_io_ins_left[43] ,
    \ces_3_1_io_ins_left[42] ,
    \ces_3_1_io_ins_left[41] ,
    \ces_3_1_io_ins_left[40] ,
    \ces_3_1_io_ins_left[39] ,
    \ces_3_1_io_ins_left[38] ,
    \ces_3_1_io_ins_left[37] ,
    \ces_3_1_io_ins_left[36] ,
    \ces_3_1_io_ins_left[35] ,
    \ces_3_1_io_ins_left[34] ,
    \ces_3_1_io_ins_left[33] ,
    \ces_3_1_io_ins_left[32] ,
    \ces_3_1_io_ins_left[31] ,
    \ces_3_1_io_ins_left[30] ,
    \ces_3_1_io_ins_left[29] ,
    \ces_3_1_io_ins_left[28] ,
    \ces_3_1_io_ins_left[27] ,
    \ces_3_1_io_ins_left[26] ,
    \ces_3_1_io_ins_left[25] ,
    \ces_3_1_io_ins_left[24] ,
    \ces_3_1_io_ins_left[23] ,
    \ces_3_1_io_ins_left[22] ,
    \ces_3_1_io_ins_left[21] ,
    \ces_3_1_io_ins_left[20] ,
    \ces_3_1_io_ins_left[19] ,
    \ces_3_1_io_ins_left[18] ,
    \ces_3_1_io_ins_left[17] ,
    \ces_3_1_io_ins_left[16] ,
    \ces_3_1_io_ins_left[15] ,
    \ces_3_1_io_ins_left[14] ,
    \ces_3_1_io_ins_left[13] ,
    \ces_3_1_io_ins_left[12] ,
    \ces_3_1_io_ins_left[11] ,
    \ces_3_1_io_ins_left[10] ,
    \ces_3_1_io_ins_left[9] ,
    \ces_3_1_io_ins_left[8] ,
    \ces_3_1_io_ins_left[7] ,
    \ces_3_1_io_ins_left[6] ,
    \ces_3_1_io_ins_left[5] ,
    \ces_3_1_io_ins_left[4] ,
    \ces_3_1_io_ins_left[3] ,
    \ces_3_1_io_ins_left[2] ,
    \ces_3_1_io_ins_left[1] ,
    \ces_3_1_io_ins_left[0] }),
    .io_ins_right({\ces_3_0_io_outs_right[63] ,
    \ces_3_0_io_outs_right[62] ,
    \ces_3_0_io_outs_right[61] ,
    \ces_3_0_io_outs_right[60] ,
    \ces_3_0_io_outs_right[59] ,
    \ces_3_0_io_outs_right[58] ,
    \ces_3_0_io_outs_right[57] ,
    \ces_3_0_io_outs_right[56] ,
    \ces_3_0_io_outs_right[55] ,
    \ces_3_0_io_outs_right[54] ,
    \ces_3_0_io_outs_right[53] ,
    \ces_3_0_io_outs_right[52] ,
    \ces_3_0_io_outs_right[51] ,
    \ces_3_0_io_outs_right[50] ,
    \ces_3_0_io_outs_right[49] ,
    \ces_3_0_io_outs_right[48] ,
    \ces_3_0_io_outs_right[47] ,
    \ces_3_0_io_outs_right[46] ,
    \ces_3_0_io_outs_right[45] ,
    \ces_3_0_io_outs_right[44] ,
    \ces_3_0_io_outs_right[43] ,
    \ces_3_0_io_outs_right[42] ,
    \ces_3_0_io_outs_right[41] ,
    \ces_3_0_io_outs_right[40] ,
    \ces_3_0_io_outs_right[39] ,
    \ces_3_0_io_outs_right[38] ,
    \ces_3_0_io_outs_right[37] ,
    \ces_3_0_io_outs_right[36] ,
    \ces_3_0_io_outs_right[35] ,
    \ces_3_0_io_outs_right[34] ,
    \ces_3_0_io_outs_right[33] ,
    \ces_3_0_io_outs_right[32] ,
    \ces_3_0_io_outs_right[31] ,
    \ces_3_0_io_outs_right[30] ,
    \ces_3_0_io_outs_right[29] ,
    \ces_3_0_io_outs_right[28] ,
    \ces_3_0_io_outs_right[27] ,
    \ces_3_0_io_outs_right[26] ,
    \ces_3_0_io_outs_right[25] ,
    \ces_3_0_io_outs_right[24] ,
    \ces_3_0_io_outs_right[23] ,
    \ces_3_0_io_outs_right[22] ,
    \ces_3_0_io_outs_right[21] ,
    \ces_3_0_io_outs_right[20] ,
    \ces_3_0_io_outs_right[19] ,
    \ces_3_0_io_outs_right[18] ,
    \ces_3_0_io_outs_right[17] ,
    \ces_3_0_io_outs_right[16] ,
    \ces_3_0_io_outs_right[15] ,
    \ces_3_0_io_outs_right[14] ,
    \ces_3_0_io_outs_right[13] ,
    \ces_3_0_io_outs_right[12] ,
    \ces_3_0_io_outs_right[11] ,
    \ces_3_0_io_outs_right[10] ,
    \ces_3_0_io_outs_right[9] ,
    \ces_3_0_io_outs_right[8] ,
    \ces_3_0_io_outs_right[7] ,
    \ces_3_0_io_outs_right[6] ,
    \ces_3_0_io_outs_right[5] ,
    \ces_3_0_io_outs_right[4] ,
    \ces_3_0_io_outs_right[3] ,
    \ces_3_0_io_outs_right[2] ,
    \ces_3_0_io_outs_right[1] ,
    \ces_3_0_io_outs_right[0] }),
    .io_ins_up({\ces_2_1_io_outs_up[63] ,
    \ces_2_1_io_outs_up[62] ,
    \ces_2_1_io_outs_up[61] ,
    \ces_2_1_io_outs_up[60] ,
    \ces_2_1_io_outs_up[59] ,
    \ces_2_1_io_outs_up[58] ,
    \ces_2_1_io_outs_up[57] ,
    \ces_2_1_io_outs_up[56] ,
    \ces_2_1_io_outs_up[55] ,
    \ces_2_1_io_outs_up[54] ,
    \ces_2_1_io_outs_up[53] ,
    \ces_2_1_io_outs_up[52] ,
    \ces_2_1_io_outs_up[51] ,
    \ces_2_1_io_outs_up[50] ,
    \ces_2_1_io_outs_up[49] ,
    \ces_2_1_io_outs_up[48] ,
    \ces_2_1_io_outs_up[47] ,
    \ces_2_1_io_outs_up[46] ,
    \ces_2_1_io_outs_up[45] ,
    \ces_2_1_io_outs_up[44] ,
    \ces_2_1_io_outs_up[43] ,
    \ces_2_1_io_outs_up[42] ,
    \ces_2_1_io_outs_up[41] ,
    \ces_2_1_io_outs_up[40] ,
    \ces_2_1_io_outs_up[39] ,
    \ces_2_1_io_outs_up[38] ,
    \ces_2_1_io_outs_up[37] ,
    \ces_2_1_io_outs_up[36] ,
    \ces_2_1_io_outs_up[35] ,
    \ces_2_1_io_outs_up[34] ,
    \ces_2_1_io_outs_up[33] ,
    \ces_2_1_io_outs_up[32] ,
    \ces_2_1_io_outs_up[31] ,
    \ces_2_1_io_outs_up[30] ,
    \ces_2_1_io_outs_up[29] ,
    \ces_2_1_io_outs_up[28] ,
    \ces_2_1_io_outs_up[27] ,
    \ces_2_1_io_outs_up[26] ,
    \ces_2_1_io_outs_up[25] ,
    \ces_2_1_io_outs_up[24] ,
    \ces_2_1_io_outs_up[23] ,
    \ces_2_1_io_outs_up[22] ,
    \ces_2_1_io_outs_up[21] ,
    \ces_2_1_io_outs_up[20] ,
    \ces_2_1_io_outs_up[19] ,
    \ces_2_1_io_outs_up[18] ,
    \ces_2_1_io_outs_up[17] ,
    \ces_2_1_io_outs_up[16] ,
    \ces_2_1_io_outs_up[15] ,
    \ces_2_1_io_outs_up[14] ,
    \ces_2_1_io_outs_up[13] ,
    \ces_2_1_io_outs_up[12] ,
    \ces_2_1_io_outs_up[11] ,
    \ces_2_1_io_outs_up[10] ,
    \ces_2_1_io_outs_up[9] ,
    \ces_2_1_io_outs_up[8] ,
    \ces_2_1_io_outs_up[7] ,
    \ces_2_1_io_outs_up[6] ,
    \ces_2_1_io_outs_up[5] ,
    \ces_2_1_io_outs_up[4] ,
    \ces_2_1_io_outs_up[3] ,
    \ces_2_1_io_outs_up[2] ,
    \ces_2_1_io_outs_up[1] ,
    \ces_2_1_io_outs_up[0] }),
    .io_outs_down({\ces_2_1_io_ins_down[63] ,
    \ces_2_1_io_ins_down[62] ,
    \ces_2_1_io_ins_down[61] ,
    \ces_2_1_io_ins_down[60] ,
    \ces_2_1_io_ins_down[59] ,
    \ces_2_1_io_ins_down[58] ,
    \ces_2_1_io_ins_down[57] ,
    \ces_2_1_io_ins_down[56] ,
    \ces_2_1_io_ins_down[55] ,
    \ces_2_1_io_ins_down[54] ,
    \ces_2_1_io_ins_down[53] ,
    \ces_2_1_io_ins_down[52] ,
    \ces_2_1_io_ins_down[51] ,
    \ces_2_1_io_ins_down[50] ,
    \ces_2_1_io_ins_down[49] ,
    \ces_2_1_io_ins_down[48] ,
    \ces_2_1_io_ins_down[47] ,
    \ces_2_1_io_ins_down[46] ,
    \ces_2_1_io_ins_down[45] ,
    \ces_2_1_io_ins_down[44] ,
    \ces_2_1_io_ins_down[43] ,
    \ces_2_1_io_ins_down[42] ,
    \ces_2_1_io_ins_down[41] ,
    \ces_2_1_io_ins_down[40] ,
    \ces_2_1_io_ins_down[39] ,
    \ces_2_1_io_ins_down[38] ,
    \ces_2_1_io_ins_down[37] ,
    \ces_2_1_io_ins_down[36] ,
    \ces_2_1_io_ins_down[35] ,
    \ces_2_1_io_ins_down[34] ,
    \ces_2_1_io_ins_down[33] ,
    \ces_2_1_io_ins_down[32] ,
    \ces_2_1_io_ins_down[31] ,
    \ces_2_1_io_ins_down[30] ,
    \ces_2_1_io_ins_down[29] ,
    \ces_2_1_io_ins_down[28] ,
    \ces_2_1_io_ins_down[27] ,
    \ces_2_1_io_ins_down[26] ,
    \ces_2_1_io_ins_down[25] ,
    \ces_2_1_io_ins_down[24] ,
    \ces_2_1_io_ins_down[23] ,
    \ces_2_1_io_ins_down[22] ,
    \ces_2_1_io_ins_down[21] ,
    \ces_2_1_io_ins_down[20] ,
    \ces_2_1_io_ins_down[19] ,
    \ces_2_1_io_ins_down[18] ,
    \ces_2_1_io_ins_down[17] ,
    \ces_2_1_io_ins_down[16] ,
    \ces_2_1_io_ins_down[15] ,
    \ces_2_1_io_ins_down[14] ,
    \ces_2_1_io_ins_down[13] ,
    \ces_2_1_io_ins_down[12] ,
    \ces_2_1_io_ins_down[11] ,
    \ces_2_1_io_ins_down[10] ,
    \ces_2_1_io_ins_down[9] ,
    \ces_2_1_io_ins_down[8] ,
    \ces_2_1_io_ins_down[7] ,
    \ces_2_1_io_ins_down[6] ,
    \ces_2_1_io_ins_down[5] ,
    \ces_2_1_io_ins_down[4] ,
    \ces_2_1_io_ins_down[3] ,
    \ces_2_1_io_ins_down[2] ,
    \ces_2_1_io_ins_down[1] ,
    \ces_2_1_io_ins_down[0] }),
    .io_outs_left({\ces_3_0_io_ins_left[63] ,
    \ces_3_0_io_ins_left[62] ,
    \ces_3_0_io_ins_left[61] ,
    \ces_3_0_io_ins_left[60] ,
    \ces_3_0_io_ins_left[59] ,
    \ces_3_0_io_ins_left[58] ,
    \ces_3_0_io_ins_left[57] ,
    \ces_3_0_io_ins_left[56] ,
    \ces_3_0_io_ins_left[55] ,
    \ces_3_0_io_ins_left[54] ,
    \ces_3_0_io_ins_left[53] ,
    \ces_3_0_io_ins_left[52] ,
    \ces_3_0_io_ins_left[51] ,
    \ces_3_0_io_ins_left[50] ,
    \ces_3_0_io_ins_left[49] ,
    \ces_3_0_io_ins_left[48] ,
    \ces_3_0_io_ins_left[47] ,
    \ces_3_0_io_ins_left[46] ,
    \ces_3_0_io_ins_left[45] ,
    \ces_3_0_io_ins_left[44] ,
    \ces_3_0_io_ins_left[43] ,
    \ces_3_0_io_ins_left[42] ,
    \ces_3_0_io_ins_left[41] ,
    \ces_3_0_io_ins_left[40] ,
    \ces_3_0_io_ins_left[39] ,
    \ces_3_0_io_ins_left[38] ,
    \ces_3_0_io_ins_left[37] ,
    \ces_3_0_io_ins_left[36] ,
    \ces_3_0_io_ins_left[35] ,
    \ces_3_0_io_ins_left[34] ,
    \ces_3_0_io_ins_left[33] ,
    \ces_3_0_io_ins_left[32] ,
    \ces_3_0_io_ins_left[31] ,
    \ces_3_0_io_ins_left[30] ,
    \ces_3_0_io_ins_left[29] ,
    \ces_3_0_io_ins_left[28] ,
    \ces_3_0_io_ins_left[27] ,
    \ces_3_0_io_ins_left[26] ,
    \ces_3_0_io_ins_left[25] ,
    \ces_3_0_io_ins_left[24] ,
    \ces_3_0_io_ins_left[23] ,
    \ces_3_0_io_ins_left[22] ,
    \ces_3_0_io_ins_left[21] ,
    \ces_3_0_io_ins_left[20] ,
    \ces_3_0_io_ins_left[19] ,
    \ces_3_0_io_ins_left[18] ,
    \ces_3_0_io_ins_left[17] ,
    \ces_3_0_io_ins_left[16] ,
    \ces_3_0_io_ins_left[15] ,
    \ces_3_0_io_ins_left[14] ,
    \ces_3_0_io_ins_left[13] ,
    \ces_3_0_io_ins_left[12] ,
    \ces_3_0_io_ins_left[11] ,
    \ces_3_0_io_ins_left[10] ,
    \ces_3_0_io_ins_left[9] ,
    \ces_3_0_io_ins_left[8] ,
    \ces_3_0_io_ins_left[7] ,
    \ces_3_0_io_ins_left[6] ,
    \ces_3_0_io_ins_left[5] ,
    \ces_3_0_io_ins_left[4] ,
    \ces_3_0_io_ins_left[3] ,
    \ces_3_0_io_ins_left[2] ,
    \ces_3_0_io_ins_left[1] ,
    \ces_3_0_io_ins_left[0] }),
    .io_outs_right({\ces_3_1_io_outs_right[63] ,
    \ces_3_1_io_outs_right[62] ,
    \ces_3_1_io_outs_right[61] ,
    \ces_3_1_io_outs_right[60] ,
    \ces_3_1_io_outs_right[59] ,
    \ces_3_1_io_outs_right[58] ,
    \ces_3_1_io_outs_right[57] ,
    \ces_3_1_io_outs_right[56] ,
    \ces_3_1_io_outs_right[55] ,
    \ces_3_1_io_outs_right[54] ,
    \ces_3_1_io_outs_right[53] ,
    \ces_3_1_io_outs_right[52] ,
    \ces_3_1_io_outs_right[51] ,
    \ces_3_1_io_outs_right[50] ,
    \ces_3_1_io_outs_right[49] ,
    \ces_3_1_io_outs_right[48] ,
    \ces_3_1_io_outs_right[47] ,
    \ces_3_1_io_outs_right[46] ,
    \ces_3_1_io_outs_right[45] ,
    \ces_3_1_io_outs_right[44] ,
    \ces_3_1_io_outs_right[43] ,
    \ces_3_1_io_outs_right[42] ,
    \ces_3_1_io_outs_right[41] ,
    \ces_3_1_io_outs_right[40] ,
    \ces_3_1_io_outs_right[39] ,
    \ces_3_1_io_outs_right[38] ,
    \ces_3_1_io_outs_right[37] ,
    \ces_3_1_io_outs_right[36] ,
    \ces_3_1_io_outs_right[35] ,
    \ces_3_1_io_outs_right[34] ,
    \ces_3_1_io_outs_right[33] ,
    \ces_3_1_io_outs_right[32] ,
    \ces_3_1_io_outs_right[31] ,
    \ces_3_1_io_outs_right[30] ,
    \ces_3_1_io_outs_right[29] ,
    \ces_3_1_io_outs_right[28] ,
    \ces_3_1_io_outs_right[27] ,
    \ces_3_1_io_outs_right[26] ,
    \ces_3_1_io_outs_right[25] ,
    \ces_3_1_io_outs_right[24] ,
    \ces_3_1_io_outs_right[23] ,
    \ces_3_1_io_outs_right[22] ,
    \ces_3_1_io_outs_right[21] ,
    \ces_3_1_io_outs_right[20] ,
    \ces_3_1_io_outs_right[19] ,
    \ces_3_1_io_outs_right[18] ,
    \ces_3_1_io_outs_right[17] ,
    \ces_3_1_io_outs_right[16] ,
    \ces_3_1_io_outs_right[15] ,
    \ces_3_1_io_outs_right[14] ,
    \ces_3_1_io_outs_right[13] ,
    \ces_3_1_io_outs_right[12] ,
    \ces_3_1_io_outs_right[11] ,
    \ces_3_1_io_outs_right[10] ,
    \ces_3_1_io_outs_right[9] ,
    \ces_3_1_io_outs_right[8] ,
    \ces_3_1_io_outs_right[7] ,
    \ces_3_1_io_outs_right[6] ,
    \ces_3_1_io_outs_right[5] ,
    \ces_3_1_io_outs_right[4] ,
    \ces_3_1_io_outs_right[3] ,
    \ces_3_1_io_outs_right[2] ,
    \ces_3_1_io_outs_right[1] ,
    \ces_3_1_io_outs_right[0] }),
    .io_outs_up({\ces_3_1_io_outs_up[63] ,
    \ces_3_1_io_outs_up[62] ,
    \ces_3_1_io_outs_up[61] ,
    \ces_3_1_io_outs_up[60] ,
    \ces_3_1_io_outs_up[59] ,
    \ces_3_1_io_outs_up[58] ,
    \ces_3_1_io_outs_up[57] ,
    \ces_3_1_io_outs_up[56] ,
    \ces_3_1_io_outs_up[55] ,
    \ces_3_1_io_outs_up[54] ,
    \ces_3_1_io_outs_up[53] ,
    \ces_3_1_io_outs_up[52] ,
    \ces_3_1_io_outs_up[51] ,
    \ces_3_1_io_outs_up[50] ,
    \ces_3_1_io_outs_up[49] ,
    \ces_3_1_io_outs_up[48] ,
    \ces_3_1_io_outs_up[47] ,
    \ces_3_1_io_outs_up[46] ,
    \ces_3_1_io_outs_up[45] ,
    \ces_3_1_io_outs_up[44] ,
    \ces_3_1_io_outs_up[43] ,
    \ces_3_1_io_outs_up[42] ,
    \ces_3_1_io_outs_up[41] ,
    \ces_3_1_io_outs_up[40] ,
    \ces_3_1_io_outs_up[39] ,
    \ces_3_1_io_outs_up[38] ,
    \ces_3_1_io_outs_up[37] ,
    \ces_3_1_io_outs_up[36] ,
    \ces_3_1_io_outs_up[35] ,
    \ces_3_1_io_outs_up[34] ,
    \ces_3_1_io_outs_up[33] ,
    \ces_3_1_io_outs_up[32] ,
    \ces_3_1_io_outs_up[31] ,
    \ces_3_1_io_outs_up[30] ,
    \ces_3_1_io_outs_up[29] ,
    \ces_3_1_io_outs_up[28] ,
    \ces_3_1_io_outs_up[27] ,
    \ces_3_1_io_outs_up[26] ,
    \ces_3_1_io_outs_up[25] ,
    \ces_3_1_io_outs_up[24] ,
    \ces_3_1_io_outs_up[23] ,
    \ces_3_1_io_outs_up[22] ,
    \ces_3_1_io_outs_up[21] ,
    \ces_3_1_io_outs_up[20] ,
    \ces_3_1_io_outs_up[19] ,
    \ces_3_1_io_outs_up[18] ,
    \ces_3_1_io_outs_up[17] ,
    \ces_3_1_io_outs_up[16] ,
    \ces_3_1_io_outs_up[15] ,
    \ces_3_1_io_outs_up[14] ,
    \ces_3_1_io_outs_up[13] ,
    \ces_3_1_io_outs_up[12] ,
    \ces_3_1_io_outs_up[11] ,
    \ces_3_1_io_outs_up[10] ,
    \ces_3_1_io_outs_up[9] ,
    \ces_3_1_io_outs_up[8] ,
    \ces_3_1_io_outs_up[7] ,
    \ces_3_1_io_outs_up[6] ,
    \ces_3_1_io_outs_up[5] ,
    \ces_3_1_io_outs_up[4] ,
    \ces_3_1_io_outs_up[3] ,
    \ces_3_1_io_outs_up[2] ,
    \ces_3_1_io_outs_up[1] ,
    \ces_3_1_io_outs_up[0] }));
 Element ces_3_2 (.clock(clknet_3_1_0_clock),
    .io_lsbIns_1(ces_3_1_io_lsbOuts_1),
    .io_lsbIns_2(ces_3_1_io_lsbOuts_2),
    .io_lsbIns_3(ces_3_1_io_lsbOuts_3),
    .io_lsbIns_4(ces_3_1_io_lsbOuts_4),
    .io_lsbIns_5(ces_3_1_io_lsbOuts_5),
    .io_lsbIns_6(ces_3_1_io_lsbOuts_6),
    .io_lsbIns_7(ces_3_1_io_lsbOuts_7),
    .io_lsbOuts_0(ces_3_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_2_io_lsbOuts_7),
    .io_ins_down({\ces_3_2_io_ins_down[63] ,
    \ces_3_2_io_ins_down[62] ,
    \ces_3_2_io_ins_down[61] ,
    \ces_3_2_io_ins_down[60] ,
    \ces_3_2_io_ins_down[59] ,
    \ces_3_2_io_ins_down[58] ,
    \ces_3_2_io_ins_down[57] ,
    \ces_3_2_io_ins_down[56] ,
    \ces_3_2_io_ins_down[55] ,
    \ces_3_2_io_ins_down[54] ,
    \ces_3_2_io_ins_down[53] ,
    \ces_3_2_io_ins_down[52] ,
    \ces_3_2_io_ins_down[51] ,
    \ces_3_2_io_ins_down[50] ,
    \ces_3_2_io_ins_down[49] ,
    \ces_3_2_io_ins_down[48] ,
    \ces_3_2_io_ins_down[47] ,
    \ces_3_2_io_ins_down[46] ,
    \ces_3_2_io_ins_down[45] ,
    \ces_3_2_io_ins_down[44] ,
    \ces_3_2_io_ins_down[43] ,
    \ces_3_2_io_ins_down[42] ,
    \ces_3_2_io_ins_down[41] ,
    \ces_3_2_io_ins_down[40] ,
    \ces_3_2_io_ins_down[39] ,
    \ces_3_2_io_ins_down[38] ,
    \ces_3_2_io_ins_down[37] ,
    \ces_3_2_io_ins_down[36] ,
    \ces_3_2_io_ins_down[35] ,
    \ces_3_2_io_ins_down[34] ,
    \ces_3_2_io_ins_down[33] ,
    \ces_3_2_io_ins_down[32] ,
    \ces_3_2_io_ins_down[31] ,
    \ces_3_2_io_ins_down[30] ,
    \ces_3_2_io_ins_down[29] ,
    \ces_3_2_io_ins_down[28] ,
    \ces_3_2_io_ins_down[27] ,
    \ces_3_2_io_ins_down[26] ,
    \ces_3_2_io_ins_down[25] ,
    \ces_3_2_io_ins_down[24] ,
    \ces_3_2_io_ins_down[23] ,
    \ces_3_2_io_ins_down[22] ,
    \ces_3_2_io_ins_down[21] ,
    \ces_3_2_io_ins_down[20] ,
    \ces_3_2_io_ins_down[19] ,
    \ces_3_2_io_ins_down[18] ,
    \ces_3_2_io_ins_down[17] ,
    \ces_3_2_io_ins_down[16] ,
    \ces_3_2_io_ins_down[15] ,
    \ces_3_2_io_ins_down[14] ,
    \ces_3_2_io_ins_down[13] ,
    \ces_3_2_io_ins_down[12] ,
    \ces_3_2_io_ins_down[11] ,
    \ces_3_2_io_ins_down[10] ,
    \ces_3_2_io_ins_down[9] ,
    \ces_3_2_io_ins_down[8] ,
    \ces_3_2_io_ins_down[7] ,
    \ces_3_2_io_ins_down[6] ,
    \ces_3_2_io_ins_down[5] ,
    \ces_3_2_io_ins_down[4] ,
    \ces_3_2_io_ins_down[3] ,
    \ces_3_2_io_ins_down[2] ,
    \ces_3_2_io_ins_down[1] ,
    \ces_3_2_io_ins_down[0] }),
    .io_ins_left({\ces_3_2_io_ins_left[63] ,
    \ces_3_2_io_ins_left[62] ,
    \ces_3_2_io_ins_left[61] ,
    \ces_3_2_io_ins_left[60] ,
    \ces_3_2_io_ins_left[59] ,
    \ces_3_2_io_ins_left[58] ,
    \ces_3_2_io_ins_left[57] ,
    \ces_3_2_io_ins_left[56] ,
    \ces_3_2_io_ins_left[55] ,
    \ces_3_2_io_ins_left[54] ,
    \ces_3_2_io_ins_left[53] ,
    \ces_3_2_io_ins_left[52] ,
    \ces_3_2_io_ins_left[51] ,
    \ces_3_2_io_ins_left[50] ,
    \ces_3_2_io_ins_left[49] ,
    \ces_3_2_io_ins_left[48] ,
    \ces_3_2_io_ins_left[47] ,
    \ces_3_2_io_ins_left[46] ,
    \ces_3_2_io_ins_left[45] ,
    \ces_3_2_io_ins_left[44] ,
    \ces_3_2_io_ins_left[43] ,
    \ces_3_2_io_ins_left[42] ,
    \ces_3_2_io_ins_left[41] ,
    \ces_3_2_io_ins_left[40] ,
    \ces_3_2_io_ins_left[39] ,
    \ces_3_2_io_ins_left[38] ,
    \ces_3_2_io_ins_left[37] ,
    \ces_3_2_io_ins_left[36] ,
    \ces_3_2_io_ins_left[35] ,
    \ces_3_2_io_ins_left[34] ,
    \ces_3_2_io_ins_left[33] ,
    \ces_3_2_io_ins_left[32] ,
    \ces_3_2_io_ins_left[31] ,
    \ces_3_2_io_ins_left[30] ,
    \ces_3_2_io_ins_left[29] ,
    \ces_3_2_io_ins_left[28] ,
    \ces_3_2_io_ins_left[27] ,
    \ces_3_2_io_ins_left[26] ,
    \ces_3_2_io_ins_left[25] ,
    \ces_3_2_io_ins_left[24] ,
    \ces_3_2_io_ins_left[23] ,
    \ces_3_2_io_ins_left[22] ,
    \ces_3_2_io_ins_left[21] ,
    \ces_3_2_io_ins_left[20] ,
    \ces_3_2_io_ins_left[19] ,
    \ces_3_2_io_ins_left[18] ,
    \ces_3_2_io_ins_left[17] ,
    \ces_3_2_io_ins_left[16] ,
    \ces_3_2_io_ins_left[15] ,
    \ces_3_2_io_ins_left[14] ,
    \ces_3_2_io_ins_left[13] ,
    \ces_3_2_io_ins_left[12] ,
    \ces_3_2_io_ins_left[11] ,
    \ces_3_2_io_ins_left[10] ,
    \ces_3_2_io_ins_left[9] ,
    \ces_3_2_io_ins_left[8] ,
    \ces_3_2_io_ins_left[7] ,
    \ces_3_2_io_ins_left[6] ,
    \ces_3_2_io_ins_left[5] ,
    \ces_3_2_io_ins_left[4] ,
    \ces_3_2_io_ins_left[3] ,
    \ces_3_2_io_ins_left[2] ,
    \ces_3_2_io_ins_left[1] ,
    \ces_3_2_io_ins_left[0] }),
    .io_ins_right({\ces_3_1_io_outs_right[63] ,
    \ces_3_1_io_outs_right[62] ,
    \ces_3_1_io_outs_right[61] ,
    \ces_3_1_io_outs_right[60] ,
    \ces_3_1_io_outs_right[59] ,
    \ces_3_1_io_outs_right[58] ,
    \ces_3_1_io_outs_right[57] ,
    \ces_3_1_io_outs_right[56] ,
    \ces_3_1_io_outs_right[55] ,
    \ces_3_1_io_outs_right[54] ,
    \ces_3_1_io_outs_right[53] ,
    \ces_3_1_io_outs_right[52] ,
    \ces_3_1_io_outs_right[51] ,
    \ces_3_1_io_outs_right[50] ,
    \ces_3_1_io_outs_right[49] ,
    \ces_3_1_io_outs_right[48] ,
    \ces_3_1_io_outs_right[47] ,
    \ces_3_1_io_outs_right[46] ,
    \ces_3_1_io_outs_right[45] ,
    \ces_3_1_io_outs_right[44] ,
    \ces_3_1_io_outs_right[43] ,
    \ces_3_1_io_outs_right[42] ,
    \ces_3_1_io_outs_right[41] ,
    \ces_3_1_io_outs_right[40] ,
    \ces_3_1_io_outs_right[39] ,
    \ces_3_1_io_outs_right[38] ,
    \ces_3_1_io_outs_right[37] ,
    \ces_3_1_io_outs_right[36] ,
    \ces_3_1_io_outs_right[35] ,
    \ces_3_1_io_outs_right[34] ,
    \ces_3_1_io_outs_right[33] ,
    \ces_3_1_io_outs_right[32] ,
    \ces_3_1_io_outs_right[31] ,
    \ces_3_1_io_outs_right[30] ,
    \ces_3_1_io_outs_right[29] ,
    \ces_3_1_io_outs_right[28] ,
    \ces_3_1_io_outs_right[27] ,
    \ces_3_1_io_outs_right[26] ,
    \ces_3_1_io_outs_right[25] ,
    \ces_3_1_io_outs_right[24] ,
    \ces_3_1_io_outs_right[23] ,
    \ces_3_1_io_outs_right[22] ,
    \ces_3_1_io_outs_right[21] ,
    \ces_3_1_io_outs_right[20] ,
    \ces_3_1_io_outs_right[19] ,
    \ces_3_1_io_outs_right[18] ,
    \ces_3_1_io_outs_right[17] ,
    \ces_3_1_io_outs_right[16] ,
    \ces_3_1_io_outs_right[15] ,
    \ces_3_1_io_outs_right[14] ,
    \ces_3_1_io_outs_right[13] ,
    \ces_3_1_io_outs_right[12] ,
    \ces_3_1_io_outs_right[11] ,
    \ces_3_1_io_outs_right[10] ,
    \ces_3_1_io_outs_right[9] ,
    \ces_3_1_io_outs_right[8] ,
    \ces_3_1_io_outs_right[7] ,
    \ces_3_1_io_outs_right[6] ,
    \ces_3_1_io_outs_right[5] ,
    \ces_3_1_io_outs_right[4] ,
    \ces_3_1_io_outs_right[3] ,
    \ces_3_1_io_outs_right[2] ,
    \ces_3_1_io_outs_right[1] ,
    \ces_3_1_io_outs_right[0] }),
    .io_ins_up({\ces_2_2_io_outs_up[63] ,
    \ces_2_2_io_outs_up[62] ,
    \ces_2_2_io_outs_up[61] ,
    \ces_2_2_io_outs_up[60] ,
    \ces_2_2_io_outs_up[59] ,
    \ces_2_2_io_outs_up[58] ,
    \ces_2_2_io_outs_up[57] ,
    \ces_2_2_io_outs_up[56] ,
    \ces_2_2_io_outs_up[55] ,
    \ces_2_2_io_outs_up[54] ,
    \ces_2_2_io_outs_up[53] ,
    \ces_2_2_io_outs_up[52] ,
    \ces_2_2_io_outs_up[51] ,
    \ces_2_2_io_outs_up[50] ,
    \ces_2_2_io_outs_up[49] ,
    \ces_2_2_io_outs_up[48] ,
    \ces_2_2_io_outs_up[47] ,
    \ces_2_2_io_outs_up[46] ,
    \ces_2_2_io_outs_up[45] ,
    \ces_2_2_io_outs_up[44] ,
    \ces_2_2_io_outs_up[43] ,
    \ces_2_2_io_outs_up[42] ,
    \ces_2_2_io_outs_up[41] ,
    \ces_2_2_io_outs_up[40] ,
    \ces_2_2_io_outs_up[39] ,
    \ces_2_2_io_outs_up[38] ,
    \ces_2_2_io_outs_up[37] ,
    \ces_2_2_io_outs_up[36] ,
    \ces_2_2_io_outs_up[35] ,
    \ces_2_2_io_outs_up[34] ,
    \ces_2_2_io_outs_up[33] ,
    \ces_2_2_io_outs_up[32] ,
    \ces_2_2_io_outs_up[31] ,
    \ces_2_2_io_outs_up[30] ,
    \ces_2_2_io_outs_up[29] ,
    \ces_2_2_io_outs_up[28] ,
    \ces_2_2_io_outs_up[27] ,
    \ces_2_2_io_outs_up[26] ,
    \ces_2_2_io_outs_up[25] ,
    \ces_2_2_io_outs_up[24] ,
    \ces_2_2_io_outs_up[23] ,
    \ces_2_2_io_outs_up[22] ,
    \ces_2_2_io_outs_up[21] ,
    \ces_2_2_io_outs_up[20] ,
    \ces_2_2_io_outs_up[19] ,
    \ces_2_2_io_outs_up[18] ,
    \ces_2_2_io_outs_up[17] ,
    \ces_2_2_io_outs_up[16] ,
    \ces_2_2_io_outs_up[15] ,
    \ces_2_2_io_outs_up[14] ,
    \ces_2_2_io_outs_up[13] ,
    \ces_2_2_io_outs_up[12] ,
    \ces_2_2_io_outs_up[11] ,
    \ces_2_2_io_outs_up[10] ,
    \ces_2_2_io_outs_up[9] ,
    \ces_2_2_io_outs_up[8] ,
    \ces_2_2_io_outs_up[7] ,
    \ces_2_2_io_outs_up[6] ,
    \ces_2_2_io_outs_up[5] ,
    \ces_2_2_io_outs_up[4] ,
    \ces_2_2_io_outs_up[3] ,
    \ces_2_2_io_outs_up[2] ,
    \ces_2_2_io_outs_up[1] ,
    \ces_2_2_io_outs_up[0] }),
    .io_outs_down({\ces_2_2_io_ins_down[63] ,
    \ces_2_2_io_ins_down[62] ,
    \ces_2_2_io_ins_down[61] ,
    \ces_2_2_io_ins_down[60] ,
    \ces_2_2_io_ins_down[59] ,
    \ces_2_2_io_ins_down[58] ,
    \ces_2_2_io_ins_down[57] ,
    \ces_2_2_io_ins_down[56] ,
    \ces_2_2_io_ins_down[55] ,
    \ces_2_2_io_ins_down[54] ,
    \ces_2_2_io_ins_down[53] ,
    \ces_2_2_io_ins_down[52] ,
    \ces_2_2_io_ins_down[51] ,
    \ces_2_2_io_ins_down[50] ,
    \ces_2_2_io_ins_down[49] ,
    \ces_2_2_io_ins_down[48] ,
    \ces_2_2_io_ins_down[47] ,
    \ces_2_2_io_ins_down[46] ,
    \ces_2_2_io_ins_down[45] ,
    \ces_2_2_io_ins_down[44] ,
    \ces_2_2_io_ins_down[43] ,
    \ces_2_2_io_ins_down[42] ,
    \ces_2_2_io_ins_down[41] ,
    \ces_2_2_io_ins_down[40] ,
    \ces_2_2_io_ins_down[39] ,
    \ces_2_2_io_ins_down[38] ,
    \ces_2_2_io_ins_down[37] ,
    \ces_2_2_io_ins_down[36] ,
    \ces_2_2_io_ins_down[35] ,
    \ces_2_2_io_ins_down[34] ,
    \ces_2_2_io_ins_down[33] ,
    \ces_2_2_io_ins_down[32] ,
    \ces_2_2_io_ins_down[31] ,
    \ces_2_2_io_ins_down[30] ,
    \ces_2_2_io_ins_down[29] ,
    \ces_2_2_io_ins_down[28] ,
    \ces_2_2_io_ins_down[27] ,
    \ces_2_2_io_ins_down[26] ,
    \ces_2_2_io_ins_down[25] ,
    \ces_2_2_io_ins_down[24] ,
    \ces_2_2_io_ins_down[23] ,
    \ces_2_2_io_ins_down[22] ,
    \ces_2_2_io_ins_down[21] ,
    \ces_2_2_io_ins_down[20] ,
    \ces_2_2_io_ins_down[19] ,
    \ces_2_2_io_ins_down[18] ,
    \ces_2_2_io_ins_down[17] ,
    \ces_2_2_io_ins_down[16] ,
    \ces_2_2_io_ins_down[15] ,
    \ces_2_2_io_ins_down[14] ,
    \ces_2_2_io_ins_down[13] ,
    \ces_2_2_io_ins_down[12] ,
    \ces_2_2_io_ins_down[11] ,
    \ces_2_2_io_ins_down[10] ,
    \ces_2_2_io_ins_down[9] ,
    \ces_2_2_io_ins_down[8] ,
    \ces_2_2_io_ins_down[7] ,
    \ces_2_2_io_ins_down[6] ,
    \ces_2_2_io_ins_down[5] ,
    \ces_2_2_io_ins_down[4] ,
    \ces_2_2_io_ins_down[3] ,
    \ces_2_2_io_ins_down[2] ,
    \ces_2_2_io_ins_down[1] ,
    \ces_2_2_io_ins_down[0] }),
    .io_outs_left({\ces_3_1_io_ins_left[63] ,
    \ces_3_1_io_ins_left[62] ,
    \ces_3_1_io_ins_left[61] ,
    \ces_3_1_io_ins_left[60] ,
    \ces_3_1_io_ins_left[59] ,
    \ces_3_1_io_ins_left[58] ,
    \ces_3_1_io_ins_left[57] ,
    \ces_3_1_io_ins_left[56] ,
    \ces_3_1_io_ins_left[55] ,
    \ces_3_1_io_ins_left[54] ,
    \ces_3_1_io_ins_left[53] ,
    \ces_3_1_io_ins_left[52] ,
    \ces_3_1_io_ins_left[51] ,
    \ces_3_1_io_ins_left[50] ,
    \ces_3_1_io_ins_left[49] ,
    \ces_3_1_io_ins_left[48] ,
    \ces_3_1_io_ins_left[47] ,
    \ces_3_1_io_ins_left[46] ,
    \ces_3_1_io_ins_left[45] ,
    \ces_3_1_io_ins_left[44] ,
    \ces_3_1_io_ins_left[43] ,
    \ces_3_1_io_ins_left[42] ,
    \ces_3_1_io_ins_left[41] ,
    \ces_3_1_io_ins_left[40] ,
    \ces_3_1_io_ins_left[39] ,
    \ces_3_1_io_ins_left[38] ,
    \ces_3_1_io_ins_left[37] ,
    \ces_3_1_io_ins_left[36] ,
    \ces_3_1_io_ins_left[35] ,
    \ces_3_1_io_ins_left[34] ,
    \ces_3_1_io_ins_left[33] ,
    \ces_3_1_io_ins_left[32] ,
    \ces_3_1_io_ins_left[31] ,
    \ces_3_1_io_ins_left[30] ,
    \ces_3_1_io_ins_left[29] ,
    \ces_3_1_io_ins_left[28] ,
    \ces_3_1_io_ins_left[27] ,
    \ces_3_1_io_ins_left[26] ,
    \ces_3_1_io_ins_left[25] ,
    \ces_3_1_io_ins_left[24] ,
    \ces_3_1_io_ins_left[23] ,
    \ces_3_1_io_ins_left[22] ,
    \ces_3_1_io_ins_left[21] ,
    \ces_3_1_io_ins_left[20] ,
    \ces_3_1_io_ins_left[19] ,
    \ces_3_1_io_ins_left[18] ,
    \ces_3_1_io_ins_left[17] ,
    \ces_3_1_io_ins_left[16] ,
    \ces_3_1_io_ins_left[15] ,
    \ces_3_1_io_ins_left[14] ,
    \ces_3_1_io_ins_left[13] ,
    \ces_3_1_io_ins_left[12] ,
    \ces_3_1_io_ins_left[11] ,
    \ces_3_1_io_ins_left[10] ,
    \ces_3_1_io_ins_left[9] ,
    \ces_3_1_io_ins_left[8] ,
    \ces_3_1_io_ins_left[7] ,
    \ces_3_1_io_ins_left[6] ,
    \ces_3_1_io_ins_left[5] ,
    \ces_3_1_io_ins_left[4] ,
    \ces_3_1_io_ins_left[3] ,
    \ces_3_1_io_ins_left[2] ,
    \ces_3_1_io_ins_left[1] ,
    \ces_3_1_io_ins_left[0] }),
    .io_outs_right({\ces_3_2_io_outs_right[63] ,
    \ces_3_2_io_outs_right[62] ,
    \ces_3_2_io_outs_right[61] ,
    \ces_3_2_io_outs_right[60] ,
    \ces_3_2_io_outs_right[59] ,
    \ces_3_2_io_outs_right[58] ,
    \ces_3_2_io_outs_right[57] ,
    \ces_3_2_io_outs_right[56] ,
    \ces_3_2_io_outs_right[55] ,
    \ces_3_2_io_outs_right[54] ,
    \ces_3_2_io_outs_right[53] ,
    \ces_3_2_io_outs_right[52] ,
    \ces_3_2_io_outs_right[51] ,
    \ces_3_2_io_outs_right[50] ,
    \ces_3_2_io_outs_right[49] ,
    \ces_3_2_io_outs_right[48] ,
    \ces_3_2_io_outs_right[47] ,
    \ces_3_2_io_outs_right[46] ,
    \ces_3_2_io_outs_right[45] ,
    \ces_3_2_io_outs_right[44] ,
    \ces_3_2_io_outs_right[43] ,
    \ces_3_2_io_outs_right[42] ,
    \ces_3_2_io_outs_right[41] ,
    \ces_3_2_io_outs_right[40] ,
    \ces_3_2_io_outs_right[39] ,
    \ces_3_2_io_outs_right[38] ,
    \ces_3_2_io_outs_right[37] ,
    \ces_3_2_io_outs_right[36] ,
    \ces_3_2_io_outs_right[35] ,
    \ces_3_2_io_outs_right[34] ,
    \ces_3_2_io_outs_right[33] ,
    \ces_3_2_io_outs_right[32] ,
    \ces_3_2_io_outs_right[31] ,
    \ces_3_2_io_outs_right[30] ,
    \ces_3_2_io_outs_right[29] ,
    \ces_3_2_io_outs_right[28] ,
    \ces_3_2_io_outs_right[27] ,
    \ces_3_2_io_outs_right[26] ,
    \ces_3_2_io_outs_right[25] ,
    \ces_3_2_io_outs_right[24] ,
    \ces_3_2_io_outs_right[23] ,
    \ces_3_2_io_outs_right[22] ,
    \ces_3_2_io_outs_right[21] ,
    \ces_3_2_io_outs_right[20] ,
    \ces_3_2_io_outs_right[19] ,
    \ces_3_2_io_outs_right[18] ,
    \ces_3_2_io_outs_right[17] ,
    \ces_3_2_io_outs_right[16] ,
    \ces_3_2_io_outs_right[15] ,
    \ces_3_2_io_outs_right[14] ,
    \ces_3_2_io_outs_right[13] ,
    \ces_3_2_io_outs_right[12] ,
    \ces_3_2_io_outs_right[11] ,
    \ces_3_2_io_outs_right[10] ,
    \ces_3_2_io_outs_right[9] ,
    \ces_3_2_io_outs_right[8] ,
    \ces_3_2_io_outs_right[7] ,
    \ces_3_2_io_outs_right[6] ,
    \ces_3_2_io_outs_right[5] ,
    \ces_3_2_io_outs_right[4] ,
    \ces_3_2_io_outs_right[3] ,
    \ces_3_2_io_outs_right[2] ,
    \ces_3_2_io_outs_right[1] ,
    \ces_3_2_io_outs_right[0] }),
    .io_outs_up({\ces_3_2_io_outs_up[63] ,
    \ces_3_2_io_outs_up[62] ,
    \ces_3_2_io_outs_up[61] ,
    \ces_3_2_io_outs_up[60] ,
    \ces_3_2_io_outs_up[59] ,
    \ces_3_2_io_outs_up[58] ,
    \ces_3_2_io_outs_up[57] ,
    \ces_3_2_io_outs_up[56] ,
    \ces_3_2_io_outs_up[55] ,
    \ces_3_2_io_outs_up[54] ,
    \ces_3_2_io_outs_up[53] ,
    \ces_3_2_io_outs_up[52] ,
    \ces_3_2_io_outs_up[51] ,
    \ces_3_2_io_outs_up[50] ,
    \ces_3_2_io_outs_up[49] ,
    \ces_3_2_io_outs_up[48] ,
    \ces_3_2_io_outs_up[47] ,
    \ces_3_2_io_outs_up[46] ,
    \ces_3_2_io_outs_up[45] ,
    \ces_3_2_io_outs_up[44] ,
    \ces_3_2_io_outs_up[43] ,
    \ces_3_2_io_outs_up[42] ,
    \ces_3_2_io_outs_up[41] ,
    \ces_3_2_io_outs_up[40] ,
    \ces_3_2_io_outs_up[39] ,
    \ces_3_2_io_outs_up[38] ,
    \ces_3_2_io_outs_up[37] ,
    \ces_3_2_io_outs_up[36] ,
    \ces_3_2_io_outs_up[35] ,
    \ces_3_2_io_outs_up[34] ,
    \ces_3_2_io_outs_up[33] ,
    \ces_3_2_io_outs_up[32] ,
    \ces_3_2_io_outs_up[31] ,
    \ces_3_2_io_outs_up[30] ,
    \ces_3_2_io_outs_up[29] ,
    \ces_3_2_io_outs_up[28] ,
    \ces_3_2_io_outs_up[27] ,
    \ces_3_2_io_outs_up[26] ,
    \ces_3_2_io_outs_up[25] ,
    \ces_3_2_io_outs_up[24] ,
    \ces_3_2_io_outs_up[23] ,
    \ces_3_2_io_outs_up[22] ,
    \ces_3_2_io_outs_up[21] ,
    \ces_3_2_io_outs_up[20] ,
    \ces_3_2_io_outs_up[19] ,
    \ces_3_2_io_outs_up[18] ,
    \ces_3_2_io_outs_up[17] ,
    \ces_3_2_io_outs_up[16] ,
    \ces_3_2_io_outs_up[15] ,
    \ces_3_2_io_outs_up[14] ,
    \ces_3_2_io_outs_up[13] ,
    \ces_3_2_io_outs_up[12] ,
    \ces_3_2_io_outs_up[11] ,
    \ces_3_2_io_outs_up[10] ,
    \ces_3_2_io_outs_up[9] ,
    \ces_3_2_io_outs_up[8] ,
    \ces_3_2_io_outs_up[7] ,
    \ces_3_2_io_outs_up[6] ,
    \ces_3_2_io_outs_up[5] ,
    \ces_3_2_io_outs_up[4] ,
    \ces_3_2_io_outs_up[3] ,
    \ces_3_2_io_outs_up[2] ,
    \ces_3_2_io_outs_up[1] ,
    \ces_3_2_io_outs_up[0] }));
 Element ces_3_3 (.clock(clknet_3_1_0_clock),
    .io_lsbIns_1(ces_3_2_io_lsbOuts_1),
    .io_lsbIns_2(ces_3_2_io_lsbOuts_2),
    .io_lsbIns_3(ces_3_2_io_lsbOuts_3),
    .io_lsbIns_4(ces_3_2_io_lsbOuts_4),
    .io_lsbIns_5(ces_3_2_io_lsbOuts_5),
    .io_lsbIns_6(ces_3_2_io_lsbOuts_6),
    .io_lsbIns_7(ces_3_2_io_lsbOuts_7),
    .io_lsbOuts_0(ces_3_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_3_io_lsbOuts_7),
    .io_ins_down({\ces_3_3_io_ins_down[63] ,
    \ces_3_3_io_ins_down[62] ,
    \ces_3_3_io_ins_down[61] ,
    \ces_3_3_io_ins_down[60] ,
    \ces_3_3_io_ins_down[59] ,
    \ces_3_3_io_ins_down[58] ,
    \ces_3_3_io_ins_down[57] ,
    \ces_3_3_io_ins_down[56] ,
    \ces_3_3_io_ins_down[55] ,
    \ces_3_3_io_ins_down[54] ,
    \ces_3_3_io_ins_down[53] ,
    \ces_3_3_io_ins_down[52] ,
    \ces_3_3_io_ins_down[51] ,
    \ces_3_3_io_ins_down[50] ,
    \ces_3_3_io_ins_down[49] ,
    \ces_3_3_io_ins_down[48] ,
    \ces_3_3_io_ins_down[47] ,
    \ces_3_3_io_ins_down[46] ,
    \ces_3_3_io_ins_down[45] ,
    \ces_3_3_io_ins_down[44] ,
    \ces_3_3_io_ins_down[43] ,
    \ces_3_3_io_ins_down[42] ,
    \ces_3_3_io_ins_down[41] ,
    \ces_3_3_io_ins_down[40] ,
    \ces_3_3_io_ins_down[39] ,
    \ces_3_3_io_ins_down[38] ,
    \ces_3_3_io_ins_down[37] ,
    \ces_3_3_io_ins_down[36] ,
    \ces_3_3_io_ins_down[35] ,
    \ces_3_3_io_ins_down[34] ,
    \ces_3_3_io_ins_down[33] ,
    \ces_3_3_io_ins_down[32] ,
    \ces_3_3_io_ins_down[31] ,
    \ces_3_3_io_ins_down[30] ,
    \ces_3_3_io_ins_down[29] ,
    \ces_3_3_io_ins_down[28] ,
    \ces_3_3_io_ins_down[27] ,
    \ces_3_3_io_ins_down[26] ,
    \ces_3_3_io_ins_down[25] ,
    \ces_3_3_io_ins_down[24] ,
    \ces_3_3_io_ins_down[23] ,
    \ces_3_3_io_ins_down[22] ,
    \ces_3_3_io_ins_down[21] ,
    \ces_3_3_io_ins_down[20] ,
    \ces_3_3_io_ins_down[19] ,
    \ces_3_3_io_ins_down[18] ,
    \ces_3_3_io_ins_down[17] ,
    \ces_3_3_io_ins_down[16] ,
    \ces_3_3_io_ins_down[15] ,
    \ces_3_3_io_ins_down[14] ,
    \ces_3_3_io_ins_down[13] ,
    \ces_3_3_io_ins_down[12] ,
    \ces_3_3_io_ins_down[11] ,
    \ces_3_3_io_ins_down[10] ,
    \ces_3_3_io_ins_down[9] ,
    \ces_3_3_io_ins_down[8] ,
    \ces_3_3_io_ins_down[7] ,
    \ces_3_3_io_ins_down[6] ,
    \ces_3_3_io_ins_down[5] ,
    \ces_3_3_io_ins_down[4] ,
    \ces_3_3_io_ins_down[3] ,
    \ces_3_3_io_ins_down[2] ,
    \ces_3_3_io_ins_down[1] ,
    \ces_3_3_io_ins_down[0] }),
    .io_ins_left({\ces_3_3_io_ins_left[63] ,
    \ces_3_3_io_ins_left[62] ,
    \ces_3_3_io_ins_left[61] ,
    \ces_3_3_io_ins_left[60] ,
    \ces_3_3_io_ins_left[59] ,
    \ces_3_3_io_ins_left[58] ,
    \ces_3_3_io_ins_left[57] ,
    \ces_3_3_io_ins_left[56] ,
    \ces_3_3_io_ins_left[55] ,
    \ces_3_3_io_ins_left[54] ,
    \ces_3_3_io_ins_left[53] ,
    \ces_3_3_io_ins_left[52] ,
    \ces_3_3_io_ins_left[51] ,
    \ces_3_3_io_ins_left[50] ,
    \ces_3_3_io_ins_left[49] ,
    \ces_3_3_io_ins_left[48] ,
    \ces_3_3_io_ins_left[47] ,
    \ces_3_3_io_ins_left[46] ,
    \ces_3_3_io_ins_left[45] ,
    \ces_3_3_io_ins_left[44] ,
    \ces_3_3_io_ins_left[43] ,
    \ces_3_3_io_ins_left[42] ,
    \ces_3_3_io_ins_left[41] ,
    \ces_3_3_io_ins_left[40] ,
    \ces_3_3_io_ins_left[39] ,
    \ces_3_3_io_ins_left[38] ,
    \ces_3_3_io_ins_left[37] ,
    \ces_3_3_io_ins_left[36] ,
    \ces_3_3_io_ins_left[35] ,
    \ces_3_3_io_ins_left[34] ,
    \ces_3_3_io_ins_left[33] ,
    \ces_3_3_io_ins_left[32] ,
    \ces_3_3_io_ins_left[31] ,
    \ces_3_3_io_ins_left[30] ,
    \ces_3_3_io_ins_left[29] ,
    \ces_3_3_io_ins_left[28] ,
    \ces_3_3_io_ins_left[27] ,
    \ces_3_3_io_ins_left[26] ,
    \ces_3_3_io_ins_left[25] ,
    \ces_3_3_io_ins_left[24] ,
    \ces_3_3_io_ins_left[23] ,
    \ces_3_3_io_ins_left[22] ,
    \ces_3_3_io_ins_left[21] ,
    \ces_3_3_io_ins_left[20] ,
    \ces_3_3_io_ins_left[19] ,
    \ces_3_3_io_ins_left[18] ,
    \ces_3_3_io_ins_left[17] ,
    \ces_3_3_io_ins_left[16] ,
    \ces_3_3_io_ins_left[15] ,
    \ces_3_3_io_ins_left[14] ,
    \ces_3_3_io_ins_left[13] ,
    \ces_3_3_io_ins_left[12] ,
    \ces_3_3_io_ins_left[11] ,
    \ces_3_3_io_ins_left[10] ,
    \ces_3_3_io_ins_left[9] ,
    \ces_3_3_io_ins_left[8] ,
    \ces_3_3_io_ins_left[7] ,
    \ces_3_3_io_ins_left[6] ,
    \ces_3_3_io_ins_left[5] ,
    \ces_3_3_io_ins_left[4] ,
    \ces_3_3_io_ins_left[3] ,
    \ces_3_3_io_ins_left[2] ,
    \ces_3_3_io_ins_left[1] ,
    \ces_3_3_io_ins_left[0] }),
    .io_ins_right({\ces_3_2_io_outs_right[63] ,
    \ces_3_2_io_outs_right[62] ,
    \ces_3_2_io_outs_right[61] ,
    \ces_3_2_io_outs_right[60] ,
    \ces_3_2_io_outs_right[59] ,
    \ces_3_2_io_outs_right[58] ,
    \ces_3_2_io_outs_right[57] ,
    \ces_3_2_io_outs_right[56] ,
    \ces_3_2_io_outs_right[55] ,
    \ces_3_2_io_outs_right[54] ,
    \ces_3_2_io_outs_right[53] ,
    \ces_3_2_io_outs_right[52] ,
    \ces_3_2_io_outs_right[51] ,
    \ces_3_2_io_outs_right[50] ,
    \ces_3_2_io_outs_right[49] ,
    \ces_3_2_io_outs_right[48] ,
    \ces_3_2_io_outs_right[47] ,
    \ces_3_2_io_outs_right[46] ,
    \ces_3_2_io_outs_right[45] ,
    \ces_3_2_io_outs_right[44] ,
    \ces_3_2_io_outs_right[43] ,
    \ces_3_2_io_outs_right[42] ,
    \ces_3_2_io_outs_right[41] ,
    \ces_3_2_io_outs_right[40] ,
    \ces_3_2_io_outs_right[39] ,
    \ces_3_2_io_outs_right[38] ,
    \ces_3_2_io_outs_right[37] ,
    \ces_3_2_io_outs_right[36] ,
    \ces_3_2_io_outs_right[35] ,
    \ces_3_2_io_outs_right[34] ,
    \ces_3_2_io_outs_right[33] ,
    \ces_3_2_io_outs_right[32] ,
    \ces_3_2_io_outs_right[31] ,
    \ces_3_2_io_outs_right[30] ,
    \ces_3_2_io_outs_right[29] ,
    \ces_3_2_io_outs_right[28] ,
    \ces_3_2_io_outs_right[27] ,
    \ces_3_2_io_outs_right[26] ,
    \ces_3_2_io_outs_right[25] ,
    \ces_3_2_io_outs_right[24] ,
    \ces_3_2_io_outs_right[23] ,
    \ces_3_2_io_outs_right[22] ,
    \ces_3_2_io_outs_right[21] ,
    \ces_3_2_io_outs_right[20] ,
    \ces_3_2_io_outs_right[19] ,
    \ces_3_2_io_outs_right[18] ,
    \ces_3_2_io_outs_right[17] ,
    \ces_3_2_io_outs_right[16] ,
    \ces_3_2_io_outs_right[15] ,
    \ces_3_2_io_outs_right[14] ,
    \ces_3_2_io_outs_right[13] ,
    \ces_3_2_io_outs_right[12] ,
    \ces_3_2_io_outs_right[11] ,
    \ces_3_2_io_outs_right[10] ,
    \ces_3_2_io_outs_right[9] ,
    \ces_3_2_io_outs_right[8] ,
    \ces_3_2_io_outs_right[7] ,
    \ces_3_2_io_outs_right[6] ,
    \ces_3_2_io_outs_right[5] ,
    \ces_3_2_io_outs_right[4] ,
    \ces_3_2_io_outs_right[3] ,
    \ces_3_2_io_outs_right[2] ,
    \ces_3_2_io_outs_right[1] ,
    \ces_3_2_io_outs_right[0] }),
    .io_ins_up({\ces_2_3_io_outs_up[63] ,
    \ces_2_3_io_outs_up[62] ,
    \ces_2_3_io_outs_up[61] ,
    \ces_2_3_io_outs_up[60] ,
    \ces_2_3_io_outs_up[59] ,
    \ces_2_3_io_outs_up[58] ,
    \ces_2_3_io_outs_up[57] ,
    \ces_2_3_io_outs_up[56] ,
    \ces_2_3_io_outs_up[55] ,
    \ces_2_3_io_outs_up[54] ,
    \ces_2_3_io_outs_up[53] ,
    \ces_2_3_io_outs_up[52] ,
    \ces_2_3_io_outs_up[51] ,
    \ces_2_3_io_outs_up[50] ,
    \ces_2_3_io_outs_up[49] ,
    \ces_2_3_io_outs_up[48] ,
    \ces_2_3_io_outs_up[47] ,
    \ces_2_3_io_outs_up[46] ,
    \ces_2_3_io_outs_up[45] ,
    \ces_2_3_io_outs_up[44] ,
    \ces_2_3_io_outs_up[43] ,
    \ces_2_3_io_outs_up[42] ,
    \ces_2_3_io_outs_up[41] ,
    \ces_2_3_io_outs_up[40] ,
    \ces_2_3_io_outs_up[39] ,
    \ces_2_3_io_outs_up[38] ,
    \ces_2_3_io_outs_up[37] ,
    \ces_2_3_io_outs_up[36] ,
    \ces_2_3_io_outs_up[35] ,
    \ces_2_3_io_outs_up[34] ,
    \ces_2_3_io_outs_up[33] ,
    \ces_2_3_io_outs_up[32] ,
    \ces_2_3_io_outs_up[31] ,
    \ces_2_3_io_outs_up[30] ,
    \ces_2_3_io_outs_up[29] ,
    \ces_2_3_io_outs_up[28] ,
    \ces_2_3_io_outs_up[27] ,
    \ces_2_3_io_outs_up[26] ,
    \ces_2_3_io_outs_up[25] ,
    \ces_2_3_io_outs_up[24] ,
    \ces_2_3_io_outs_up[23] ,
    \ces_2_3_io_outs_up[22] ,
    \ces_2_3_io_outs_up[21] ,
    \ces_2_3_io_outs_up[20] ,
    \ces_2_3_io_outs_up[19] ,
    \ces_2_3_io_outs_up[18] ,
    \ces_2_3_io_outs_up[17] ,
    \ces_2_3_io_outs_up[16] ,
    \ces_2_3_io_outs_up[15] ,
    \ces_2_3_io_outs_up[14] ,
    \ces_2_3_io_outs_up[13] ,
    \ces_2_3_io_outs_up[12] ,
    \ces_2_3_io_outs_up[11] ,
    \ces_2_3_io_outs_up[10] ,
    \ces_2_3_io_outs_up[9] ,
    \ces_2_3_io_outs_up[8] ,
    \ces_2_3_io_outs_up[7] ,
    \ces_2_3_io_outs_up[6] ,
    \ces_2_3_io_outs_up[5] ,
    \ces_2_3_io_outs_up[4] ,
    \ces_2_3_io_outs_up[3] ,
    \ces_2_3_io_outs_up[2] ,
    \ces_2_3_io_outs_up[1] ,
    \ces_2_3_io_outs_up[0] }),
    .io_outs_down({\ces_2_3_io_ins_down[63] ,
    \ces_2_3_io_ins_down[62] ,
    \ces_2_3_io_ins_down[61] ,
    \ces_2_3_io_ins_down[60] ,
    \ces_2_3_io_ins_down[59] ,
    \ces_2_3_io_ins_down[58] ,
    \ces_2_3_io_ins_down[57] ,
    \ces_2_3_io_ins_down[56] ,
    \ces_2_3_io_ins_down[55] ,
    \ces_2_3_io_ins_down[54] ,
    \ces_2_3_io_ins_down[53] ,
    \ces_2_3_io_ins_down[52] ,
    \ces_2_3_io_ins_down[51] ,
    \ces_2_3_io_ins_down[50] ,
    \ces_2_3_io_ins_down[49] ,
    \ces_2_3_io_ins_down[48] ,
    \ces_2_3_io_ins_down[47] ,
    \ces_2_3_io_ins_down[46] ,
    \ces_2_3_io_ins_down[45] ,
    \ces_2_3_io_ins_down[44] ,
    \ces_2_3_io_ins_down[43] ,
    \ces_2_3_io_ins_down[42] ,
    \ces_2_3_io_ins_down[41] ,
    \ces_2_3_io_ins_down[40] ,
    \ces_2_3_io_ins_down[39] ,
    \ces_2_3_io_ins_down[38] ,
    \ces_2_3_io_ins_down[37] ,
    \ces_2_3_io_ins_down[36] ,
    \ces_2_3_io_ins_down[35] ,
    \ces_2_3_io_ins_down[34] ,
    \ces_2_3_io_ins_down[33] ,
    \ces_2_3_io_ins_down[32] ,
    \ces_2_3_io_ins_down[31] ,
    \ces_2_3_io_ins_down[30] ,
    \ces_2_3_io_ins_down[29] ,
    \ces_2_3_io_ins_down[28] ,
    \ces_2_3_io_ins_down[27] ,
    \ces_2_3_io_ins_down[26] ,
    \ces_2_3_io_ins_down[25] ,
    \ces_2_3_io_ins_down[24] ,
    \ces_2_3_io_ins_down[23] ,
    \ces_2_3_io_ins_down[22] ,
    \ces_2_3_io_ins_down[21] ,
    \ces_2_3_io_ins_down[20] ,
    \ces_2_3_io_ins_down[19] ,
    \ces_2_3_io_ins_down[18] ,
    \ces_2_3_io_ins_down[17] ,
    \ces_2_3_io_ins_down[16] ,
    \ces_2_3_io_ins_down[15] ,
    \ces_2_3_io_ins_down[14] ,
    \ces_2_3_io_ins_down[13] ,
    \ces_2_3_io_ins_down[12] ,
    \ces_2_3_io_ins_down[11] ,
    \ces_2_3_io_ins_down[10] ,
    \ces_2_3_io_ins_down[9] ,
    \ces_2_3_io_ins_down[8] ,
    \ces_2_3_io_ins_down[7] ,
    \ces_2_3_io_ins_down[6] ,
    \ces_2_3_io_ins_down[5] ,
    \ces_2_3_io_ins_down[4] ,
    \ces_2_3_io_ins_down[3] ,
    \ces_2_3_io_ins_down[2] ,
    \ces_2_3_io_ins_down[1] ,
    \ces_2_3_io_ins_down[0] }),
    .io_outs_left({\ces_3_2_io_ins_left[63] ,
    \ces_3_2_io_ins_left[62] ,
    \ces_3_2_io_ins_left[61] ,
    \ces_3_2_io_ins_left[60] ,
    \ces_3_2_io_ins_left[59] ,
    \ces_3_2_io_ins_left[58] ,
    \ces_3_2_io_ins_left[57] ,
    \ces_3_2_io_ins_left[56] ,
    \ces_3_2_io_ins_left[55] ,
    \ces_3_2_io_ins_left[54] ,
    \ces_3_2_io_ins_left[53] ,
    \ces_3_2_io_ins_left[52] ,
    \ces_3_2_io_ins_left[51] ,
    \ces_3_2_io_ins_left[50] ,
    \ces_3_2_io_ins_left[49] ,
    \ces_3_2_io_ins_left[48] ,
    \ces_3_2_io_ins_left[47] ,
    \ces_3_2_io_ins_left[46] ,
    \ces_3_2_io_ins_left[45] ,
    \ces_3_2_io_ins_left[44] ,
    \ces_3_2_io_ins_left[43] ,
    \ces_3_2_io_ins_left[42] ,
    \ces_3_2_io_ins_left[41] ,
    \ces_3_2_io_ins_left[40] ,
    \ces_3_2_io_ins_left[39] ,
    \ces_3_2_io_ins_left[38] ,
    \ces_3_2_io_ins_left[37] ,
    \ces_3_2_io_ins_left[36] ,
    \ces_3_2_io_ins_left[35] ,
    \ces_3_2_io_ins_left[34] ,
    \ces_3_2_io_ins_left[33] ,
    \ces_3_2_io_ins_left[32] ,
    \ces_3_2_io_ins_left[31] ,
    \ces_3_2_io_ins_left[30] ,
    \ces_3_2_io_ins_left[29] ,
    \ces_3_2_io_ins_left[28] ,
    \ces_3_2_io_ins_left[27] ,
    \ces_3_2_io_ins_left[26] ,
    \ces_3_2_io_ins_left[25] ,
    \ces_3_2_io_ins_left[24] ,
    \ces_3_2_io_ins_left[23] ,
    \ces_3_2_io_ins_left[22] ,
    \ces_3_2_io_ins_left[21] ,
    \ces_3_2_io_ins_left[20] ,
    \ces_3_2_io_ins_left[19] ,
    \ces_3_2_io_ins_left[18] ,
    \ces_3_2_io_ins_left[17] ,
    \ces_3_2_io_ins_left[16] ,
    \ces_3_2_io_ins_left[15] ,
    \ces_3_2_io_ins_left[14] ,
    \ces_3_2_io_ins_left[13] ,
    \ces_3_2_io_ins_left[12] ,
    \ces_3_2_io_ins_left[11] ,
    \ces_3_2_io_ins_left[10] ,
    \ces_3_2_io_ins_left[9] ,
    \ces_3_2_io_ins_left[8] ,
    \ces_3_2_io_ins_left[7] ,
    \ces_3_2_io_ins_left[6] ,
    \ces_3_2_io_ins_left[5] ,
    \ces_3_2_io_ins_left[4] ,
    \ces_3_2_io_ins_left[3] ,
    \ces_3_2_io_ins_left[2] ,
    \ces_3_2_io_ins_left[1] ,
    \ces_3_2_io_ins_left[0] }),
    .io_outs_right({\ces_3_3_io_outs_right[63] ,
    \ces_3_3_io_outs_right[62] ,
    \ces_3_3_io_outs_right[61] ,
    \ces_3_3_io_outs_right[60] ,
    \ces_3_3_io_outs_right[59] ,
    \ces_3_3_io_outs_right[58] ,
    \ces_3_3_io_outs_right[57] ,
    \ces_3_3_io_outs_right[56] ,
    \ces_3_3_io_outs_right[55] ,
    \ces_3_3_io_outs_right[54] ,
    \ces_3_3_io_outs_right[53] ,
    \ces_3_3_io_outs_right[52] ,
    \ces_3_3_io_outs_right[51] ,
    \ces_3_3_io_outs_right[50] ,
    \ces_3_3_io_outs_right[49] ,
    \ces_3_3_io_outs_right[48] ,
    \ces_3_3_io_outs_right[47] ,
    \ces_3_3_io_outs_right[46] ,
    \ces_3_3_io_outs_right[45] ,
    \ces_3_3_io_outs_right[44] ,
    \ces_3_3_io_outs_right[43] ,
    \ces_3_3_io_outs_right[42] ,
    \ces_3_3_io_outs_right[41] ,
    \ces_3_3_io_outs_right[40] ,
    \ces_3_3_io_outs_right[39] ,
    \ces_3_3_io_outs_right[38] ,
    \ces_3_3_io_outs_right[37] ,
    \ces_3_3_io_outs_right[36] ,
    \ces_3_3_io_outs_right[35] ,
    \ces_3_3_io_outs_right[34] ,
    \ces_3_3_io_outs_right[33] ,
    \ces_3_3_io_outs_right[32] ,
    \ces_3_3_io_outs_right[31] ,
    \ces_3_3_io_outs_right[30] ,
    \ces_3_3_io_outs_right[29] ,
    \ces_3_3_io_outs_right[28] ,
    \ces_3_3_io_outs_right[27] ,
    \ces_3_3_io_outs_right[26] ,
    \ces_3_3_io_outs_right[25] ,
    \ces_3_3_io_outs_right[24] ,
    \ces_3_3_io_outs_right[23] ,
    \ces_3_3_io_outs_right[22] ,
    \ces_3_3_io_outs_right[21] ,
    \ces_3_3_io_outs_right[20] ,
    \ces_3_3_io_outs_right[19] ,
    \ces_3_3_io_outs_right[18] ,
    \ces_3_3_io_outs_right[17] ,
    \ces_3_3_io_outs_right[16] ,
    \ces_3_3_io_outs_right[15] ,
    \ces_3_3_io_outs_right[14] ,
    \ces_3_3_io_outs_right[13] ,
    \ces_3_3_io_outs_right[12] ,
    \ces_3_3_io_outs_right[11] ,
    \ces_3_3_io_outs_right[10] ,
    \ces_3_3_io_outs_right[9] ,
    \ces_3_3_io_outs_right[8] ,
    \ces_3_3_io_outs_right[7] ,
    \ces_3_3_io_outs_right[6] ,
    \ces_3_3_io_outs_right[5] ,
    \ces_3_3_io_outs_right[4] ,
    \ces_3_3_io_outs_right[3] ,
    \ces_3_3_io_outs_right[2] ,
    \ces_3_3_io_outs_right[1] ,
    \ces_3_3_io_outs_right[0] }),
    .io_outs_up({\ces_3_3_io_outs_up[63] ,
    \ces_3_3_io_outs_up[62] ,
    \ces_3_3_io_outs_up[61] ,
    \ces_3_3_io_outs_up[60] ,
    \ces_3_3_io_outs_up[59] ,
    \ces_3_3_io_outs_up[58] ,
    \ces_3_3_io_outs_up[57] ,
    \ces_3_3_io_outs_up[56] ,
    \ces_3_3_io_outs_up[55] ,
    \ces_3_3_io_outs_up[54] ,
    \ces_3_3_io_outs_up[53] ,
    \ces_3_3_io_outs_up[52] ,
    \ces_3_3_io_outs_up[51] ,
    \ces_3_3_io_outs_up[50] ,
    \ces_3_3_io_outs_up[49] ,
    \ces_3_3_io_outs_up[48] ,
    \ces_3_3_io_outs_up[47] ,
    \ces_3_3_io_outs_up[46] ,
    \ces_3_3_io_outs_up[45] ,
    \ces_3_3_io_outs_up[44] ,
    \ces_3_3_io_outs_up[43] ,
    \ces_3_3_io_outs_up[42] ,
    \ces_3_3_io_outs_up[41] ,
    \ces_3_3_io_outs_up[40] ,
    \ces_3_3_io_outs_up[39] ,
    \ces_3_3_io_outs_up[38] ,
    \ces_3_3_io_outs_up[37] ,
    \ces_3_3_io_outs_up[36] ,
    \ces_3_3_io_outs_up[35] ,
    \ces_3_3_io_outs_up[34] ,
    \ces_3_3_io_outs_up[33] ,
    \ces_3_3_io_outs_up[32] ,
    \ces_3_3_io_outs_up[31] ,
    \ces_3_3_io_outs_up[30] ,
    \ces_3_3_io_outs_up[29] ,
    \ces_3_3_io_outs_up[28] ,
    \ces_3_3_io_outs_up[27] ,
    \ces_3_3_io_outs_up[26] ,
    \ces_3_3_io_outs_up[25] ,
    \ces_3_3_io_outs_up[24] ,
    \ces_3_3_io_outs_up[23] ,
    \ces_3_3_io_outs_up[22] ,
    \ces_3_3_io_outs_up[21] ,
    \ces_3_3_io_outs_up[20] ,
    \ces_3_3_io_outs_up[19] ,
    \ces_3_3_io_outs_up[18] ,
    \ces_3_3_io_outs_up[17] ,
    \ces_3_3_io_outs_up[16] ,
    \ces_3_3_io_outs_up[15] ,
    \ces_3_3_io_outs_up[14] ,
    \ces_3_3_io_outs_up[13] ,
    \ces_3_3_io_outs_up[12] ,
    \ces_3_3_io_outs_up[11] ,
    \ces_3_3_io_outs_up[10] ,
    \ces_3_3_io_outs_up[9] ,
    \ces_3_3_io_outs_up[8] ,
    \ces_3_3_io_outs_up[7] ,
    \ces_3_3_io_outs_up[6] ,
    \ces_3_3_io_outs_up[5] ,
    \ces_3_3_io_outs_up[4] ,
    \ces_3_3_io_outs_up[3] ,
    \ces_3_3_io_outs_up[2] ,
    \ces_3_3_io_outs_up[1] ,
    \ces_3_3_io_outs_up[0] }));
 Element ces_3_4 (.clock(clknet_3_3_0_clock),
    .io_lsbIns_1(ces_3_3_io_lsbOuts_1),
    .io_lsbIns_2(ces_3_3_io_lsbOuts_2),
    .io_lsbIns_3(ces_3_3_io_lsbOuts_3),
    .io_lsbIns_4(ces_3_3_io_lsbOuts_4),
    .io_lsbIns_5(ces_3_3_io_lsbOuts_5),
    .io_lsbIns_6(ces_3_3_io_lsbOuts_6),
    .io_lsbIns_7(ces_3_3_io_lsbOuts_7),
    .io_lsbOuts_0(ces_3_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_4_io_lsbOuts_7),
    .io_ins_down({\ces_3_4_io_ins_down[63] ,
    \ces_3_4_io_ins_down[62] ,
    \ces_3_4_io_ins_down[61] ,
    \ces_3_4_io_ins_down[60] ,
    \ces_3_4_io_ins_down[59] ,
    \ces_3_4_io_ins_down[58] ,
    \ces_3_4_io_ins_down[57] ,
    \ces_3_4_io_ins_down[56] ,
    \ces_3_4_io_ins_down[55] ,
    \ces_3_4_io_ins_down[54] ,
    \ces_3_4_io_ins_down[53] ,
    \ces_3_4_io_ins_down[52] ,
    \ces_3_4_io_ins_down[51] ,
    \ces_3_4_io_ins_down[50] ,
    \ces_3_4_io_ins_down[49] ,
    \ces_3_4_io_ins_down[48] ,
    \ces_3_4_io_ins_down[47] ,
    \ces_3_4_io_ins_down[46] ,
    \ces_3_4_io_ins_down[45] ,
    \ces_3_4_io_ins_down[44] ,
    \ces_3_4_io_ins_down[43] ,
    \ces_3_4_io_ins_down[42] ,
    \ces_3_4_io_ins_down[41] ,
    \ces_3_4_io_ins_down[40] ,
    \ces_3_4_io_ins_down[39] ,
    \ces_3_4_io_ins_down[38] ,
    \ces_3_4_io_ins_down[37] ,
    \ces_3_4_io_ins_down[36] ,
    \ces_3_4_io_ins_down[35] ,
    \ces_3_4_io_ins_down[34] ,
    \ces_3_4_io_ins_down[33] ,
    \ces_3_4_io_ins_down[32] ,
    \ces_3_4_io_ins_down[31] ,
    \ces_3_4_io_ins_down[30] ,
    \ces_3_4_io_ins_down[29] ,
    \ces_3_4_io_ins_down[28] ,
    \ces_3_4_io_ins_down[27] ,
    \ces_3_4_io_ins_down[26] ,
    \ces_3_4_io_ins_down[25] ,
    \ces_3_4_io_ins_down[24] ,
    \ces_3_4_io_ins_down[23] ,
    \ces_3_4_io_ins_down[22] ,
    \ces_3_4_io_ins_down[21] ,
    \ces_3_4_io_ins_down[20] ,
    \ces_3_4_io_ins_down[19] ,
    \ces_3_4_io_ins_down[18] ,
    \ces_3_4_io_ins_down[17] ,
    \ces_3_4_io_ins_down[16] ,
    \ces_3_4_io_ins_down[15] ,
    \ces_3_4_io_ins_down[14] ,
    \ces_3_4_io_ins_down[13] ,
    \ces_3_4_io_ins_down[12] ,
    \ces_3_4_io_ins_down[11] ,
    \ces_3_4_io_ins_down[10] ,
    \ces_3_4_io_ins_down[9] ,
    \ces_3_4_io_ins_down[8] ,
    \ces_3_4_io_ins_down[7] ,
    \ces_3_4_io_ins_down[6] ,
    \ces_3_4_io_ins_down[5] ,
    \ces_3_4_io_ins_down[4] ,
    \ces_3_4_io_ins_down[3] ,
    \ces_3_4_io_ins_down[2] ,
    \ces_3_4_io_ins_down[1] ,
    \ces_3_4_io_ins_down[0] }),
    .io_ins_left({\ces_3_4_io_ins_left[63] ,
    \ces_3_4_io_ins_left[62] ,
    \ces_3_4_io_ins_left[61] ,
    \ces_3_4_io_ins_left[60] ,
    \ces_3_4_io_ins_left[59] ,
    \ces_3_4_io_ins_left[58] ,
    \ces_3_4_io_ins_left[57] ,
    \ces_3_4_io_ins_left[56] ,
    \ces_3_4_io_ins_left[55] ,
    \ces_3_4_io_ins_left[54] ,
    \ces_3_4_io_ins_left[53] ,
    \ces_3_4_io_ins_left[52] ,
    \ces_3_4_io_ins_left[51] ,
    \ces_3_4_io_ins_left[50] ,
    \ces_3_4_io_ins_left[49] ,
    \ces_3_4_io_ins_left[48] ,
    \ces_3_4_io_ins_left[47] ,
    \ces_3_4_io_ins_left[46] ,
    \ces_3_4_io_ins_left[45] ,
    \ces_3_4_io_ins_left[44] ,
    \ces_3_4_io_ins_left[43] ,
    \ces_3_4_io_ins_left[42] ,
    \ces_3_4_io_ins_left[41] ,
    \ces_3_4_io_ins_left[40] ,
    \ces_3_4_io_ins_left[39] ,
    \ces_3_4_io_ins_left[38] ,
    \ces_3_4_io_ins_left[37] ,
    \ces_3_4_io_ins_left[36] ,
    \ces_3_4_io_ins_left[35] ,
    \ces_3_4_io_ins_left[34] ,
    \ces_3_4_io_ins_left[33] ,
    \ces_3_4_io_ins_left[32] ,
    \ces_3_4_io_ins_left[31] ,
    \ces_3_4_io_ins_left[30] ,
    \ces_3_4_io_ins_left[29] ,
    \ces_3_4_io_ins_left[28] ,
    \ces_3_4_io_ins_left[27] ,
    \ces_3_4_io_ins_left[26] ,
    \ces_3_4_io_ins_left[25] ,
    \ces_3_4_io_ins_left[24] ,
    \ces_3_4_io_ins_left[23] ,
    \ces_3_4_io_ins_left[22] ,
    \ces_3_4_io_ins_left[21] ,
    \ces_3_4_io_ins_left[20] ,
    \ces_3_4_io_ins_left[19] ,
    \ces_3_4_io_ins_left[18] ,
    \ces_3_4_io_ins_left[17] ,
    \ces_3_4_io_ins_left[16] ,
    \ces_3_4_io_ins_left[15] ,
    \ces_3_4_io_ins_left[14] ,
    \ces_3_4_io_ins_left[13] ,
    \ces_3_4_io_ins_left[12] ,
    \ces_3_4_io_ins_left[11] ,
    \ces_3_4_io_ins_left[10] ,
    \ces_3_4_io_ins_left[9] ,
    \ces_3_4_io_ins_left[8] ,
    \ces_3_4_io_ins_left[7] ,
    \ces_3_4_io_ins_left[6] ,
    \ces_3_4_io_ins_left[5] ,
    \ces_3_4_io_ins_left[4] ,
    \ces_3_4_io_ins_left[3] ,
    \ces_3_4_io_ins_left[2] ,
    \ces_3_4_io_ins_left[1] ,
    \ces_3_4_io_ins_left[0] }),
    .io_ins_right({\ces_3_3_io_outs_right[63] ,
    \ces_3_3_io_outs_right[62] ,
    \ces_3_3_io_outs_right[61] ,
    \ces_3_3_io_outs_right[60] ,
    \ces_3_3_io_outs_right[59] ,
    \ces_3_3_io_outs_right[58] ,
    \ces_3_3_io_outs_right[57] ,
    \ces_3_3_io_outs_right[56] ,
    \ces_3_3_io_outs_right[55] ,
    \ces_3_3_io_outs_right[54] ,
    \ces_3_3_io_outs_right[53] ,
    \ces_3_3_io_outs_right[52] ,
    \ces_3_3_io_outs_right[51] ,
    \ces_3_3_io_outs_right[50] ,
    \ces_3_3_io_outs_right[49] ,
    \ces_3_3_io_outs_right[48] ,
    \ces_3_3_io_outs_right[47] ,
    \ces_3_3_io_outs_right[46] ,
    \ces_3_3_io_outs_right[45] ,
    \ces_3_3_io_outs_right[44] ,
    \ces_3_3_io_outs_right[43] ,
    \ces_3_3_io_outs_right[42] ,
    \ces_3_3_io_outs_right[41] ,
    \ces_3_3_io_outs_right[40] ,
    \ces_3_3_io_outs_right[39] ,
    \ces_3_3_io_outs_right[38] ,
    \ces_3_3_io_outs_right[37] ,
    \ces_3_3_io_outs_right[36] ,
    \ces_3_3_io_outs_right[35] ,
    \ces_3_3_io_outs_right[34] ,
    \ces_3_3_io_outs_right[33] ,
    \ces_3_3_io_outs_right[32] ,
    \ces_3_3_io_outs_right[31] ,
    \ces_3_3_io_outs_right[30] ,
    \ces_3_3_io_outs_right[29] ,
    \ces_3_3_io_outs_right[28] ,
    \ces_3_3_io_outs_right[27] ,
    \ces_3_3_io_outs_right[26] ,
    \ces_3_3_io_outs_right[25] ,
    \ces_3_3_io_outs_right[24] ,
    \ces_3_3_io_outs_right[23] ,
    \ces_3_3_io_outs_right[22] ,
    \ces_3_3_io_outs_right[21] ,
    \ces_3_3_io_outs_right[20] ,
    \ces_3_3_io_outs_right[19] ,
    \ces_3_3_io_outs_right[18] ,
    \ces_3_3_io_outs_right[17] ,
    \ces_3_3_io_outs_right[16] ,
    \ces_3_3_io_outs_right[15] ,
    \ces_3_3_io_outs_right[14] ,
    \ces_3_3_io_outs_right[13] ,
    \ces_3_3_io_outs_right[12] ,
    \ces_3_3_io_outs_right[11] ,
    \ces_3_3_io_outs_right[10] ,
    \ces_3_3_io_outs_right[9] ,
    \ces_3_3_io_outs_right[8] ,
    \ces_3_3_io_outs_right[7] ,
    \ces_3_3_io_outs_right[6] ,
    \ces_3_3_io_outs_right[5] ,
    \ces_3_3_io_outs_right[4] ,
    \ces_3_3_io_outs_right[3] ,
    \ces_3_3_io_outs_right[2] ,
    \ces_3_3_io_outs_right[1] ,
    \ces_3_3_io_outs_right[0] }),
    .io_ins_up({\ces_2_4_io_outs_up[63] ,
    \ces_2_4_io_outs_up[62] ,
    \ces_2_4_io_outs_up[61] ,
    \ces_2_4_io_outs_up[60] ,
    \ces_2_4_io_outs_up[59] ,
    \ces_2_4_io_outs_up[58] ,
    \ces_2_4_io_outs_up[57] ,
    \ces_2_4_io_outs_up[56] ,
    \ces_2_4_io_outs_up[55] ,
    \ces_2_4_io_outs_up[54] ,
    \ces_2_4_io_outs_up[53] ,
    \ces_2_4_io_outs_up[52] ,
    \ces_2_4_io_outs_up[51] ,
    \ces_2_4_io_outs_up[50] ,
    \ces_2_4_io_outs_up[49] ,
    \ces_2_4_io_outs_up[48] ,
    \ces_2_4_io_outs_up[47] ,
    \ces_2_4_io_outs_up[46] ,
    \ces_2_4_io_outs_up[45] ,
    \ces_2_4_io_outs_up[44] ,
    \ces_2_4_io_outs_up[43] ,
    \ces_2_4_io_outs_up[42] ,
    \ces_2_4_io_outs_up[41] ,
    \ces_2_4_io_outs_up[40] ,
    \ces_2_4_io_outs_up[39] ,
    \ces_2_4_io_outs_up[38] ,
    \ces_2_4_io_outs_up[37] ,
    \ces_2_4_io_outs_up[36] ,
    \ces_2_4_io_outs_up[35] ,
    \ces_2_4_io_outs_up[34] ,
    \ces_2_4_io_outs_up[33] ,
    \ces_2_4_io_outs_up[32] ,
    \ces_2_4_io_outs_up[31] ,
    \ces_2_4_io_outs_up[30] ,
    \ces_2_4_io_outs_up[29] ,
    \ces_2_4_io_outs_up[28] ,
    \ces_2_4_io_outs_up[27] ,
    \ces_2_4_io_outs_up[26] ,
    \ces_2_4_io_outs_up[25] ,
    \ces_2_4_io_outs_up[24] ,
    \ces_2_4_io_outs_up[23] ,
    \ces_2_4_io_outs_up[22] ,
    \ces_2_4_io_outs_up[21] ,
    \ces_2_4_io_outs_up[20] ,
    \ces_2_4_io_outs_up[19] ,
    \ces_2_4_io_outs_up[18] ,
    \ces_2_4_io_outs_up[17] ,
    \ces_2_4_io_outs_up[16] ,
    \ces_2_4_io_outs_up[15] ,
    \ces_2_4_io_outs_up[14] ,
    \ces_2_4_io_outs_up[13] ,
    \ces_2_4_io_outs_up[12] ,
    \ces_2_4_io_outs_up[11] ,
    \ces_2_4_io_outs_up[10] ,
    \ces_2_4_io_outs_up[9] ,
    \ces_2_4_io_outs_up[8] ,
    \ces_2_4_io_outs_up[7] ,
    \ces_2_4_io_outs_up[6] ,
    \ces_2_4_io_outs_up[5] ,
    \ces_2_4_io_outs_up[4] ,
    \ces_2_4_io_outs_up[3] ,
    \ces_2_4_io_outs_up[2] ,
    \ces_2_4_io_outs_up[1] ,
    \ces_2_4_io_outs_up[0] }),
    .io_outs_down({\ces_2_4_io_ins_down[63] ,
    \ces_2_4_io_ins_down[62] ,
    \ces_2_4_io_ins_down[61] ,
    \ces_2_4_io_ins_down[60] ,
    \ces_2_4_io_ins_down[59] ,
    \ces_2_4_io_ins_down[58] ,
    \ces_2_4_io_ins_down[57] ,
    \ces_2_4_io_ins_down[56] ,
    \ces_2_4_io_ins_down[55] ,
    \ces_2_4_io_ins_down[54] ,
    \ces_2_4_io_ins_down[53] ,
    \ces_2_4_io_ins_down[52] ,
    \ces_2_4_io_ins_down[51] ,
    \ces_2_4_io_ins_down[50] ,
    \ces_2_4_io_ins_down[49] ,
    \ces_2_4_io_ins_down[48] ,
    \ces_2_4_io_ins_down[47] ,
    \ces_2_4_io_ins_down[46] ,
    \ces_2_4_io_ins_down[45] ,
    \ces_2_4_io_ins_down[44] ,
    \ces_2_4_io_ins_down[43] ,
    \ces_2_4_io_ins_down[42] ,
    \ces_2_4_io_ins_down[41] ,
    \ces_2_4_io_ins_down[40] ,
    \ces_2_4_io_ins_down[39] ,
    \ces_2_4_io_ins_down[38] ,
    \ces_2_4_io_ins_down[37] ,
    \ces_2_4_io_ins_down[36] ,
    \ces_2_4_io_ins_down[35] ,
    \ces_2_4_io_ins_down[34] ,
    \ces_2_4_io_ins_down[33] ,
    \ces_2_4_io_ins_down[32] ,
    \ces_2_4_io_ins_down[31] ,
    \ces_2_4_io_ins_down[30] ,
    \ces_2_4_io_ins_down[29] ,
    \ces_2_4_io_ins_down[28] ,
    \ces_2_4_io_ins_down[27] ,
    \ces_2_4_io_ins_down[26] ,
    \ces_2_4_io_ins_down[25] ,
    \ces_2_4_io_ins_down[24] ,
    \ces_2_4_io_ins_down[23] ,
    \ces_2_4_io_ins_down[22] ,
    \ces_2_4_io_ins_down[21] ,
    \ces_2_4_io_ins_down[20] ,
    \ces_2_4_io_ins_down[19] ,
    \ces_2_4_io_ins_down[18] ,
    \ces_2_4_io_ins_down[17] ,
    \ces_2_4_io_ins_down[16] ,
    \ces_2_4_io_ins_down[15] ,
    \ces_2_4_io_ins_down[14] ,
    \ces_2_4_io_ins_down[13] ,
    \ces_2_4_io_ins_down[12] ,
    \ces_2_4_io_ins_down[11] ,
    \ces_2_4_io_ins_down[10] ,
    \ces_2_4_io_ins_down[9] ,
    \ces_2_4_io_ins_down[8] ,
    \ces_2_4_io_ins_down[7] ,
    \ces_2_4_io_ins_down[6] ,
    \ces_2_4_io_ins_down[5] ,
    \ces_2_4_io_ins_down[4] ,
    \ces_2_4_io_ins_down[3] ,
    \ces_2_4_io_ins_down[2] ,
    \ces_2_4_io_ins_down[1] ,
    \ces_2_4_io_ins_down[0] }),
    .io_outs_left({\ces_3_3_io_ins_left[63] ,
    \ces_3_3_io_ins_left[62] ,
    \ces_3_3_io_ins_left[61] ,
    \ces_3_3_io_ins_left[60] ,
    \ces_3_3_io_ins_left[59] ,
    \ces_3_3_io_ins_left[58] ,
    \ces_3_3_io_ins_left[57] ,
    \ces_3_3_io_ins_left[56] ,
    \ces_3_3_io_ins_left[55] ,
    \ces_3_3_io_ins_left[54] ,
    \ces_3_3_io_ins_left[53] ,
    \ces_3_3_io_ins_left[52] ,
    \ces_3_3_io_ins_left[51] ,
    \ces_3_3_io_ins_left[50] ,
    \ces_3_3_io_ins_left[49] ,
    \ces_3_3_io_ins_left[48] ,
    \ces_3_3_io_ins_left[47] ,
    \ces_3_3_io_ins_left[46] ,
    \ces_3_3_io_ins_left[45] ,
    \ces_3_3_io_ins_left[44] ,
    \ces_3_3_io_ins_left[43] ,
    \ces_3_3_io_ins_left[42] ,
    \ces_3_3_io_ins_left[41] ,
    \ces_3_3_io_ins_left[40] ,
    \ces_3_3_io_ins_left[39] ,
    \ces_3_3_io_ins_left[38] ,
    \ces_3_3_io_ins_left[37] ,
    \ces_3_3_io_ins_left[36] ,
    \ces_3_3_io_ins_left[35] ,
    \ces_3_3_io_ins_left[34] ,
    \ces_3_3_io_ins_left[33] ,
    \ces_3_3_io_ins_left[32] ,
    \ces_3_3_io_ins_left[31] ,
    \ces_3_3_io_ins_left[30] ,
    \ces_3_3_io_ins_left[29] ,
    \ces_3_3_io_ins_left[28] ,
    \ces_3_3_io_ins_left[27] ,
    \ces_3_3_io_ins_left[26] ,
    \ces_3_3_io_ins_left[25] ,
    \ces_3_3_io_ins_left[24] ,
    \ces_3_3_io_ins_left[23] ,
    \ces_3_3_io_ins_left[22] ,
    \ces_3_3_io_ins_left[21] ,
    \ces_3_3_io_ins_left[20] ,
    \ces_3_3_io_ins_left[19] ,
    \ces_3_3_io_ins_left[18] ,
    \ces_3_3_io_ins_left[17] ,
    \ces_3_3_io_ins_left[16] ,
    \ces_3_3_io_ins_left[15] ,
    \ces_3_3_io_ins_left[14] ,
    \ces_3_3_io_ins_left[13] ,
    \ces_3_3_io_ins_left[12] ,
    \ces_3_3_io_ins_left[11] ,
    \ces_3_3_io_ins_left[10] ,
    \ces_3_3_io_ins_left[9] ,
    \ces_3_3_io_ins_left[8] ,
    \ces_3_3_io_ins_left[7] ,
    \ces_3_3_io_ins_left[6] ,
    \ces_3_3_io_ins_left[5] ,
    \ces_3_3_io_ins_left[4] ,
    \ces_3_3_io_ins_left[3] ,
    \ces_3_3_io_ins_left[2] ,
    \ces_3_3_io_ins_left[1] ,
    \ces_3_3_io_ins_left[0] }),
    .io_outs_right({\ces_3_4_io_outs_right[63] ,
    \ces_3_4_io_outs_right[62] ,
    \ces_3_4_io_outs_right[61] ,
    \ces_3_4_io_outs_right[60] ,
    \ces_3_4_io_outs_right[59] ,
    \ces_3_4_io_outs_right[58] ,
    \ces_3_4_io_outs_right[57] ,
    \ces_3_4_io_outs_right[56] ,
    \ces_3_4_io_outs_right[55] ,
    \ces_3_4_io_outs_right[54] ,
    \ces_3_4_io_outs_right[53] ,
    \ces_3_4_io_outs_right[52] ,
    \ces_3_4_io_outs_right[51] ,
    \ces_3_4_io_outs_right[50] ,
    \ces_3_4_io_outs_right[49] ,
    \ces_3_4_io_outs_right[48] ,
    \ces_3_4_io_outs_right[47] ,
    \ces_3_4_io_outs_right[46] ,
    \ces_3_4_io_outs_right[45] ,
    \ces_3_4_io_outs_right[44] ,
    \ces_3_4_io_outs_right[43] ,
    \ces_3_4_io_outs_right[42] ,
    \ces_3_4_io_outs_right[41] ,
    \ces_3_4_io_outs_right[40] ,
    \ces_3_4_io_outs_right[39] ,
    \ces_3_4_io_outs_right[38] ,
    \ces_3_4_io_outs_right[37] ,
    \ces_3_4_io_outs_right[36] ,
    \ces_3_4_io_outs_right[35] ,
    \ces_3_4_io_outs_right[34] ,
    \ces_3_4_io_outs_right[33] ,
    \ces_3_4_io_outs_right[32] ,
    \ces_3_4_io_outs_right[31] ,
    \ces_3_4_io_outs_right[30] ,
    \ces_3_4_io_outs_right[29] ,
    \ces_3_4_io_outs_right[28] ,
    \ces_3_4_io_outs_right[27] ,
    \ces_3_4_io_outs_right[26] ,
    \ces_3_4_io_outs_right[25] ,
    \ces_3_4_io_outs_right[24] ,
    \ces_3_4_io_outs_right[23] ,
    \ces_3_4_io_outs_right[22] ,
    \ces_3_4_io_outs_right[21] ,
    \ces_3_4_io_outs_right[20] ,
    \ces_3_4_io_outs_right[19] ,
    \ces_3_4_io_outs_right[18] ,
    \ces_3_4_io_outs_right[17] ,
    \ces_3_4_io_outs_right[16] ,
    \ces_3_4_io_outs_right[15] ,
    \ces_3_4_io_outs_right[14] ,
    \ces_3_4_io_outs_right[13] ,
    \ces_3_4_io_outs_right[12] ,
    \ces_3_4_io_outs_right[11] ,
    \ces_3_4_io_outs_right[10] ,
    \ces_3_4_io_outs_right[9] ,
    \ces_3_4_io_outs_right[8] ,
    \ces_3_4_io_outs_right[7] ,
    \ces_3_4_io_outs_right[6] ,
    \ces_3_4_io_outs_right[5] ,
    \ces_3_4_io_outs_right[4] ,
    \ces_3_4_io_outs_right[3] ,
    \ces_3_4_io_outs_right[2] ,
    \ces_3_4_io_outs_right[1] ,
    \ces_3_4_io_outs_right[0] }),
    .io_outs_up({\ces_3_4_io_outs_up[63] ,
    \ces_3_4_io_outs_up[62] ,
    \ces_3_4_io_outs_up[61] ,
    \ces_3_4_io_outs_up[60] ,
    \ces_3_4_io_outs_up[59] ,
    \ces_3_4_io_outs_up[58] ,
    \ces_3_4_io_outs_up[57] ,
    \ces_3_4_io_outs_up[56] ,
    \ces_3_4_io_outs_up[55] ,
    \ces_3_4_io_outs_up[54] ,
    \ces_3_4_io_outs_up[53] ,
    \ces_3_4_io_outs_up[52] ,
    \ces_3_4_io_outs_up[51] ,
    \ces_3_4_io_outs_up[50] ,
    \ces_3_4_io_outs_up[49] ,
    \ces_3_4_io_outs_up[48] ,
    \ces_3_4_io_outs_up[47] ,
    \ces_3_4_io_outs_up[46] ,
    \ces_3_4_io_outs_up[45] ,
    \ces_3_4_io_outs_up[44] ,
    \ces_3_4_io_outs_up[43] ,
    \ces_3_4_io_outs_up[42] ,
    \ces_3_4_io_outs_up[41] ,
    \ces_3_4_io_outs_up[40] ,
    \ces_3_4_io_outs_up[39] ,
    \ces_3_4_io_outs_up[38] ,
    \ces_3_4_io_outs_up[37] ,
    \ces_3_4_io_outs_up[36] ,
    \ces_3_4_io_outs_up[35] ,
    \ces_3_4_io_outs_up[34] ,
    \ces_3_4_io_outs_up[33] ,
    \ces_3_4_io_outs_up[32] ,
    \ces_3_4_io_outs_up[31] ,
    \ces_3_4_io_outs_up[30] ,
    \ces_3_4_io_outs_up[29] ,
    \ces_3_4_io_outs_up[28] ,
    \ces_3_4_io_outs_up[27] ,
    \ces_3_4_io_outs_up[26] ,
    \ces_3_4_io_outs_up[25] ,
    \ces_3_4_io_outs_up[24] ,
    \ces_3_4_io_outs_up[23] ,
    \ces_3_4_io_outs_up[22] ,
    \ces_3_4_io_outs_up[21] ,
    \ces_3_4_io_outs_up[20] ,
    \ces_3_4_io_outs_up[19] ,
    \ces_3_4_io_outs_up[18] ,
    \ces_3_4_io_outs_up[17] ,
    \ces_3_4_io_outs_up[16] ,
    \ces_3_4_io_outs_up[15] ,
    \ces_3_4_io_outs_up[14] ,
    \ces_3_4_io_outs_up[13] ,
    \ces_3_4_io_outs_up[12] ,
    \ces_3_4_io_outs_up[11] ,
    \ces_3_4_io_outs_up[10] ,
    \ces_3_4_io_outs_up[9] ,
    \ces_3_4_io_outs_up[8] ,
    \ces_3_4_io_outs_up[7] ,
    \ces_3_4_io_outs_up[6] ,
    \ces_3_4_io_outs_up[5] ,
    \ces_3_4_io_outs_up[4] ,
    \ces_3_4_io_outs_up[3] ,
    \ces_3_4_io_outs_up[2] ,
    \ces_3_4_io_outs_up[1] ,
    \ces_3_4_io_outs_up[0] }));
 Element ces_3_5 (.clock(clknet_3_3_0_clock),
    .io_lsbIns_1(ces_3_4_io_lsbOuts_1),
    .io_lsbIns_2(ces_3_4_io_lsbOuts_2),
    .io_lsbIns_3(ces_3_4_io_lsbOuts_3),
    .io_lsbIns_4(ces_3_4_io_lsbOuts_4),
    .io_lsbIns_5(ces_3_4_io_lsbOuts_5),
    .io_lsbIns_6(ces_3_4_io_lsbOuts_6),
    .io_lsbIns_7(ces_3_4_io_lsbOuts_7),
    .io_lsbOuts_0(ces_3_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_5_io_lsbOuts_7),
    .io_ins_down({\ces_3_5_io_ins_down[63] ,
    \ces_3_5_io_ins_down[62] ,
    \ces_3_5_io_ins_down[61] ,
    \ces_3_5_io_ins_down[60] ,
    \ces_3_5_io_ins_down[59] ,
    \ces_3_5_io_ins_down[58] ,
    \ces_3_5_io_ins_down[57] ,
    \ces_3_5_io_ins_down[56] ,
    \ces_3_5_io_ins_down[55] ,
    \ces_3_5_io_ins_down[54] ,
    \ces_3_5_io_ins_down[53] ,
    \ces_3_5_io_ins_down[52] ,
    \ces_3_5_io_ins_down[51] ,
    \ces_3_5_io_ins_down[50] ,
    \ces_3_5_io_ins_down[49] ,
    \ces_3_5_io_ins_down[48] ,
    \ces_3_5_io_ins_down[47] ,
    \ces_3_5_io_ins_down[46] ,
    \ces_3_5_io_ins_down[45] ,
    \ces_3_5_io_ins_down[44] ,
    \ces_3_5_io_ins_down[43] ,
    \ces_3_5_io_ins_down[42] ,
    \ces_3_5_io_ins_down[41] ,
    \ces_3_5_io_ins_down[40] ,
    \ces_3_5_io_ins_down[39] ,
    \ces_3_5_io_ins_down[38] ,
    \ces_3_5_io_ins_down[37] ,
    \ces_3_5_io_ins_down[36] ,
    \ces_3_5_io_ins_down[35] ,
    \ces_3_5_io_ins_down[34] ,
    \ces_3_5_io_ins_down[33] ,
    \ces_3_5_io_ins_down[32] ,
    \ces_3_5_io_ins_down[31] ,
    \ces_3_5_io_ins_down[30] ,
    \ces_3_5_io_ins_down[29] ,
    \ces_3_5_io_ins_down[28] ,
    \ces_3_5_io_ins_down[27] ,
    \ces_3_5_io_ins_down[26] ,
    \ces_3_5_io_ins_down[25] ,
    \ces_3_5_io_ins_down[24] ,
    \ces_3_5_io_ins_down[23] ,
    \ces_3_5_io_ins_down[22] ,
    \ces_3_5_io_ins_down[21] ,
    \ces_3_5_io_ins_down[20] ,
    \ces_3_5_io_ins_down[19] ,
    \ces_3_5_io_ins_down[18] ,
    \ces_3_5_io_ins_down[17] ,
    \ces_3_5_io_ins_down[16] ,
    \ces_3_5_io_ins_down[15] ,
    \ces_3_5_io_ins_down[14] ,
    \ces_3_5_io_ins_down[13] ,
    \ces_3_5_io_ins_down[12] ,
    \ces_3_5_io_ins_down[11] ,
    \ces_3_5_io_ins_down[10] ,
    \ces_3_5_io_ins_down[9] ,
    \ces_3_5_io_ins_down[8] ,
    \ces_3_5_io_ins_down[7] ,
    \ces_3_5_io_ins_down[6] ,
    \ces_3_5_io_ins_down[5] ,
    \ces_3_5_io_ins_down[4] ,
    \ces_3_5_io_ins_down[3] ,
    \ces_3_5_io_ins_down[2] ,
    \ces_3_5_io_ins_down[1] ,
    \ces_3_5_io_ins_down[0] }),
    .io_ins_left({\ces_3_5_io_ins_left[63] ,
    \ces_3_5_io_ins_left[62] ,
    \ces_3_5_io_ins_left[61] ,
    \ces_3_5_io_ins_left[60] ,
    \ces_3_5_io_ins_left[59] ,
    \ces_3_5_io_ins_left[58] ,
    \ces_3_5_io_ins_left[57] ,
    \ces_3_5_io_ins_left[56] ,
    \ces_3_5_io_ins_left[55] ,
    \ces_3_5_io_ins_left[54] ,
    \ces_3_5_io_ins_left[53] ,
    \ces_3_5_io_ins_left[52] ,
    \ces_3_5_io_ins_left[51] ,
    \ces_3_5_io_ins_left[50] ,
    \ces_3_5_io_ins_left[49] ,
    \ces_3_5_io_ins_left[48] ,
    \ces_3_5_io_ins_left[47] ,
    \ces_3_5_io_ins_left[46] ,
    \ces_3_5_io_ins_left[45] ,
    \ces_3_5_io_ins_left[44] ,
    \ces_3_5_io_ins_left[43] ,
    \ces_3_5_io_ins_left[42] ,
    \ces_3_5_io_ins_left[41] ,
    \ces_3_5_io_ins_left[40] ,
    \ces_3_5_io_ins_left[39] ,
    \ces_3_5_io_ins_left[38] ,
    \ces_3_5_io_ins_left[37] ,
    \ces_3_5_io_ins_left[36] ,
    \ces_3_5_io_ins_left[35] ,
    \ces_3_5_io_ins_left[34] ,
    \ces_3_5_io_ins_left[33] ,
    \ces_3_5_io_ins_left[32] ,
    \ces_3_5_io_ins_left[31] ,
    \ces_3_5_io_ins_left[30] ,
    \ces_3_5_io_ins_left[29] ,
    \ces_3_5_io_ins_left[28] ,
    \ces_3_5_io_ins_left[27] ,
    \ces_3_5_io_ins_left[26] ,
    \ces_3_5_io_ins_left[25] ,
    \ces_3_5_io_ins_left[24] ,
    \ces_3_5_io_ins_left[23] ,
    \ces_3_5_io_ins_left[22] ,
    \ces_3_5_io_ins_left[21] ,
    \ces_3_5_io_ins_left[20] ,
    \ces_3_5_io_ins_left[19] ,
    \ces_3_5_io_ins_left[18] ,
    \ces_3_5_io_ins_left[17] ,
    \ces_3_5_io_ins_left[16] ,
    \ces_3_5_io_ins_left[15] ,
    \ces_3_5_io_ins_left[14] ,
    \ces_3_5_io_ins_left[13] ,
    \ces_3_5_io_ins_left[12] ,
    \ces_3_5_io_ins_left[11] ,
    \ces_3_5_io_ins_left[10] ,
    \ces_3_5_io_ins_left[9] ,
    \ces_3_5_io_ins_left[8] ,
    \ces_3_5_io_ins_left[7] ,
    \ces_3_5_io_ins_left[6] ,
    \ces_3_5_io_ins_left[5] ,
    \ces_3_5_io_ins_left[4] ,
    \ces_3_5_io_ins_left[3] ,
    \ces_3_5_io_ins_left[2] ,
    \ces_3_5_io_ins_left[1] ,
    \ces_3_5_io_ins_left[0] }),
    .io_ins_right({\ces_3_4_io_outs_right[63] ,
    \ces_3_4_io_outs_right[62] ,
    \ces_3_4_io_outs_right[61] ,
    \ces_3_4_io_outs_right[60] ,
    \ces_3_4_io_outs_right[59] ,
    \ces_3_4_io_outs_right[58] ,
    \ces_3_4_io_outs_right[57] ,
    \ces_3_4_io_outs_right[56] ,
    \ces_3_4_io_outs_right[55] ,
    \ces_3_4_io_outs_right[54] ,
    \ces_3_4_io_outs_right[53] ,
    \ces_3_4_io_outs_right[52] ,
    \ces_3_4_io_outs_right[51] ,
    \ces_3_4_io_outs_right[50] ,
    \ces_3_4_io_outs_right[49] ,
    \ces_3_4_io_outs_right[48] ,
    \ces_3_4_io_outs_right[47] ,
    \ces_3_4_io_outs_right[46] ,
    \ces_3_4_io_outs_right[45] ,
    \ces_3_4_io_outs_right[44] ,
    \ces_3_4_io_outs_right[43] ,
    \ces_3_4_io_outs_right[42] ,
    \ces_3_4_io_outs_right[41] ,
    \ces_3_4_io_outs_right[40] ,
    \ces_3_4_io_outs_right[39] ,
    \ces_3_4_io_outs_right[38] ,
    \ces_3_4_io_outs_right[37] ,
    \ces_3_4_io_outs_right[36] ,
    \ces_3_4_io_outs_right[35] ,
    \ces_3_4_io_outs_right[34] ,
    \ces_3_4_io_outs_right[33] ,
    \ces_3_4_io_outs_right[32] ,
    \ces_3_4_io_outs_right[31] ,
    \ces_3_4_io_outs_right[30] ,
    \ces_3_4_io_outs_right[29] ,
    \ces_3_4_io_outs_right[28] ,
    \ces_3_4_io_outs_right[27] ,
    \ces_3_4_io_outs_right[26] ,
    \ces_3_4_io_outs_right[25] ,
    \ces_3_4_io_outs_right[24] ,
    \ces_3_4_io_outs_right[23] ,
    \ces_3_4_io_outs_right[22] ,
    \ces_3_4_io_outs_right[21] ,
    \ces_3_4_io_outs_right[20] ,
    \ces_3_4_io_outs_right[19] ,
    \ces_3_4_io_outs_right[18] ,
    \ces_3_4_io_outs_right[17] ,
    \ces_3_4_io_outs_right[16] ,
    \ces_3_4_io_outs_right[15] ,
    \ces_3_4_io_outs_right[14] ,
    \ces_3_4_io_outs_right[13] ,
    \ces_3_4_io_outs_right[12] ,
    \ces_3_4_io_outs_right[11] ,
    \ces_3_4_io_outs_right[10] ,
    \ces_3_4_io_outs_right[9] ,
    \ces_3_4_io_outs_right[8] ,
    \ces_3_4_io_outs_right[7] ,
    \ces_3_4_io_outs_right[6] ,
    \ces_3_4_io_outs_right[5] ,
    \ces_3_4_io_outs_right[4] ,
    \ces_3_4_io_outs_right[3] ,
    \ces_3_4_io_outs_right[2] ,
    \ces_3_4_io_outs_right[1] ,
    \ces_3_4_io_outs_right[0] }),
    .io_ins_up({\ces_2_5_io_outs_up[63] ,
    \ces_2_5_io_outs_up[62] ,
    \ces_2_5_io_outs_up[61] ,
    \ces_2_5_io_outs_up[60] ,
    \ces_2_5_io_outs_up[59] ,
    \ces_2_5_io_outs_up[58] ,
    \ces_2_5_io_outs_up[57] ,
    \ces_2_5_io_outs_up[56] ,
    \ces_2_5_io_outs_up[55] ,
    \ces_2_5_io_outs_up[54] ,
    \ces_2_5_io_outs_up[53] ,
    \ces_2_5_io_outs_up[52] ,
    \ces_2_5_io_outs_up[51] ,
    \ces_2_5_io_outs_up[50] ,
    \ces_2_5_io_outs_up[49] ,
    \ces_2_5_io_outs_up[48] ,
    \ces_2_5_io_outs_up[47] ,
    \ces_2_5_io_outs_up[46] ,
    \ces_2_5_io_outs_up[45] ,
    \ces_2_5_io_outs_up[44] ,
    \ces_2_5_io_outs_up[43] ,
    \ces_2_5_io_outs_up[42] ,
    \ces_2_5_io_outs_up[41] ,
    \ces_2_5_io_outs_up[40] ,
    \ces_2_5_io_outs_up[39] ,
    \ces_2_5_io_outs_up[38] ,
    \ces_2_5_io_outs_up[37] ,
    \ces_2_5_io_outs_up[36] ,
    \ces_2_5_io_outs_up[35] ,
    \ces_2_5_io_outs_up[34] ,
    \ces_2_5_io_outs_up[33] ,
    \ces_2_5_io_outs_up[32] ,
    \ces_2_5_io_outs_up[31] ,
    \ces_2_5_io_outs_up[30] ,
    \ces_2_5_io_outs_up[29] ,
    \ces_2_5_io_outs_up[28] ,
    \ces_2_5_io_outs_up[27] ,
    \ces_2_5_io_outs_up[26] ,
    \ces_2_5_io_outs_up[25] ,
    \ces_2_5_io_outs_up[24] ,
    \ces_2_5_io_outs_up[23] ,
    \ces_2_5_io_outs_up[22] ,
    \ces_2_5_io_outs_up[21] ,
    \ces_2_5_io_outs_up[20] ,
    \ces_2_5_io_outs_up[19] ,
    \ces_2_5_io_outs_up[18] ,
    \ces_2_5_io_outs_up[17] ,
    \ces_2_5_io_outs_up[16] ,
    \ces_2_5_io_outs_up[15] ,
    \ces_2_5_io_outs_up[14] ,
    \ces_2_5_io_outs_up[13] ,
    \ces_2_5_io_outs_up[12] ,
    \ces_2_5_io_outs_up[11] ,
    \ces_2_5_io_outs_up[10] ,
    \ces_2_5_io_outs_up[9] ,
    \ces_2_5_io_outs_up[8] ,
    \ces_2_5_io_outs_up[7] ,
    \ces_2_5_io_outs_up[6] ,
    \ces_2_5_io_outs_up[5] ,
    \ces_2_5_io_outs_up[4] ,
    \ces_2_5_io_outs_up[3] ,
    \ces_2_5_io_outs_up[2] ,
    \ces_2_5_io_outs_up[1] ,
    \ces_2_5_io_outs_up[0] }),
    .io_outs_down({\ces_2_5_io_ins_down[63] ,
    \ces_2_5_io_ins_down[62] ,
    \ces_2_5_io_ins_down[61] ,
    \ces_2_5_io_ins_down[60] ,
    \ces_2_5_io_ins_down[59] ,
    \ces_2_5_io_ins_down[58] ,
    \ces_2_5_io_ins_down[57] ,
    \ces_2_5_io_ins_down[56] ,
    \ces_2_5_io_ins_down[55] ,
    \ces_2_5_io_ins_down[54] ,
    \ces_2_5_io_ins_down[53] ,
    \ces_2_5_io_ins_down[52] ,
    \ces_2_5_io_ins_down[51] ,
    \ces_2_5_io_ins_down[50] ,
    \ces_2_5_io_ins_down[49] ,
    \ces_2_5_io_ins_down[48] ,
    \ces_2_5_io_ins_down[47] ,
    \ces_2_5_io_ins_down[46] ,
    \ces_2_5_io_ins_down[45] ,
    \ces_2_5_io_ins_down[44] ,
    \ces_2_5_io_ins_down[43] ,
    \ces_2_5_io_ins_down[42] ,
    \ces_2_5_io_ins_down[41] ,
    \ces_2_5_io_ins_down[40] ,
    \ces_2_5_io_ins_down[39] ,
    \ces_2_5_io_ins_down[38] ,
    \ces_2_5_io_ins_down[37] ,
    \ces_2_5_io_ins_down[36] ,
    \ces_2_5_io_ins_down[35] ,
    \ces_2_5_io_ins_down[34] ,
    \ces_2_5_io_ins_down[33] ,
    \ces_2_5_io_ins_down[32] ,
    \ces_2_5_io_ins_down[31] ,
    \ces_2_5_io_ins_down[30] ,
    \ces_2_5_io_ins_down[29] ,
    \ces_2_5_io_ins_down[28] ,
    \ces_2_5_io_ins_down[27] ,
    \ces_2_5_io_ins_down[26] ,
    \ces_2_5_io_ins_down[25] ,
    \ces_2_5_io_ins_down[24] ,
    \ces_2_5_io_ins_down[23] ,
    \ces_2_5_io_ins_down[22] ,
    \ces_2_5_io_ins_down[21] ,
    \ces_2_5_io_ins_down[20] ,
    \ces_2_5_io_ins_down[19] ,
    \ces_2_5_io_ins_down[18] ,
    \ces_2_5_io_ins_down[17] ,
    \ces_2_5_io_ins_down[16] ,
    \ces_2_5_io_ins_down[15] ,
    \ces_2_5_io_ins_down[14] ,
    \ces_2_5_io_ins_down[13] ,
    \ces_2_5_io_ins_down[12] ,
    \ces_2_5_io_ins_down[11] ,
    \ces_2_5_io_ins_down[10] ,
    \ces_2_5_io_ins_down[9] ,
    \ces_2_5_io_ins_down[8] ,
    \ces_2_5_io_ins_down[7] ,
    \ces_2_5_io_ins_down[6] ,
    \ces_2_5_io_ins_down[5] ,
    \ces_2_5_io_ins_down[4] ,
    \ces_2_5_io_ins_down[3] ,
    \ces_2_5_io_ins_down[2] ,
    \ces_2_5_io_ins_down[1] ,
    \ces_2_5_io_ins_down[0] }),
    .io_outs_left({\ces_3_4_io_ins_left[63] ,
    \ces_3_4_io_ins_left[62] ,
    \ces_3_4_io_ins_left[61] ,
    \ces_3_4_io_ins_left[60] ,
    \ces_3_4_io_ins_left[59] ,
    \ces_3_4_io_ins_left[58] ,
    \ces_3_4_io_ins_left[57] ,
    \ces_3_4_io_ins_left[56] ,
    \ces_3_4_io_ins_left[55] ,
    \ces_3_4_io_ins_left[54] ,
    \ces_3_4_io_ins_left[53] ,
    \ces_3_4_io_ins_left[52] ,
    \ces_3_4_io_ins_left[51] ,
    \ces_3_4_io_ins_left[50] ,
    \ces_3_4_io_ins_left[49] ,
    \ces_3_4_io_ins_left[48] ,
    \ces_3_4_io_ins_left[47] ,
    \ces_3_4_io_ins_left[46] ,
    \ces_3_4_io_ins_left[45] ,
    \ces_3_4_io_ins_left[44] ,
    \ces_3_4_io_ins_left[43] ,
    \ces_3_4_io_ins_left[42] ,
    \ces_3_4_io_ins_left[41] ,
    \ces_3_4_io_ins_left[40] ,
    \ces_3_4_io_ins_left[39] ,
    \ces_3_4_io_ins_left[38] ,
    \ces_3_4_io_ins_left[37] ,
    \ces_3_4_io_ins_left[36] ,
    \ces_3_4_io_ins_left[35] ,
    \ces_3_4_io_ins_left[34] ,
    \ces_3_4_io_ins_left[33] ,
    \ces_3_4_io_ins_left[32] ,
    \ces_3_4_io_ins_left[31] ,
    \ces_3_4_io_ins_left[30] ,
    \ces_3_4_io_ins_left[29] ,
    \ces_3_4_io_ins_left[28] ,
    \ces_3_4_io_ins_left[27] ,
    \ces_3_4_io_ins_left[26] ,
    \ces_3_4_io_ins_left[25] ,
    \ces_3_4_io_ins_left[24] ,
    \ces_3_4_io_ins_left[23] ,
    \ces_3_4_io_ins_left[22] ,
    \ces_3_4_io_ins_left[21] ,
    \ces_3_4_io_ins_left[20] ,
    \ces_3_4_io_ins_left[19] ,
    \ces_3_4_io_ins_left[18] ,
    \ces_3_4_io_ins_left[17] ,
    \ces_3_4_io_ins_left[16] ,
    \ces_3_4_io_ins_left[15] ,
    \ces_3_4_io_ins_left[14] ,
    \ces_3_4_io_ins_left[13] ,
    \ces_3_4_io_ins_left[12] ,
    \ces_3_4_io_ins_left[11] ,
    \ces_3_4_io_ins_left[10] ,
    \ces_3_4_io_ins_left[9] ,
    \ces_3_4_io_ins_left[8] ,
    \ces_3_4_io_ins_left[7] ,
    \ces_3_4_io_ins_left[6] ,
    \ces_3_4_io_ins_left[5] ,
    \ces_3_4_io_ins_left[4] ,
    \ces_3_4_io_ins_left[3] ,
    \ces_3_4_io_ins_left[2] ,
    \ces_3_4_io_ins_left[1] ,
    \ces_3_4_io_ins_left[0] }),
    .io_outs_right({\ces_3_5_io_outs_right[63] ,
    \ces_3_5_io_outs_right[62] ,
    \ces_3_5_io_outs_right[61] ,
    \ces_3_5_io_outs_right[60] ,
    \ces_3_5_io_outs_right[59] ,
    \ces_3_5_io_outs_right[58] ,
    \ces_3_5_io_outs_right[57] ,
    \ces_3_5_io_outs_right[56] ,
    \ces_3_5_io_outs_right[55] ,
    \ces_3_5_io_outs_right[54] ,
    \ces_3_5_io_outs_right[53] ,
    \ces_3_5_io_outs_right[52] ,
    \ces_3_5_io_outs_right[51] ,
    \ces_3_5_io_outs_right[50] ,
    \ces_3_5_io_outs_right[49] ,
    \ces_3_5_io_outs_right[48] ,
    \ces_3_5_io_outs_right[47] ,
    \ces_3_5_io_outs_right[46] ,
    \ces_3_5_io_outs_right[45] ,
    \ces_3_5_io_outs_right[44] ,
    \ces_3_5_io_outs_right[43] ,
    \ces_3_5_io_outs_right[42] ,
    \ces_3_5_io_outs_right[41] ,
    \ces_3_5_io_outs_right[40] ,
    \ces_3_5_io_outs_right[39] ,
    \ces_3_5_io_outs_right[38] ,
    \ces_3_5_io_outs_right[37] ,
    \ces_3_5_io_outs_right[36] ,
    \ces_3_5_io_outs_right[35] ,
    \ces_3_5_io_outs_right[34] ,
    \ces_3_5_io_outs_right[33] ,
    \ces_3_5_io_outs_right[32] ,
    \ces_3_5_io_outs_right[31] ,
    \ces_3_5_io_outs_right[30] ,
    \ces_3_5_io_outs_right[29] ,
    \ces_3_5_io_outs_right[28] ,
    \ces_3_5_io_outs_right[27] ,
    \ces_3_5_io_outs_right[26] ,
    \ces_3_5_io_outs_right[25] ,
    \ces_3_5_io_outs_right[24] ,
    \ces_3_5_io_outs_right[23] ,
    \ces_3_5_io_outs_right[22] ,
    \ces_3_5_io_outs_right[21] ,
    \ces_3_5_io_outs_right[20] ,
    \ces_3_5_io_outs_right[19] ,
    \ces_3_5_io_outs_right[18] ,
    \ces_3_5_io_outs_right[17] ,
    \ces_3_5_io_outs_right[16] ,
    \ces_3_5_io_outs_right[15] ,
    \ces_3_5_io_outs_right[14] ,
    \ces_3_5_io_outs_right[13] ,
    \ces_3_5_io_outs_right[12] ,
    \ces_3_5_io_outs_right[11] ,
    \ces_3_5_io_outs_right[10] ,
    \ces_3_5_io_outs_right[9] ,
    \ces_3_5_io_outs_right[8] ,
    \ces_3_5_io_outs_right[7] ,
    \ces_3_5_io_outs_right[6] ,
    \ces_3_5_io_outs_right[5] ,
    \ces_3_5_io_outs_right[4] ,
    \ces_3_5_io_outs_right[3] ,
    \ces_3_5_io_outs_right[2] ,
    \ces_3_5_io_outs_right[1] ,
    \ces_3_5_io_outs_right[0] }),
    .io_outs_up({\ces_3_5_io_outs_up[63] ,
    \ces_3_5_io_outs_up[62] ,
    \ces_3_5_io_outs_up[61] ,
    \ces_3_5_io_outs_up[60] ,
    \ces_3_5_io_outs_up[59] ,
    \ces_3_5_io_outs_up[58] ,
    \ces_3_5_io_outs_up[57] ,
    \ces_3_5_io_outs_up[56] ,
    \ces_3_5_io_outs_up[55] ,
    \ces_3_5_io_outs_up[54] ,
    \ces_3_5_io_outs_up[53] ,
    \ces_3_5_io_outs_up[52] ,
    \ces_3_5_io_outs_up[51] ,
    \ces_3_5_io_outs_up[50] ,
    \ces_3_5_io_outs_up[49] ,
    \ces_3_5_io_outs_up[48] ,
    \ces_3_5_io_outs_up[47] ,
    \ces_3_5_io_outs_up[46] ,
    \ces_3_5_io_outs_up[45] ,
    \ces_3_5_io_outs_up[44] ,
    \ces_3_5_io_outs_up[43] ,
    \ces_3_5_io_outs_up[42] ,
    \ces_3_5_io_outs_up[41] ,
    \ces_3_5_io_outs_up[40] ,
    \ces_3_5_io_outs_up[39] ,
    \ces_3_5_io_outs_up[38] ,
    \ces_3_5_io_outs_up[37] ,
    \ces_3_5_io_outs_up[36] ,
    \ces_3_5_io_outs_up[35] ,
    \ces_3_5_io_outs_up[34] ,
    \ces_3_5_io_outs_up[33] ,
    \ces_3_5_io_outs_up[32] ,
    \ces_3_5_io_outs_up[31] ,
    \ces_3_5_io_outs_up[30] ,
    \ces_3_5_io_outs_up[29] ,
    \ces_3_5_io_outs_up[28] ,
    \ces_3_5_io_outs_up[27] ,
    \ces_3_5_io_outs_up[26] ,
    \ces_3_5_io_outs_up[25] ,
    \ces_3_5_io_outs_up[24] ,
    \ces_3_5_io_outs_up[23] ,
    \ces_3_5_io_outs_up[22] ,
    \ces_3_5_io_outs_up[21] ,
    \ces_3_5_io_outs_up[20] ,
    \ces_3_5_io_outs_up[19] ,
    \ces_3_5_io_outs_up[18] ,
    \ces_3_5_io_outs_up[17] ,
    \ces_3_5_io_outs_up[16] ,
    \ces_3_5_io_outs_up[15] ,
    \ces_3_5_io_outs_up[14] ,
    \ces_3_5_io_outs_up[13] ,
    \ces_3_5_io_outs_up[12] ,
    \ces_3_5_io_outs_up[11] ,
    \ces_3_5_io_outs_up[10] ,
    \ces_3_5_io_outs_up[9] ,
    \ces_3_5_io_outs_up[8] ,
    \ces_3_5_io_outs_up[7] ,
    \ces_3_5_io_outs_up[6] ,
    \ces_3_5_io_outs_up[5] ,
    \ces_3_5_io_outs_up[4] ,
    \ces_3_5_io_outs_up[3] ,
    \ces_3_5_io_outs_up[2] ,
    \ces_3_5_io_outs_up[1] ,
    \ces_3_5_io_outs_up[0] }));
 Element ces_3_6 (.clock(clknet_3_3_0_clock),
    .io_lsbIns_1(ces_3_5_io_lsbOuts_1),
    .io_lsbIns_2(ces_3_5_io_lsbOuts_2),
    .io_lsbIns_3(ces_3_5_io_lsbOuts_3),
    .io_lsbIns_4(ces_3_5_io_lsbOuts_4),
    .io_lsbIns_5(ces_3_5_io_lsbOuts_5),
    .io_lsbIns_6(ces_3_5_io_lsbOuts_6),
    .io_lsbIns_7(ces_3_5_io_lsbOuts_7),
    .io_lsbOuts_0(ces_3_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_6_io_lsbOuts_7),
    .io_ins_down({\ces_3_6_io_ins_down[63] ,
    \ces_3_6_io_ins_down[62] ,
    \ces_3_6_io_ins_down[61] ,
    \ces_3_6_io_ins_down[60] ,
    \ces_3_6_io_ins_down[59] ,
    \ces_3_6_io_ins_down[58] ,
    \ces_3_6_io_ins_down[57] ,
    \ces_3_6_io_ins_down[56] ,
    \ces_3_6_io_ins_down[55] ,
    \ces_3_6_io_ins_down[54] ,
    \ces_3_6_io_ins_down[53] ,
    \ces_3_6_io_ins_down[52] ,
    \ces_3_6_io_ins_down[51] ,
    \ces_3_6_io_ins_down[50] ,
    \ces_3_6_io_ins_down[49] ,
    \ces_3_6_io_ins_down[48] ,
    \ces_3_6_io_ins_down[47] ,
    \ces_3_6_io_ins_down[46] ,
    \ces_3_6_io_ins_down[45] ,
    \ces_3_6_io_ins_down[44] ,
    \ces_3_6_io_ins_down[43] ,
    \ces_3_6_io_ins_down[42] ,
    \ces_3_6_io_ins_down[41] ,
    \ces_3_6_io_ins_down[40] ,
    \ces_3_6_io_ins_down[39] ,
    \ces_3_6_io_ins_down[38] ,
    \ces_3_6_io_ins_down[37] ,
    \ces_3_6_io_ins_down[36] ,
    \ces_3_6_io_ins_down[35] ,
    \ces_3_6_io_ins_down[34] ,
    \ces_3_6_io_ins_down[33] ,
    \ces_3_6_io_ins_down[32] ,
    \ces_3_6_io_ins_down[31] ,
    \ces_3_6_io_ins_down[30] ,
    \ces_3_6_io_ins_down[29] ,
    \ces_3_6_io_ins_down[28] ,
    \ces_3_6_io_ins_down[27] ,
    \ces_3_6_io_ins_down[26] ,
    \ces_3_6_io_ins_down[25] ,
    \ces_3_6_io_ins_down[24] ,
    \ces_3_6_io_ins_down[23] ,
    \ces_3_6_io_ins_down[22] ,
    \ces_3_6_io_ins_down[21] ,
    \ces_3_6_io_ins_down[20] ,
    \ces_3_6_io_ins_down[19] ,
    \ces_3_6_io_ins_down[18] ,
    \ces_3_6_io_ins_down[17] ,
    \ces_3_6_io_ins_down[16] ,
    \ces_3_6_io_ins_down[15] ,
    \ces_3_6_io_ins_down[14] ,
    \ces_3_6_io_ins_down[13] ,
    \ces_3_6_io_ins_down[12] ,
    \ces_3_6_io_ins_down[11] ,
    \ces_3_6_io_ins_down[10] ,
    \ces_3_6_io_ins_down[9] ,
    \ces_3_6_io_ins_down[8] ,
    \ces_3_6_io_ins_down[7] ,
    \ces_3_6_io_ins_down[6] ,
    \ces_3_6_io_ins_down[5] ,
    \ces_3_6_io_ins_down[4] ,
    \ces_3_6_io_ins_down[3] ,
    \ces_3_6_io_ins_down[2] ,
    \ces_3_6_io_ins_down[1] ,
    \ces_3_6_io_ins_down[0] }),
    .io_ins_left({\ces_3_6_io_ins_left[63] ,
    \ces_3_6_io_ins_left[62] ,
    \ces_3_6_io_ins_left[61] ,
    \ces_3_6_io_ins_left[60] ,
    \ces_3_6_io_ins_left[59] ,
    \ces_3_6_io_ins_left[58] ,
    \ces_3_6_io_ins_left[57] ,
    \ces_3_6_io_ins_left[56] ,
    \ces_3_6_io_ins_left[55] ,
    \ces_3_6_io_ins_left[54] ,
    \ces_3_6_io_ins_left[53] ,
    \ces_3_6_io_ins_left[52] ,
    \ces_3_6_io_ins_left[51] ,
    \ces_3_6_io_ins_left[50] ,
    \ces_3_6_io_ins_left[49] ,
    \ces_3_6_io_ins_left[48] ,
    \ces_3_6_io_ins_left[47] ,
    \ces_3_6_io_ins_left[46] ,
    \ces_3_6_io_ins_left[45] ,
    \ces_3_6_io_ins_left[44] ,
    \ces_3_6_io_ins_left[43] ,
    \ces_3_6_io_ins_left[42] ,
    \ces_3_6_io_ins_left[41] ,
    \ces_3_6_io_ins_left[40] ,
    \ces_3_6_io_ins_left[39] ,
    \ces_3_6_io_ins_left[38] ,
    \ces_3_6_io_ins_left[37] ,
    \ces_3_6_io_ins_left[36] ,
    \ces_3_6_io_ins_left[35] ,
    \ces_3_6_io_ins_left[34] ,
    \ces_3_6_io_ins_left[33] ,
    \ces_3_6_io_ins_left[32] ,
    \ces_3_6_io_ins_left[31] ,
    \ces_3_6_io_ins_left[30] ,
    \ces_3_6_io_ins_left[29] ,
    \ces_3_6_io_ins_left[28] ,
    \ces_3_6_io_ins_left[27] ,
    \ces_3_6_io_ins_left[26] ,
    \ces_3_6_io_ins_left[25] ,
    \ces_3_6_io_ins_left[24] ,
    \ces_3_6_io_ins_left[23] ,
    \ces_3_6_io_ins_left[22] ,
    \ces_3_6_io_ins_left[21] ,
    \ces_3_6_io_ins_left[20] ,
    \ces_3_6_io_ins_left[19] ,
    \ces_3_6_io_ins_left[18] ,
    \ces_3_6_io_ins_left[17] ,
    \ces_3_6_io_ins_left[16] ,
    \ces_3_6_io_ins_left[15] ,
    \ces_3_6_io_ins_left[14] ,
    \ces_3_6_io_ins_left[13] ,
    \ces_3_6_io_ins_left[12] ,
    \ces_3_6_io_ins_left[11] ,
    \ces_3_6_io_ins_left[10] ,
    \ces_3_6_io_ins_left[9] ,
    \ces_3_6_io_ins_left[8] ,
    \ces_3_6_io_ins_left[7] ,
    \ces_3_6_io_ins_left[6] ,
    \ces_3_6_io_ins_left[5] ,
    \ces_3_6_io_ins_left[4] ,
    \ces_3_6_io_ins_left[3] ,
    \ces_3_6_io_ins_left[2] ,
    \ces_3_6_io_ins_left[1] ,
    \ces_3_6_io_ins_left[0] }),
    .io_ins_right({\ces_3_5_io_outs_right[63] ,
    \ces_3_5_io_outs_right[62] ,
    \ces_3_5_io_outs_right[61] ,
    \ces_3_5_io_outs_right[60] ,
    \ces_3_5_io_outs_right[59] ,
    \ces_3_5_io_outs_right[58] ,
    \ces_3_5_io_outs_right[57] ,
    \ces_3_5_io_outs_right[56] ,
    \ces_3_5_io_outs_right[55] ,
    \ces_3_5_io_outs_right[54] ,
    \ces_3_5_io_outs_right[53] ,
    \ces_3_5_io_outs_right[52] ,
    \ces_3_5_io_outs_right[51] ,
    \ces_3_5_io_outs_right[50] ,
    \ces_3_5_io_outs_right[49] ,
    \ces_3_5_io_outs_right[48] ,
    \ces_3_5_io_outs_right[47] ,
    \ces_3_5_io_outs_right[46] ,
    \ces_3_5_io_outs_right[45] ,
    \ces_3_5_io_outs_right[44] ,
    \ces_3_5_io_outs_right[43] ,
    \ces_3_5_io_outs_right[42] ,
    \ces_3_5_io_outs_right[41] ,
    \ces_3_5_io_outs_right[40] ,
    \ces_3_5_io_outs_right[39] ,
    \ces_3_5_io_outs_right[38] ,
    \ces_3_5_io_outs_right[37] ,
    \ces_3_5_io_outs_right[36] ,
    \ces_3_5_io_outs_right[35] ,
    \ces_3_5_io_outs_right[34] ,
    \ces_3_5_io_outs_right[33] ,
    \ces_3_5_io_outs_right[32] ,
    \ces_3_5_io_outs_right[31] ,
    \ces_3_5_io_outs_right[30] ,
    \ces_3_5_io_outs_right[29] ,
    \ces_3_5_io_outs_right[28] ,
    \ces_3_5_io_outs_right[27] ,
    \ces_3_5_io_outs_right[26] ,
    \ces_3_5_io_outs_right[25] ,
    \ces_3_5_io_outs_right[24] ,
    \ces_3_5_io_outs_right[23] ,
    \ces_3_5_io_outs_right[22] ,
    \ces_3_5_io_outs_right[21] ,
    \ces_3_5_io_outs_right[20] ,
    \ces_3_5_io_outs_right[19] ,
    \ces_3_5_io_outs_right[18] ,
    \ces_3_5_io_outs_right[17] ,
    \ces_3_5_io_outs_right[16] ,
    \ces_3_5_io_outs_right[15] ,
    \ces_3_5_io_outs_right[14] ,
    \ces_3_5_io_outs_right[13] ,
    \ces_3_5_io_outs_right[12] ,
    \ces_3_5_io_outs_right[11] ,
    \ces_3_5_io_outs_right[10] ,
    \ces_3_5_io_outs_right[9] ,
    \ces_3_5_io_outs_right[8] ,
    \ces_3_5_io_outs_right[7] ,
    \ces_3_5_io_outs_right[6] ,
    \ces_3_5_io_outs_right[5] ,
    \ces_3_5_io_outs_right[4] ,
    \ces_3_5_io_outs_right[3] ,
    \ces_3_5_io_outs_right[2] ,
    \ces_3_5_io_outs_right[1] ,
    \ces_3_5_io_outs_right[0] }),
    .io_ins_up({\ces_2_6_io_outs_up[63] ,
    \ces_2_6_io_outs_up[62] ,
    \ces_2_6_io_outs_up[61] ,
    \ces_2_6_io_outs_up[60] ,
    \ces_2_6_io_outs_up[59] ,
    \ces_2_6_io_outs_up[58] ,
    \ces_2_6_io_outs_up[57] ,
    \ces_2_6_io_outs_up[56] ,
    \ces_2_6_io_outs_up[55] ,
    \ces_2_6_io_outs_up[54] ,
    \ces_2_6_io_outs_up[53] ,
    \ces_2_6_io_outs_up[52] ,
    \ces_2_6_io_outs_up[51] ,
    \ces_2_6_io_outs_up[50] ,
    \ces_2_6_io_outs_up[49] ,
    \ces_2_6_io_outs_up[48] ,
    \ces_2_6_io_outs_up[47] ,
    \ces_2_6_io_outs_up[46] ,
    \ces_2_6_io_outs_up[45] ,
    \ces_2_6_io_outs_up[44] ,
    \ces_2_6_io_outs_up[43] ,
    \ces_2_6_io_outs_up[42] ,
    \ces_2_6_io_outs_up[41] ,
    \ces_2_6_io_outs_up[40] ,
    \ces_2_6_io_outs_up[39] ,
    \ces_2_6_io_outs_up[38] ,
    \ces_2_6_io_outs_up[37] ,
    \ces_2_6_io_outs_up[36] ,
    \ces_2_6_io_outs_up[35] ,
    \ces_2_6_io_outs_up[34] ,
    \ces_2_6_io_outs_up[33] ,
    \ces_2_6_io_outs_up[32] ,
    \ces_2_6_io_outs_up[31] ,
    \ces_2_6_io_outs_up[30] ,
    \ces_2_6_io_outs_up[29] ,
    \ces_2_6_io_outs_up[28] ,
    \ces_2_6_io_outs_up[27] ,
    \ces_2_6_io_outs_up[26] ,
    \ces_2_6_io_outs_up[25] ,
    \ces_2_6_io_outs_up[24] ,
    \ces_2_6_io_outs_up[23] ,
    \ces_2_6_io_outs_up[22] ,
    \ces_2_6_io_outs_up[21] ,
    \ces_2_6_io_outs_up[20] ,
    \ces_2_6_io_outs_up[19] ,
    \ces_2_6_io_outs_up[18] ,
    \ces_2_6_io_outs_up[17] ,
    \ces_2_6_io_outs_up[16] ,
    \ces_2_6_io_outs_up[15] ,
    \ces_2_6_io_outs_up[14] ,
    \ces_2_6_io_outs_up[13] ,
    \ces_2_6_io_outs_up[12] ,
    \ces_2_6_io_outs_up[11] ,
    \ces_2_6_io_outs_up[10] ,
    \ces_2_6_io_outs_up[9] ,
    \ces_2_6_io_outs_up[8] ,
    \ces_2_6_io_outs_up[7] ,
    \ces_2_6_io_outs_up[6] ,
    \ces_2_6_io_outs_up[5] ,
    \ces_2_6_io_outs_up[4] ,
    \ces_2_6_io_outs_up[3] ,
    \ces_2_6_io_outs_up[2] ,
    \ces_2_6_io_outs_up[1] ,
    \ces_2_6_io_outs_up[0] }),
    .io_outs_down({\ces_2_6_io_ins_down[63] ,
    \ces_2_6_io_ins_down[62] ,
    \ces_2_6_io_ins_down[61] ,
    \ces_2_6_io_ins_down[60] ,
    \ces_2_6_io_ins_down[59] ,
    \ces_2_6_io_ins_down[58] ,
    \ces_2_6_io_ins_down[57] ,
    \ces_2_6_io_ins_down[56] ,
    \ces_2_6_io_ins_down[55] ,
    \ces_2_6_io_ins_down[54] ,
    \ces_2_6_io_ins_down[53] ,
    \ces_2_6_io_ins_down[52] ,
    \ces_2_6_io_ins_down[51] ,
    \ces_2_6_io_ins_down[50] ,
    \ces_2_6_io_ins_down[49] ,
    \ces_2_6_io_ins_down[48] ,
    \ces_2_6_io_ins_down[47] ,
    \ces_2_6_io_ins_down[46] ,
    \ces_2_6_io_ins_down[45] ,
    \ces_2_6_io_ins_down[44] ,
    \ces_2_6_io_ins_down[43] ,
    \ces_2_6_io_ins_down[42] ,
    \ces_2_6_io_ins_down[41] ,
    \ces_2_6_io_ins_down[40] ,
    \ces_2_6_io_ins_down[39] ,
    \ces_2_6_io_ins_down[38] ,
    \ces_2_6_io_ins_down[37] ,
    \ces_2_6_io_ins_down[36] ,
    \ces_2_6_io_ins_down[35] ,
    \ces_2_6_io_ins_down[34] ,
    \ces_2_6_io_ins_down[33] ,
    \ces_2_6_io_ins_down[32] ,
    \ces_2_6_io_ins_down[31] ,
    \ces_2_6_io_ins_down[30] ,
    \ces_2_6_io_ins_down[29] ,
    \ces_2_6_io_ins_down[28] ,
    \ces_2_6_io_ins_down[27] ,
    \ces_2_6_io_ins_down[26] ,
    \ces_2_6_io_ins_down[25] ,
    \ces_2_6_io_ins_down[24] ,
    \ces_2_6_io_ins_down[23] ,
    \ces_2_6_io_ins_down[22] ,
    \ces_2_6_io_ins_down[21] ,
    \ces_2_6_io_ins_down[20] ,
    \ces_2_6_io_ins_down[19] ,
    \ces_2_6_io_ins_down[18] ,
    \ces_2_6_io_ins_down[17] ,
    \ces_2_6_io_ins_down[16] ,
    \ces_2_6_io_ins_down[15] ,
    \ces_2_6_io_ins_down[14] ,
    \ces_2_6_io_ins_down[13] ,
    \ces_2_6_io_ins_down[12] ,
    \ces_2_6_io_ins_down[11] ,
    \ces_2_6_io_ins_down[10] ,
    \ces_2_6_io_ins_down[9] ,
    \ces_2_6_io_ins_down[8] ,
    \ces_2_6_io_ins_down[7] ,
    \ces_2_6_io_ins_down[6] ,
    \ces_2_6_io_ins_down[5] ,
    \ces_2_6_io_ins_down[4] ,
    \ces_2_6_io_ins_down[3] ,
    \ces_2_6_io_ins_down[2] ,
    \ces_2_6_io_ins_down[1] ,
    \ces_2_6_io_ins_down[0] }),
    .io_outs_left({\ces_3_5_io_ins_left[63] ,
    \ces_3_5_io_ins_left[62] ,
    \ces_3_5_io_ins_left[61] ,
    \ces_3_5_io_ins_left[60] ,
    \ces_3_5_io_ins_left[59] ,
    \ces_3_5_io_ins_left[58] ,
    \ces_3_5_io_ins_left[57] ,
    \ces_3_5_io_ins_left[56] ,
    \ces_3_5_io_ins_left[55] ,
    \ces_3_5_io_ins_left[54] ,
    \ces_3_5_io_ins_left[53] ,
    \ces_3_5_io_ins_left[52] ,
    \ces_3_5_io_ins_left[51] ,
    \ces_3_5_io_ins_left[50] ,
    \ces_3_5_io_ins_left[49] ,
    \ces_3_5_io_ins_left[48] ,
    \ces_3_5_io_ins_left[47] ,
    \ces_3_5_io_ins_left[46] ,
    \ces_3_5_io_ins_left[45] ,
    \ces_3_5_io_ins_left[44] ,
    \ces_3_5_io_ins_left[43] ,
    \ces_3_5_io_ins_left[42] ,
    \ces_3_5_io_ins_left[41] ,
    \ces_3_5_io_ins_left[40] ,
    \ces_3_5_io_ins_left[39] ,
    \ces_3_5_io_ins_left[38] ,
    \ces_3_5_io_ins_left[37] ,
    \ces_3_5_io_ins_left[36] ,
    \ces_3_5_io_ins_left[35] ,
    \ces_3_5_io_ins_left[34] ,
    \ces_3_5_io_ins_left[33] ,
    \ces_3_5_io_ins_left[32] ,
    \ces_3_5_io_ins_left[31] ,
    \ces_3_5_io_ins_left[30] ,
    \ces_3_5_io_ins_left[29] ,
    \ces_3_5_io_ins_left[28] ,
    \ces_3_5_io_ins_left[27] ,
    \ces_3_5_io_ins_left[26] ,
    \ces_3_5_io_ins_left[25] ,
    \ces_3_5_io_ins_left[24] ,
    \ces_3_5_io_ins_left[23] ,
    \ces_3_5_io_ins_left[22] ,
    \ces_3_5_io_ins_left[21] ,
    \ces_3_5_io_ins_left[20] ,
    \ces_3_5_io_ins_left[19] ,
    \ces_3_5_io_ins_left[18] ,
    \ces_3_5_io_ins_left[17] ,
    \ces_3_5_io_ins_left[16] ,
    \ces_3_5_io_ins_left[15] ,
    \ces_3_5_io_ins_left[14] ,
    \ces_3_5_io_ins_left[13] ,
    \ces_3_5_io_ins_left[12] ,
    \ces_3_5_io_ins_left[11] ,
    \ces_3_5_io_ins_left[10] ,
    \ces_3_5_io_ins_left[9] ,
    \ces_3_5_io_ins_left[8] ,
    \ces_3_5_io_ins_left[7] ,
    \ces_3_5_io_ins_left[6] ,
    \ces_3_5_io_ins_left[5] ,
    \ces_3_5_io_ins_left[4] ,
    \ces_3_5_io_ins_left[3] ,
    \ces_3_5_io_ins_left[2] ,
    \ces_3_5_io_ins_left[1] ,
    \ces_3_5_io_ins_left[0] }),
    .io_outs_right({\ces_3_6_io_outs_right[63] ,
    \ces_3_6_io_outs_right[62] ,
    \ces_3_6_io_outs_right[61] ,
    \ces_3_6_io_outs_right[60] ,
    \ces_3_6_io_outs_right[59] ,
    \ces_3_6_io_outs_right[58] ,
    \ces_3_6_io_outs_right[57] ,
    \ces_3_6_io_outs_right[56] ,
    \ces_3_6_io_outs_right[55] ,
    \ces_3_6_io_outs_right[54] ,
    \ces_3_6_io_outs_right[53] ,
    \ces_3_6_io_outs_right[52] ,
    \ces_3_6_io_outs_right[51] ,
    \ces_3_6_io_outs_right[50] ,
    \ces_3_6_io_outs_right[49] ,
    \ces_3_6_io_outs_right[48] ,
    \ces_3_6_io_outs_right[47] ,
    \ces_3_6_io_outs_right[46] ,
    \ces_3_6_io_outs_right[45] ,
    \ces_3_6_io_outs_right[44] ,
    \ces_3_6_io_outs_right[43] ,
    \ces_3_6_io_outs_right[42] ,
    \ces_3_6_io_outs_right[41] ,
    \ces_3_6_io_outs_right[40] ,
    \ces_3_6_io_outs_right[39] ,
    \ces_3_6_io_outs_right[38] ,
    \ces_3_6_io_outs_right[37] ,
    \ces_3_6_io_outs_right[36] ,
    \ces_3_6_io_outs_right[35] ,
    \ces_3_6_io_outs_right[34] ,
    \ces_3_6_io_outs_right[33] ,
    \ces_3_6_io_outs_right[32] ,
    \ces_3_6_io_outs_right[31] ,
    \ces_3_6_io_outs_right[30] ,
    \ces_3_6_io_outs_right[29] ,
    \ces_3_6_io_outs_right[28] ,
    \ces_3_6_io_outs_right[27] ,
    \ces_3_6_io_outs_right[26] ,
    \ces_3_6_io_outs_right[25] ,
    \ces_3_6_io_outs_right[24] ,
    \ces_3_6_io_outs_right[23] ,
    \ces_3_6_io_outs_right[22] ,
    \ces_3_6_io_outs_right[21] ,
    \ces_3_6_io_outs_right[20] ,
    \ces_3_6_io_outs_right[19] ,
    \ces_3_6_io_outs_right[18] ,
    \ces_3_6_io_outs_right[17] ,
    \ces_3_6_io_outs_right[16] ,
    \ces_3_6_io_outs_right[15] ,
    \ces_3_6_io_outs_right[14] ,
    \ces_3_6_io_outs_right[13] ,
    \ces_3_6_io_outs_right[12] ,
    \ces_3_6_io_outs_right[11] ,
    \ces_3_6_io_outs_right[10] ,
    \ces_3_6_io_outs_right[9] ,
    \ces_3_6_io_outs_right[8] ,
    \ces_3_6_io_outs_right[7] ,
    \ces_3_6_io_outs_right[6] ,
    \ces_3_6_io_outs_right[5] ,
    \ces_3_6_io_outs_right[4] ,
    \ces_3_6_io_outs_right[3] ,
    \ces_3_6_io_outs_right[2] ,
    \ces_3_6_io_outs_right[1] ,
    \ces_3_6_io_outs_right[0] }),
    .io_outs_up({\ces_3_6_io_outs_up[63] ,
    \ces_3_6_io_outs_up[62] ,
    \ces_3_6_io_outs_up[61] ,
    \ces_3_6_io_outs_up[60] ,
    \ces_3_6_io_outs_up[59] ,
    \ces_3_6_io_outs_up[58] ,
    \ces_3_6_io_outs_up[57] ,
    \ces_3_6_io_outs_up[56] ,
    \ces_3_6_io_outs_up[55] ,
    \ces_3_6_io_outs_up[54] ,
    \ces_3_6_io_outs_up[53] ,
    \ces_3_6_io_outs_up[52] ,
    \ces_3_6_io_outs_up[51] ,
    \ces_3_6_io_outs_up[50] ,
    \ces_3_6_io_outs_up[49] ,
    \ces_3_6_io_outs_up[48] ,
    \ces_3_6_io_outs_up[47] ,
    \ces_3_6_io_outs_up[46] ,
    \ces_3_6_io_outs_up[45] ,
    \ces_3_6_io_outs_up[44] ,
    \ces_3_6_io_outs_up[43] ,
    \ces_3_6_io_outs_up[42] ,
    \ces_3_6_io_outs_up[41] ,
    \ces_3_6_io_outs_up[40] ,
    \ces_3_6_io_outs_up[39] ,
    \ces_3_6_io_outs_up[38] ,
    \ces_3_6_io_outs_up[37] ,
    \ces_3_6_io_outs_up[36] ,
    \ces_3_6_io_outs_up[35] ,
    \ces_3_6_io_outs_up[34] ,
    \ces_3_6_io_outs_up[33] ,
    \ces_3_6_io_outs_up[32] ,
    \ces_3_6_io_outs_up[31] ,
    \ces_3_6_io_outs_up[30] ,
    \ces_3_6_io_outs_up[29] ,
    \ces_3_6_io_outs_up[28] ,
    \ces_3_6_io_outs_up[27] ,
    \ces_3_6_io_outs_up[26] ,
    \ces_3_6_io_outs_up[25] ,
    \ces_3_6_io_outs_up[24] ,
    \ces_3_6_io_outs_up[23] ,
    \ces_3_6_io_outs_up[22] ,
    \ces_3_6_io_outs_up[21] ,
    \ces_3_6_io_outs_up[20] ,
    \ces_3_6_io_outs_up[19] ,
    \ces_3_6_io_outs_up[18] ,
    \ces_3_6_io_outs_up[17] ,
    \ces_3_6_io_outs_up[16] ,
    \ces_3_6_io_outs_up[15] ,
    \ces_3_6_io_outs_up[14] ,
    \ces_3_6_io_outs_up[13] ,
    \ces_3_6_io_outs_up[12] ,
    \ces_3_6_io_outs_up[11] ,
    \ces_3_6_io_outs_up[10] ,
    \ces_3_6_io_outs_up[9] ,
    \ces_3_6_io_outs_up[8] ,
    \ces_3_6_io_outs_up[7] ,
    \ces_3_6_io_outs_up[6] ,
    \ces_3_6_io_outs_up[5] ,
    \ces_3_6_io_outs_up[4] ,
    \ces_3_6_io_outs_up[3] ,
    \ces_3_6_io_outs_up[2] ,
    \ces_3_6_io_outs_up[1] ,
    \ces_3_6_io_outs_up[0] }));
 Element ces_3_7 (.clock(clknet_3_3_0_clock),
    .io_lsbIns_1(ces_3_6_io_lsbOuts_1),
    .io_lsbIns_2(ces_3_6_io_lsbOuts_2),
    .io_lsbIns_3(ces_3_6_io_lsbOuts_3),
    .io_lsbIns_4(ces_3_6_io_lsbOuts_4),
    .io_lsbIns_5(ces_3_6_io_lsbOuts_5),
    .io_lsbIns_6(ces_3_6_io_lsbOuts_6),
    .io_lsbIns_7(ces_3_6_io_lsbOuts_7),
    .io_lsbOuts_0(ces_3_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_3_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_3_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_3_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_3_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_3_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_3_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_3_7_io_lsbOuts_7),
    .io_ins_down({\ces_3_7_io_ins_down[63] ,
    \ces_3_7_io_ins_down[62] ,
    \ces_3_7_io_ins_down[61] ,
    \ces_3_7_io_ins_down[60] ,
    \ces_3_7_io_ins_down[59] ,
    \ces_3_7_io_ins_down[58] ,
    \ces_3_7_io_ins_down[57] ,
    \ces_3_7_io_ins_down[56] ,
    \ces_3_7_io_ins_down[55] ,
    \ces_3_7_io_ins_down[54] ,
    \ces_3_7_io_ins_down[53] ,
    \ces_3_7_io_ins_down[52] ,
    \ces_3_7_io_ins_down[51] ,
    \ces_3_7_io_ins_down[50] ,
    \ces_3_7_io_ins_down[49] ,
    \ces_3_7_io_ins_down[48] ,
    \ces_3_7_io_ins_down[47] ,
    \ces_3_7_io_ins_down[46] ,
    \ces_3_7_io_ins_down[45] ,
    \ces_3_7_io_ins_down[44] ,
    \ces_3_7_io_ins_down[43] ,
    \ces_3_7_io_ins_down[42] ,
    \ces_3_7_io_ins_down[41] ,
    \ces_3_7_io_ins_down[40] ,
    \ces_3_7_io_ins_down[39] ,
    \ces_3_7_io_ins_down[38] ,
    \ces_3_7_io_ins_down[37] ,
    \ces_3_7_io_ins_down[36] ,
    \ces_3_7_io_ins_down[35] ,
    \ces_3_7_io_ins_down[34] ,
    \ces_3_7_io_ins_down[33] ,
    \ces_3_7_io_ins_down[32] ,
    \ces_3_7_io_ins_down[31] ,
    \ces_3_7_io_ins_down[30] ,
    \ces_3_7_io_ins_down[29] ,
    \ces_3_7_io_ins_down[28] ,
    \ces_3_7_io_ins_down[27] ,
    \ces_3_7_io_ins_down[26] ,
    \ces_3_7_io_ins_down[25] ,
    \ces_3_7_io_ins_down[24] ,
    \ces_3_7_io_ins_down[23] ,
    \ces_3_7_io_ins_down[22] ,
    \ces_3_7_io_ins_down[21] ,
    \ces_3_7_io_ins_down[20] ,
    \ces_3_7_io_ins_down[19] ,
    \ces_3_7_io_ins_down[18] ,
    \ces_3_7_io_ins_down[17] ,
    \ces_3_7_io_ins_down[16] ,
    \ces_3_7_io_ins_down[15] ,
    \ces_3_7_io_ins_down[14] ,
    \ces_3_7_io_ins_down[13] ,
    \ces_3_7_io_ins_down[12] ,
    \ces_3_7_io_ins_down[11] ,
    \ces_3_7_io_ins_down[10] ,
    \ces_3_7_io_ins_down[9] ,
    \ces_3_7_io_ins_down[8] ,
    \ces_3_7_io_ins_down[7] ,
    \ces_3_7_io_ins_down[6] ,
    \ces_3_7_io_ins_down[5] ,
    \ces_3_7_io_ins_down[4] ,
    \ces_3_7_io_ins_down[3] ,
    \ces_3_7_io_ins_down[2] ,
    \ces_3_7_io_ins_down[1] ,
    \ces_3_7_io_ins_down[0] }),
    .io_ins_left({net764,
    net763,
    net762,
    net761,
    net759,
    net758,
    net757,
    net756,
    net755,
    net754,
    net753,
    net752,
    net751,
    net750,
    net748,
    net747,
    net746,
    net745,
    net744,
    net743,
    net742,
    net741,
    net740,
    net739,
    net737,
    net736,
    net735,
    net734,
    net733,
    net732,
    net731,
    net730,
    net729,
    net728,
    net726,
    net725,
    net724,
    net723,
    net722,
    net721,
    net720,
    net719,
    net718,
    net717,
    net715,
    net714,
    net713,
    net712,
    net711,
    net710,
    net709,
    net708,
    net707,
    net706,
    net768,
    net767,
    net766,
    net765,
    net760,
    net749,
    net738,
    net727,
    net716,
    net705}),
    .io_ins_right({\ces_3_6_io_outs_right[63] ,
    \ces_3_6_io_outs_right[62] ,
    \ces_3_6_io_outs_right[61] ,
    \ces_3_6_io_outs_right[60] ,
    \ces_3_6_io_outs_right[59] ,
    \ces_3_6_io_outs_right[58] ,
    \ces_3_6_io_outs_right[57] ,
    \ces_3_6_io_outs_right[56] ,
    \ces_3_6_io_outs_right[55] ,
    \ces_3_6_io_outs_right[54] ,
    \ces_3_6_io_outs_right[53] ,
    \ces_3_6_io_outs_right[52] ,
    \ces_3_6_io_outs_right[51] ,
    \ces_3_6_io_outs_right[50] ,
    \ces_3_6_io_outs_right[49] ,
    \ces_3_6_io_outs_right[48] ,
    \ces_3_6_io_outs_right[47] ,
    \ces_3_6_io_outs_right[46] ,
    \ces_3_6_io_outs_right[45] ,
    \ces_3_6_io_outs_right[44] ,
    \ces_3_6_io_outs_right[43] ,
    \ces_3_6_io_outs_right[42] ,
    \ces_3_6_io_outs_right[41] ,
    \ces_3_6_io_outs_right[40] ,
    \ces_3_6_io_outs_right[39] ,
    \ces_3_6_io_outs_right[38] ,
    \ces_3_6_io_outs_right[37] ,
    \ces_3_6_io_outs_right[36] ,
    \ces_3_6_io_outs_right[35] ,
    \ces_3_6_io_outs_right[34] ,
    \ces_3_6_io_outs_right[33] ,
    \ces_3_6_io_outs_right[32] ,
    \ces_3_6_io_outs_right[31] ,
    \ces_3_6_io_outs_right[30] ,
    \ces_3_6_io_outs_right[29] ,
    \ces_3_6_io_outs_right[28] ,
    \ces_3_6_io_outs_right[27] ,
    \ces_3_6_io_outs_right[26] ,
    \ces_3_6_io_outs_right[25] ,
    \ces_3_6_io_outs_right[24] ,
    \ces_3_6_io_outs_right[23] ,
    \ces_3_6_io_outs_right[22] ,
    \ces_3_6_io_outs_right[21] ,
    \ces_3_6_io_outs_right[20] ,
    \ces_3_6_io_outs_right[19] ,
    \ces_3_6_io_outs_right[18] ,
    \ces_3_6_io_outs_right[17] ,
    \ces_3_6_io_outs_right[16] ,
    \ces_3_6_io_outs_right[15] ,
    \ces_3_6_io_outs_right[14] ,
    \ces_3_6_io_outs_right[13] ,
    \ces_3_6_io_outs_right[12] ,
    \ces_3_6_io_outs_right[11] ,
    \ces_3_6_io_outs_right[10] ,
    \ces_3_6_io_outs_right[9] ,
    \ces_3_6_io_outs_right[8] ,
    \ces_3_6_io_outs_right[7] ,
    \ces_3_6_io_outs_right[6] ,
    \ces_3_6_io_outs_right[5] ,
    \ces_3_6_io_outs_right[4] ,
    \ces_3_6_io_outs_right[3] ,
    \ces_3_6_io_outs_right[2] ,
    \ces_3_6_io_outs_right[1] ,
    \ces_3_6_io_outs_right[0] }),
    .io_ins_up({\ces_2_7_io_outs_up[63] ,
    \ces_2_7_io_outs_up[62] ,
    \ces_2_7_io_outs_up[61] ,
    \ces_2_7_io_outs_up[60] ,
    \ces_2_7_io_outs_up[59] ,
    \ces_2_7_io_outs_up[58] ,
    \ces_2_7_io_outs_up[57] ,
    \ces_2_7_io_outs_up[56] ,
    \ces_2_7_io_outs_up[55] ,
    \ces_2_7_io_outs_up[54] ,
    \ces_2_7_io_outs_up[53] ,
    \ces_2_7_io_outs_up[52] ,
    \ces_2_7_io_outs_up[51] ,
    \ces_2_7_io_outs_up[50] ,
    \ces_2_7_io_outs_up[49] ,
    \ces_2_7_io_outs_up[48] ,
    \ces_2_7_io_outs_up[47] ,
    \ces_2_7_io_outs_up[46] ,
    \ces_2_7_io_outs_up[45] ,
    \ces_2_7_io_outs_up[44] ,
    \ces_2_7_io_outs_up[43] ,
    \ces_2_7_io_outs_up[42] ,
    \ces_2_7_io_outs_up[41] ,
    \ces_2_7_io_outs_up[40] ,
    \ces_2_7_io_outs_up[39] ,
    \ces_2_7_io_outs_up[38] ,
    \ces_2_7_io_outs_up[37] ,
    \ces_2_7_io_outs_up[36] ,
    \ces_2_7_io_outs_up[35] ,
    \ces_2_7_io_outs_up[34] ,
    \ces_2_7_io_outs_up[33] ,
    \ces_2_7_io_outs_up[32] ,
    \ces_2_7_io_outs_up[31] ,
    \ces_2_7_io_outs_up[30] ,
    \ces_2_7_io_outs_up[29] ,
    \ces_2_7_io_outs_up[28] ,
    \ces_2_7_io_outs_up[27] ,
    \ces_2_7_io_outs_up[26] ,
    \ces_2_7_io_outs_up[25] ,
    \ces_2_7_io_outs_up[24] ,
    \ces_2_7_io_outs_up[23] ,
    \ces_2_7_io_outs_up[22] ,
    \ces_2_7_io_outs_up[21] ,
    \ces_2_7_io_outs_up[20] ,
    \ces_2_7_io_outs_up[19] ,
    \ces_2_7_io_outs_up[18] ,
    \ces_2_7_io_outs_up[17] ,
    \ces_2_7_io_outs_up[16] ,
    \ces_2_7_io_outs_up[15] ,
    \ces_2_7_io_outs_up[14] ,
    \ces_2_7_io_outs_up[13] ,
    \ces_2_7_io_outs_up[12] ,
    \ces_2_7_io_outs_up[11] ,
    \ces_2_7_io_outs_up[10] ,
    \ces_2_7_io_outs_up[9] ,
    \ces_2_7_io_outs_up[8] ,
    \ces_2_7_io_outs_up[7] ,
    \ces_2_7_io_outs_up[6] ,
    \ces_2_7_io_outs_up[5] ,
    \ces_2_7_io_outs_up[4] ,
    \ces_2_7_io_outs_up[3] ,
    \ces_2_7_io_outs_up[2] ,
    \ces_2_7_io_outs_up[1] ,
    \ces_2_7_io_outs_up[0] }),
    .io_outs_down({\ces_2_7_io_ins_down[63] ,
    \ces_2_7_io_ins_down[62] ,
    \ces_2_7_io_ins_down[61] ,
    \ces_2_7_io_ins_down[60] ,
    \ces_2_7_io_ins_down[59] ,
    \ces_2_7_io_ins_down[58] ,
    \ces_2_7_io_ins_down[57] ,
    \ces_2_7_io_ins_down[56] ,
    \ces_2_7_io_ins_down[55] ,
    \ces_2_7_io_ins_down[54] ,
    \ces_2_7_io_ins_down[53] ,
    \ces_2_7_io_ins_down[52] ,
    \ces_2_7_io_ins_down[51] ,
    \ces_2_7_io_ins_down[50] ,
    \ces_2_7_io_ins_down[49] ,
    \ces_2_7_io_ins_down[48] ,
    \ces_2_7_io_ins_down[47] ,
    \ces_2_7_io_ins_down[46] ,
    \ces_2_7_io_ins_down[45] ,
    \ces_2_7_io_ins_down[44] ,
    \ces_2_7_io_ins_down[43] ,
    \ces_2_7_io_ins_down[42] ,
    \ces_2_7_io_ins_down[41] ,
    \ces_2_7_io_ins_down[40] ,
    \ces_2_7_io_ins_down[39] ,
    \ces_2_7_io_ins_down[38] ,
    \ces_2_7_io_ins_down[37] ,
    \ces_2_7_io_ins_down[36] ,
    \ces_2_7_io_ins_down[35] ,
    \ces_2_7_io_ins_down[34] ,
    \ces_2_7_io_ins_down[33] ,
    \ces_2_7_io_ins_down[32] ,
    \ces_2_7_io_ins_down[31] ,
    \ces_2_7_io_ins_down[30] ,
    \ces_2_7_io_ins_down[29] ,
    \ces_2_7_io_ins_down[28] ,
    \ces_2_7_io_ins_down[27] ,
    \ces_2_7_io_ins_down[26] ,
    \ces_2_7_io_ins_down[25] ,
    \ces_2_7_io_ins_down[24] ,
    \ces_2_7_io_ins_down[23] ,
    \ces_2_7_io_ins_down[22] ,
    \ces_2_7_io_ins_down[21] ,
    \ces_2_7_io_ins_down[20] ,
    \ces_2_7_io_ins_down[19] ,
    \ces_2_7_io_ins_down[18] ,
    \ces_2_7_io_ins_down[17] ,
    \ces_2_7_io_ins_down[16] ,
    \ces_2_7_io_ins_down[15] ,
    \ces_2_7_io_ins_down[14] ,
    \ces_2_7_io_ins_down[13] ,
    \ces_2_7_io_ins_down[12] ,
    \ces_2_7_io_ins_down[11] ,
    \ces_2_7_io_ins_down[10] ,
    \ces_2_7_io_ins_down[9] ,
    \ces_2_7_io_ins_down[8] ,
    \ces_2_7_io_ins_down[7] ,
    \ces_2_7_io_ins_down[6] ,
    \ces_2_7_io_ins_down[5] ,
    \ces_2_7_io_ins_down[4] ,
    \ces_2_7_io_ins_down[3] ,
    \ces_2_7_io_ins_down[2] ,
    \ces_2_7_io_ins_down[1] ,
    \ces_2_7_io_ins_down[0] }),
    .io_outs_left({\ces_3_6_io_ins_left[63] ,
    \ces_3_6_io_ins_left[62] ,
    \ces_3_6_io_ins_left[61] ,
    \ces_3_6_io_ins_left[60] ,
    \ces_3_6_io_ins_left[59] ,
    \ces_3_6_io_ins_left[58] ,
    \ces_3_6_io_ins_left[57] ,
    \ces_3_6_io_ins_left[56] ,
    \ces_3_6_io_ins_left[55] ,
    \ces_3_6_io_ins_left[54] ,
    \ces_3_6_io_ins_left[53] ,
    \ces_3_6_io_ins_left[52] ,
    \ces_3_6_io_ins_left[51] ,
    \ces_3_6_io_ins_left[50] ,
    \ces_3_6_io_ins_left[49] ,
    \ces_3_6_io_ins_left[48] ,
    \ces_3_6_io_ins_left[47] ,
    \ces_3_6_io_ins_left[46] ,
    \ces_3_6_io_ins_left[45] ,
    \ces_3_6_io_ins_left[44] ,
    \ces_3_6_io_ins_left[43] ,
    \ces_3_6_io_ins_left[42] ,
    \ces_3_6_io_ins_left[41] ,
    \ces_3_6_io_ins_left[40] ,
    \ces_3_6_io_ins_left[39] ,
    \ces_3_6_io_ins_left[38] ,
    \ces_3_6_io_ins_left[37] ,
    \ces_3_6_io_ins_left[36] ,
    \ces_3_6_io_ins_left[35] ,
    \ces_3_6_io_ins_left[34] ,
    \ces_3_6_io_ins_left[33] ,
    \ces_3_6_io_ins_left[32] ,
    \ces_3_6_io_ins_left[31] ,
    \ces_3_6_io_ins_left[30] ,
    \ces_3_6_io_ins_left[29] ,
    \ces_3_6_io_ins_left[28] ,
    \ces_3_6_io_ins_left[27] ,
    \ces_3_6_io_ins_left[26] ,
    \ces_3_6_io_ins_left[25] ,
    \ces_3_6_io_ins_left[24] ,
    \ces_3_6_io_ins_left[23] ,
    \ces_3_6_io_ins_left[22] ,
    \ces_3_6_io_ins_left[21] ,
    \ces_3_6_io_ins_left[20] ,
    \ces_3_6_io_ins_left[19] ,
    \ces_3_6_io_ins_left[18] ,
    \ces_3_6_io_ins_left[17] ,
    \ces_3_6_io_ins_left[16] ,
    \ces_3_6_io_ins_left[15] ,
    \ces_3_6_io_ins_left[14] ,
    \ces_3_6_io_ins_left[13] ,
    \ces_3_6_io_ins_left[12] ,
    \ces_3_6_io_ins_left[11] ,
    \ces_3_6_io_ins_left[10] ,
    \ces_3_6_io_ins_left[9] ,
    \ces_3_6_io_ins_left[8] ,
    \ces_3_6_io_ins_left[7] ,
    \ces_3_6_io_ins_left[6] ,
    \ces_3_6_io_ins_left[5] ,
    \ces_3_6_io_ins_left[4] ,
    \ces_3_6_io_ins_left[3] ,
    \ces_3_6_io_ins_left[2] ,
    \ces_3_6_io_ins_left[1] ,
    \ces_3_6_io_ins_left[0] }),
    .io_outs_right({net3388,
    net3387,
    net3386,
    net3385,
    net3383,
    net3382,
    net3381,
    net3380,
    net3379,
    net3378,
    net3377,
    net3376,
    net3375,
    net3374,
    net3372,
    net3371,
    net3370,
    net3369,
    net3368,
    net3367,
    net3366,
    net3365,
    net3364,
    net3363,
    net3361,
    net3360,
    net3359,
    net3358,
    net3357,
    net3356,
    net3355,
    net3354,
    net3353,
    net3352,
    net3350,
    net3349,
    net3348,
    net3347,
    net3346,
    net3345,
    net3344,
    net3343,
    net3342,
    net3341,
    net3339,
    net3338,
    net3337,
    net3336,
    net3335,
    net3334,
    net3333,
    net3332,
    net3331,
    net3330,
    net3392,
    net3391,
    net3390,
    net3389,
    net3384,
    net3373,
    net3362,
    net3351,
    net3340,
    net3329}),
    .io_outs_up({\ces_3_7_io_outs_up[63] ,
    \ces_3_7_io_outs_up[62] ,
    \ces_3_7_io_outs_up[61] ,
    \ces_3_7_io_outs_up[60] ,
    \ces_3_7_io_outs_up[59] ,
    \ces_3_7_io_outs_up[58] ,
    \ces_3_7_io_outs_up[57] ,
    \ces_3_7_io_outs_up[56] ,
    \ces_3_7_io_outs_up[55] ,
    \ces_3_7_io_outs_up[54] ,
    \ces_3_7_io_outs_up[53] ,
    \ces_3_7_io_outs_up[52] ,
    \ces_3_7_io_outs_up[51] ,
    \ces_3_7_io_outs_up[50] ,
    \ces_3_7_io_outs_up[49] ,
    \ces_3_7_io_outs_up[48] ,
    \ces_3_7_io_outs_up[47] ,
    \ces_3_7_io_outs_up[46] ,
    \ces_3_7_io_outs_up[45] ,
    \ces_3_7_io_outs_up[44] ,
    \ces_3_7_io_outs_up[43] ,
    \ces_3_7_io_outs_up[42] ,
    \ces_3_7_io_outs_up[41] ,
    \ces_3_7_io_outs_up[40] ,
    \ces_3_7_io_outs_up[39] ,
    \ces_3_7_io_outs_up[38] ,
    \ces_3_7_io_outs_up[37] ,
    \ces_3_7_io_outs_up[36] ,
    \ces_3_7_io_outs_up[35] ,
    \ces_3_7_io_outs_up[34] ,
    \ces_3_7_io_outs_up[33] ,
    \ces_3_7_io_outs_up[32] ,
    \ces_3_7_io_outs_up[31] ,
    \ces_3_7_io_outs_up[30] ,
    \ces_3_7_io_outs_up[29] ,
    \ces_3_7_io_outs_up[28] ,
    \ces_3_7_io_outs_up[27] ,
    \ces_3_7_io_outs_up[26] ,
    \ces_3_7_io_outs_up[25] ,
    \ces_3_7_io_outs_up[24] ,
    \ces_3_7_io_outs_up[23] ,
    \ces_3_7_io_outs_up[22] ,
    \ces_3_7_io_outs_up[21] ,
    \ces_3_7_io_outs_up[20] ,
    \ces_3_7_io_outs_up[19] ,
    \ces_3_7_io_outs_up[18] ,
    \ces_3_7_io_outs_up[17] ,
    \ces_3_7_io_outs_up[16] ,
    \ces_3_7_io_outs_up[15] ,
    \ces_3_7_io_outs_up[14] ,
    \ces_3_7_io_outs_up[13] ,
    \ces_3_7_io_outs_up[12] ,
    \ces_3_7_io_outs_up[11] ,
    \ces_3_7_io_outs_up[10] ,
    \ces_3_7_io_outs_up[9] ,
    \ces_3_7_io_outs_up[8] ,
    \ces_3_7_io_outs_up[7] ,
    \ces_3_7_io_outs_up[6] ,
    \ces_3_7_io_outs_up[5] ,
    \ces_3_7_io_outs_up[4] ,
    \ces_3_7_io_outs_up[3] ,
    \ces_3_7_io_outs_up[2] ,
    \ces_3_7_io_outs_up[1] ,
    \ces_3_7_io_outs_up[0] }));
 Element ces_4_0 (.clock(clknet_3_4_0_clock),
    .io_lsbIns_1(net4189),
    .io_lsbIns_2(net4190),
    .io_lsbIns_3(net4191),
    .io_lsbIns_4(net4192),
    .io_lsbIns_5(net4193),
    .io_lsbIns_6(net4194),
    .io_lsbIns_7(net4195),
    .io_lsbOuts_0(ces_4_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_0_io_lsbOuts_7),
    .io_ins_down({\ces_4_0_io_ins_down[63] ,
    \ces_4_0_io_ins_down[62] ,
    \ces_4_0_io_ins_down[61] ,
    \ces_4_0_io_ins_down[60] ,
    \ces_4_0_io_ins_down[59] ,
    \ces_4_0_io_ins_down[58] ,
    \ces_4_0_io_ins_down[57] ,
    \ces_4_0_io_ins_down[56] ,
    \ces_4_0_io_ins_down[55] ,
    \ces_4_0_io_ins_down[54] ,
    \ces_4_0_io_ins_down[53] ,
    \ces_4_0_io_ins_down[52] ,
    \ces_4_0_io_ins_down[51] ,
    \ces_4_0_io_ins_down[50] ,
    \ces_4_0_io_ins_down[49] ,
    \ces_4_0_io_ins_down[48] ,
    \ces_4_0_io_ins_down[47] ,
    \ces_4_0_io_ins_down[46] ,
    \ces_4_0_io_ins_down[45] ,
    \ces_4_0_io_ins_down[44] ,
    \ces_4_0_io_ins_down[43] ,
    \ces_4_0_io_ins_down[42] ,
    \ces_4_0_io_ins_down[41] ,
    \ces_4_0_io_ins_down[40] ,
    \ces_4_0_io_ins_down[39] ,
    \ces_4_0_io_ins_down[38] ,
    \ces_4_0_io_ins_down[37] ,
    \ces_4_0_io_ins_down[36] ,
    \ces_4_0_io_ins_down[35] ,
    \ces_4_0_io_ins_down[34] ,
    \ces_4_0_io_ins_down[33] ,
    \ces_4_0_io_ins_down[32] ,
    \ces_4_0_io_ins_down[31] ,
    \ces_4_0_io_ins_down[30] ,
    \ces_4_0_io_ins_down[29] ,
    \ces_4_0_io_ins_down[28] ,
    \ces_4_0_io_ins_down[27] ,
    \ces_4_0_io_ins_down[26] ,
    \ces_4_0_io_ins_down[25] ,
    \ces_4_0_io_ins_down[24] ,
    \ces_4_0_io_ins_down[23] ,
    \ces_4_0_io_ins_down[22] ,
    \ces_4_0_io_ins_down[21] ,
    \ces_4_0_io_ins_down[20] ,
    \ces_4_0_io_ins_down[19] ,
    \ces_4_0_io_ins_down[18] ,
    \ces_4_0_io_ins_down[17] ,
    \ces_4_0_io_ins_down[16] ,
    \ces_4_0_io_ins_down[15] ,
    \ces_4_0_io_ins_down[14] ,
    \ces_4_0_io_ins_down[13] ,
    \ces_4_0_io_ins_down[12] ,
    \ces_4_0_io_ins_down[11] ,
    \ces_4_0_io_ins_down[10] ,
    \ces_4_0_io_ins_down[9] ,
    \ces_4_0_io_ins_down[8] ,
    \ces_4_0_io_ins_down[7] ,
    \ces_4_0_io_ins_down[6] ,
    \ces_4_0_io_ins_down[5] ,
    \ces_4_0_io_ins_down[4] ,
    \ces_4_0_io_ins_down[3] ,
    \ces_4_0_io_ins_down[2] ,
    \ces_4_0_io_ins_down[1] ,
    \ces_4_0_io_ins_down[0] }),
    .io_ins_left({\ces_4_0_io_ins_left[63] ,
    \ces_4_0_io_ins_left[62] ,
    \ces_4_0_io_ins_left[61] ,
    \ces_4_0_io_ins_left[60] ,
    \ces_4_0_io_ins_left[59] ,
    \ces_4_0_io_ins_left[58] ,
    \ces_4_0_io_ins_left[57] ,
    \ces_4_0_io_ins_left[56] ,
    \ces_4_0_io_ins_left[55] ,
    \ces_4_0_io_ins_left[54] ,
    \ces_4_0_io_ins_left[53] ,
    \ces_4_0_io_ins_left[52] ,
    \ces_4_0_io_ins_left[51] ,
    \ces_4_0_io_ins_left[50] ,
    \ces_4_0_io_ins_left[49] ,
    \ces_4_0_io_ins_left[48] ,
    \ces_4_0_io_ins_left[47] ,
    \ces_4_0_io_ins_left[46] ,
    \ces_4_0_io_ins_left[45] ,
    \ces_4_0_io_ins_left[44] ,
    \ces_4_0_io_ins_left[43] ,
    \ces_4_0_io_ins_left[42] ,
    \ces_4_0_io_ins_left[41] ,
    \ces_4_0_io_ins_left[40] ,
    \ces_4_0_io_ins_left[39] ,
    \ces_4_0_io_ins_left[38] ,
    \ces_4_0_io_ins_left[37] ,
    \ces_4_0_io_ins_left[36] ,
    \ces_4_0_io_ins_left[35] ,
    \ces_4_0_io_ins_left[34] ,
    \ces_4_0_io_ins_left[33] ,
    \ces_4_0_io_ins_left[32] ,
    \ces_4_0_io_ins_left[31] ,
    \ces_4_0_io_ins_left[30] ,
    \ces_4_0_io_ins_left[29] ,
    \ces_4_0_io_ins_left[28] ,
    \ces_4_0_io_ins_left[27] ,
    \ces_4_0_io_ins_left[26] ,
    \ces_4_0_io_ins_left[25] ,
    \ces_4_0_io_ins_left[24] ,
    \ces_4_0_io_ins_left[23] ,
    \ces_4_0_io_ins_left[22] ,
    \ces_4_0_io_ins_left[21] ,
    \ces_4_0_io_ins_left[20] ,
    \ces_4_0_io_ins_left[19] ,
    \ces_4_0_io_ins_left[18] ,
    \ces_4_0_io_ins_left[17] ,
    \ces_4_0_io_ins_left[16] ,
    \ces_4_0_io_ins_left[15] ,
    \ces_4_0_io_ins_left[14] ,
    \ces_4_0_io_ins_left[13] ,
    \ces_4_0_io_ins_left[12] ,
    \ces_4_0_io_ins_left[11] ,
    \ces_4_0_io_ins_left[10] ,
    \ces_4_0_io_ins_left[9] ,
    \ces_4_0_io_ins_left[8] ,
    \ces_4_0_io_ins_left[7] ,
    \ces_4_0_io_ins_left[6] ,
    \ces_4_0_io_ins_left[5] ,
    \ces_4_0_io_ins_left[4] ,
    \ces_4_0_io_ins_left[3] ,
    \ces_4_0_io_ins_left[2] ,
    \ces_4_0_io_ins_left[1] ,
    \ces_4_0_io_ins_left[0] }),
    .io_ins_right({net1340,
    net1339,
    net1338,
    net1337,
    net1335,
    net1334,
    net1333,
    net1332,
    net1331,
    net1330,
    net1329,
    net1328,
    net1327,
    net1326,
    net1324,
    net1323,
    net1322,
    net1321,
    net1320,
    net1319,
    net1318,
    net1317,
    net1316,
    net1315,
    net1313,
    net1312,
    net1311,
    net1310,
    net1309,
    net1308,
    net1307,
    net1306,
    net1305,
    net1304,
    net1302,
    net1301,
    net1300,
    net1299,
    net1298,
    net1297,
    net1296,
    net1295,
    net1294,
    net1293,
    net1291,
    net1290,
    net1289,
    net1288,
    net1287,
    net1286,
    net1285,
    net1284,
    net1283,
    net1282,
    net1344,
    net1343,
    net1342,
    net1341,
    net1336,
    net1325,
    net1314,
    net1303,
    net1292,
    net1281}),
    .io_ins_up({\ces_3_0_io_outs_up[63] ,
    \ces_3_0_io_outs_up[62] ,
    \ces_3_0_io_outs_up[61] ,
    \ces_3_0_io_outs_up[60] ,
    \ces_3_0_io_outs_up[59] ,
    \ces_3_0_io_outs_up[58] ,
    \ces_3_0_io_outs_up[57] ,
    \ces_3_0_io_outs_up[56] ,
    \ces_3_0_io_outs_up[55] ,
    \ces_3_0_io_outs_up[54] ,
    \ces_3_0_io_outs_up[53] ,
    \ces_3_0_io_outs_up[52] ,
    \ces_3_0_io_outs_up[51] ,
    \ces_3_0_io_outs_up[50] ,
    \ces_3_0_io_outs_up[49] ,
    \ces_3_0_io_outs_up[48] ,
    \ces_3_0_io_outs_up[47] ,
    \ces_3_0_io_outs_up[46] ,
    \ces_3_0_io_outs_up[45] ,
    \ces_3_0_io_outs_up[44] ,
    \ces_3_0_io_outs_up[43] ,
    \ces_3_0_io_outs_up[42] ,
    \ces_3_0_io_outs_up[41] ,
    \ces_3_0_io_outs_up[40] ,
    \ces_3_0_io_outs_up[39] ,
    \ces_3_0_io_outs_up[38] ,
    \ces_3_0_io_outs_up[37] ,
    \ces_3_0_io_outs_up[36] ,
    \ces_3_0_io_outs_up[35] ,
    \ces_3_0_io_outs_up[34] ,
    \ces_3_0_io_outs_up[33] ,
    \ces_3_0_io_outs_up[32] ,
    \ces_3_0_io_outs_up[31] ,
    \ces_3_0_io_outs_up[30] ,
    \ces_3_0_io_outs_up[29] ,
    \ces_3_0_io_outs_up[28] ,
    \ces_3_0_io_outs_up[27] ,
    \ces_3_0_io_outs_up[26] ,
    \ces_3_0_io_outs_up[25] ,
    \ces_3_0_io_outs_up[24] ,
    \ces_3_0_io_outs_up[23] ,
    \ces_3_0_io_outs_up[22] ,
    \ces_3_0_io_outs_up[21] ,
    \ces_3_0_io_outs_up[20] ,
    \ces_3_0_io_outs_up[19] ,
    \ces_3_0_io_outs_up[18] ,
    \ces_3_0_io_outs_up[17] ,
    \ces_3_0_io_outs_up[16] ,
    \ces_3_0_io_outs_up[15] ,
    \ces_3_0_io_outs_up[14] ,
    \ces_3_0_io_outs_up[13] ,
    \ces_3_0_io_outs_up[12] ,
    \ces_3_0_io_outs_up[11] ,
    \ces_3_0_io_outs_up[10] ,
    \ces_3_0_io_outs_up[9] ,
    \ces_3_0_io_outs_up[8] ,
    \ces_3_0_io_outs_up[7] ,
    \ces_3_0_io_outs_up[6] ,
    \ces_3_0_io_outs_up[5] ,
    \ces_3_0_io_outs_up[4] ,
    \ces_3_0_io_outs_up[3] ,
    \ces_3_0_io_outs_up[2] ,
    \ces_3_0_io_outs_up[1] ,
    \ces_3_0_io_outs_up[0] }),
    .io_outs_down({\ces_3_0_io_ins_down[63] ,
    \ces_3_0_io_ins_down[62] ,
    \ces_3_0_io_ins_down[61] ,
    \ces_3_0_io_ins_down[60] ,
    \ces_3_0_io_ins_down[59] ,
    \ces_3_0_io_ins_down[58] ,
    \ces_3_0_io_ins_down[57] ,
    \ces_3_0_io_ins_down[56] ,
    \ces_3_0_io_ins_down[55] ,
    \ces_3_0_io_ins_down[54] ,
    \ces_3_0_io_ins_down[53] ,
    \ces_3_0_io_ins_down[52] ,
    \ces_3_0_io_ins_down[51] ,
    \ces_3_0_io_ins_down[50] ,
    \ces_3_0_io_ins_down[49] ,
    \ces_3_0_io_ins_down[48] ,
    \ces_3_0_io_ins_down[47] ,
    \ces_3_0_io_ins_down[46] ,
    \ces_3_0_io_ins_down[45] ,
    \ces_3_0_io_ins_down[44] ,
    \ces_3_0_io_ins_down[43] ,
    \ces_3_0_io_ins_down[42] ,
    \ces_3_0_io_ins_down[41] ,
    \ces_3_0_io_ins_down[40] ,
    \ces_3_0_io_ins_down[39] ,
    \ces_3_0_io_ins_down[38] ,
    \ces_3_0_io_ins_down[37] ,
    \ces_3_0_io_ins_down[36] ,
    \ces_3_0_io_ins_down[35] ,
    \ces_3_0_io_ins_down[34] ,
    \ces_3_0_io_ins_down[33] ,
    \ces_3_0_io_ins_down[32] ,
    \ces_3_0_io_ins_down[31] ,
    \ces_3_0_io_ins_down[30] ,
    \ces_3_0_io_ins_down[29] ,
    \ces_3_0_io_ins_down[28] ,
    \ces_3_0_io_ins_down[27] ,
    \ces_3_0_io_ins_down[26] ,
    \ces_3_0_io_ins_down[25] ,
    \ces_3_0_io_ins_down[24] ,
    \ces_3_0_io_ins_down[23] ,
    \ces_3_0_io_ins_down[22] ,
    \ces_3_0_io_ins_down[21] ,
    \ces_3_0_io_ins_down[20] ,
    \ces_3_0_io_ins_down[19] ,
    \ces_3_0_io_ins_down[18] ,
    \ces_3_0_io_ins_down[17] ,
    \ces_3_0_io_ins_down[16] ,
    \ces_3_0_io_ins_down[15] ,
    \ces_3_0_io_ins_down[14] ,
    \ces_3_0_io_ins_down[13] ,
    \ces_3_0_io_ins_down[12] ,
    \ces_3_0_io_ins_down[11] ,
    \ces_3_0_io_ins_down[10] ,
    \ces_3_0_io_ins_down[9] ,
    \ces_3_0_io_ins_down[8] ,
    \ces_3_0_io_ins_down[7] ,
    \ces_3_0_io_ins_down[6] ,
    \ces_3_0_io_ins_down[5] ,
    \ces_3_0_io_ins_down[4] ,
    \ces_3_0_io_ins_down[3] ,
    \ces_3_0_io_ins_down[2] ,
    \ces_3_0_io_ins_down[1] ,
    \ces_3_0_io_ins_down[0] }),
    .io_outs_left({net2940,
    net2939,
    net2938,
    net2937,
    net2935,
    net2934,
    net2933,
    net2932,
    net2931,
    net2930,
    net2929,
    net2928,
    net2927,
    net2926,
    net2924,
    net2923,
    net2922,
    net2921,
    net2920,
    net2919,
    net2918,
    net2917,
    net2916,
    net2915,
    net2913,
    net2912,
    net2911,
    net2910,
    net2909,
    net2908,
    net2907,
    net2906,
    net2905,
    net2904,
    net2902,
    net2901,
    net2900,
    net2899,
    net2898,
    net2897,
    net2896,
    net2895,
    net2894,
    net2893,
    net2891,
    net2890,
    net2889,
    net2888,
    net2887,
    net2886,
    net2885,
    net2884,
    net2883,
    net2882,
    net2944,
    net2943,
    net2942,
    net2941,
    net2936,
    net2925,
    net2914,
    net2903,
    net2892,
    net2881}),
    .io_outs_right({\ces_4_0_io_outs_right[63] ,
    \ces_4_0_io_outs_right[62] ,
    \ces_4_0_io_outs_right[61] ,
    \ces_4_0_io_outs_right[60] ,
    \ces_4_0_io_outs_right[59] ,
    \ces_4_0_io_outs_right[58] ,
    \ces_4_0_io_outs_right[57] ,
    \ces_4_0_io_outs_right[56] ,
    \ces_4_0_io_outs_right[55] ,
    \ces_4_0_io_outs_right[54] ,
    \ces_4_0_io_outs_right[53] ,
    \ces_4_0_io_outs_right[52] ,
    \ces_4_0_io_outs_right[51] ,
    \ces_4_0_io_outs_right[50] ,
    \ces_4_0_io_outs_right[49] ,
    \ces_4_0_io_outs_right[48] ,
    \ces_4_0_io_outs_right[47] ,
    \ces_4_0_io_outs_right[46] ,
    \ces_4_0_io_outs_right[45] ,
    \ces_4_0_io_outs_right[44] ,
    \ces_4_0_io_outs_right[43] ,
    \ces_4_0_io_outs_right[42] ,
    \ces_4_0_io_outs_right[41] ,
    \ces_4_0_io_outs_right[40] ,
    \ces_4_0_io_outs_right[39] ,
    \ces_4_0_io_outs_right[38] ,
    \ces_4_0_io_outs_right[37] ,
    \ces_4_0_io_outs_right[36] ,
    \ces_4_0_io_outs_right[35] ,
    \ces_4_0_io_outs_right[34] ,
    \ces_4_0_io_outs_right[33] ,
    \ces_4_0_io_outs_right[32] ,
    \ces_4_0_io_outs_right[31] ,
    \ces_4_0_io_outs_right[30] ,
    \ces_4_0_io_outs_right[29] ,
    \ces_4_0_io_outs_right[28] ,
    \ces_4_0_io_outs_right[27] ,
    \ces_4_0_io_outs_right[26] ,
    \ces_4_0_io_outs_right[25] ,
    \ces_4_0_io_outs_right[24] ,
    \ces_4_0_io_outs_right[23] ,
    \ces_4_0_io_outs_right[22] ,
    \ces_4_0_io_outs_right[21] ,
    \ces_4_0_io_outs_right[20] ,
    \ces_4_0_io_outs_right[19] ,
    \ces_4_0_io_outs_right[18] ,
    \ces_4_0_io_outs_right[17] ,
    \ces_4_0_io_outs_right[16] ,
    \ces_4_0_io_outs_right[15] ,
    \ces_4_0_io_outs_right[14] ,
    \ces_4_0_io_outs_right[13] ,
    \ces_4_0_io_outs_right[12] ,
    \ces_4_0_io_outs_right[11] ,
    \ces_4_0_io_outs_right[10] ,
    \ces_4_0_io_outs_right[9] ,
    \ces_4_0_io_outs_right[8] ,
    \ces_4_0_io_outs_right[7] ,
    \ces_4_0_io_outs_right[6] ,
    \ces_4_0_io_outs_right[5] ,
    \ces_4_0_io_outs_right[4] ,
    \ces_4_0_io_outs_right[3] ,
    \ces_4_0_io_outs_right[2] ,
    \ces_4_0_io_outs_right[1] ,
    \ces_4_0_io_outs_right[0] }),
    .io_outs_up({\ces_4_0_io_outs_up[63] ,
    \ces_4_0_io_outs_up[62] ,
    \ces_4_0_io_outs_up[61] ,
    \ces_4_0_io_outs_up[60] ,
    \ces_4_0_io_outs_up[59] ,
    \ces_4_0_io_outs_up[58] ,
    \ces_4_0_io_outs_up[57] ,
    \ces_4_0_io_outs_up[56] ,
    \ces_4_0_io_outs_up[55] ,
    \ces_4_0_io_outs_up[54] ,
    \ces_4_0_io_outs_up[53] ,
    \ces_4_0_io_outs_up[52] ,
    \ces_4_0_io_outs_up[51] ,
    \ces_4_0_io_outs_up[50] ,
    \ces_4_0_io_outs_up[49] ,
    \ces_4_0_io_outs_up[48] ,
    \ces_4_0_io_outs_up[47] ,
    \ces_4_0_io_outs_up[46] ,
    \ces_4_0_io_outs_up[45] ,
    \ces_4_0_io_outs_up[44] ,
    \ces_4_0_io_outs_up[43] ,
    \ces_4_0_io_outs_up[42] ,
    \ces_4_0_io_outs_up[41] ,
    \ces_4_0_io_outs_up[40] ,
    \ces_4_0_io_outs_up[39] ,
    \ces_4_0_io_outs_up[38] ,
    \ces_4_0_io_outs_up[37] ,
    \ces_4_0_io_outs_up[36] ,
    \ces_4_0_io_outs_up[35] ,
    \ces_4_0_io_outs_up[34] ,
    \ces_4_0_io_outs_up[33] ,
    \ces_4_0_io_outs_up[32] ,
    \ces_4_0_io_outs_up[31] ,
    \ces_4_0_io_outs_up[30] ,
    \ces_4_0_io_outs_up[29] ,
    \ces_4_0_io_outs_up[28] ,
    \ces_4_0_io_outs_up[27] ,
    \ces_4_0_io_outs_up[26] ,
    \ces_4_0_io_outs_up[25] ,
    \ces_4_0_io_outs_up[24] ,
    \ces_4_0_io_outs_up[23] ,
    \ces_4_0_io_outs_up[22] ,
    \ces_4_0_io_outs_up[21] ,
    \ces_4_0_io_outs_up[20] ,
    \ces_4_0_io_outs_up[19] ,
    \ces_4_0_io_outs_up[18] ,
    \ces_4_0_io_outs_up[17] ,
    \ces_4_0_io_outs_up[16] ,
    \ces_4_0_io_outs_up[15] ,
    \ces_4_0_io_outs_up[14] ,
    \ces_4_0_io_outs_up[13] ,
    \ces_4_0_io_outs_up[12] ,
    \ces_4_0_io_outs_up[11] ,
    \ces_4_0_io_outs_up[10] ,
    \ces_4_0_io_outs_up[9] ,
    \ces_4_0_io_outs_up[8] ,
    \ces_4_0_io_outs_up[7] ,
    \ces_4_0_io_outs_up[6] ,
    \ces_4_0_io_outs_up[5] ,
    \ces_4_0_io_outs_up[4] ,
    \ces_4_0_io_outs_up[3] ,
    \ces_4_0_io_outs_up[2] ,
    \ces_4_0_io_outs_up[1] ,
    \ces_4_0_io_outs_up[0] }));
 Element ces_4_1 (.clock(clknet_3_4_0_clock),
    .io_lsbIns_1(ces_4_0_io_lsbOuts_1),
    .io_lsbIns_2(ces_4_0_io_lsbOuts_2),
    .io_lsbIns_3(ces_4_0_io_lsbOuts_3),
    .io_lsbIns_4(ces_4_0_io_lsbOuts_4),
    .io_lsbIns_5(ces_4_0_io_lsbOuts_5),
    .io_lsbIns_6(ces_4_0_io_lsbOuts_6),
    .io_lsbIns_7(ces_4_0_io_lsbOuts_7),
    .io_lsbOuts_0(ces_4_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_1_io_lsbOuts_7),
    .io_ins_down({\ces_4_1_io_ins_down[63] ,
    \ces_4_1_io_ins_down[62] ,
    \ces_4_1_io_ins_down[61] ,
    \ces_4_1_io_ins_down[60] ,
    \ces_4_1_io_ins_down[59] ,
    \ces_4_1_io_ins_down[58] ,
    \ces_4_1_io_ins_down[57] ,
    \ces_4_1_io_ins_down[56] ,
    \ces_4_1_io_ins_down[55] ,
    \ces_4_1_io_ins_down[54] ,
    \ces_4_1_io_ins_down[53] ,
    \ces_4_1_io_ins_down[52] ,
    \ces_4_1_io_ins_down[51] ,
    \ces_4_1_io_ins_down[50] ,
    \ces_4_1_io_ins_down[49] ,
    \ces_4_1_io_ins_down[48] ,
    \ces_4_1_io_ins_down[47] ,
    \ces_4_1_io_ins_down[46] ,
    \ces_4_1_io_ins_down[45] ,
    \ces_4_1_io_ins_down[44] ,
    \ces_4_1_io_ins_down[43] ,
    \ces_4_1_io_ins_down[42] ,
    \ces_4_1_io_ins_down[41] ,
    \ces_4_1_io_ins_down[40] ,
    \ces_4_1_io_ins_down[39] ,
    \ces_4_1_io_ins_down[38] ,
    \ces_4_1_io_ins_down[37] ,
    \ces_4_1_io_ins_down[36] ,
    \ces_4_1_io_ins_down[35] ,
    \ces_4_1_io_ins_down[34] ,
    \ces_4_1_io_ins_down[33] ,
    \ces_4_1_io_ins_down[32] ,
    \ces_4_1_io_ins_down[31] ,
    \ces_4_1_io_ins_down[30] ,
    \ces_4_1_io_ins_down[29] ,
    \ces_4_1_io_ins_down[28] ,
    \ces_4_1_io_ins_down[27] ,
    \ces_4_1_io_ins_down[26] ,
    \ces_4_1_io_ins_down[25] ,
    \ces_4_1_io_ins_down[24] ,
    \ces_4_1_io_ins_down[23] ,
    \ces_4_1_io_ins_down[22] ,
    \ces_4_1_io_ins_down[21] ,
    \ces_4_1_io_ins_down[20] ,
    \ces_4_1_io_ins_down[19] ,
    \ces_4_1_io_ins_down[18] ,
    \ces_4_1_io_ins_down[17] ,
    \ces_4_1_io_ins_down[16] ,
    \ces_4_1_io_ins_down[15] ,
    \ces_4_1_io_ins_down[14] ,
    \ces_4_1_io_ins_down[13] ,
    \ces_4_1_io_ins_down[12] ,
    \ces_4_1_io_ins_down[11] ,
    \ces_4_1_io_ins_down[10] ,
    \ces_4_1_io_ins_down[9] ,
    \ces_4_1_io_ins_down[8] ,
    \ces_4_1_io_ins_down[7] ,
    \ces_4_1_io_ins_down[6] ,
    \ces_4_1_io_ins_down[5] ,
    \ces_4_1_io_ins_down[4] ,
    \ces_4_1_io_ins_down[3] ,
    \ces_4_1_io_ins_down[2] ,
    \ces_4_1_io_ins_down[1] ,
    \ces_4_1_io_ins_down[0] }),
    .io_ins_left({\ces_4_1_io_ins_left[63] ,
    \ces_4_1_io_ins_left[62] ,
    \ces_4_1_io_ins_left[61] ,
    \ces_4_1_io_ins_left[60] ,
    \ces_4_1_io_ins_left[59] ,
    \ces_4_1_io_ins_left[58] ,
    \ces_4_1_io_ins_left[57] ,
    \ces_4_1_io_ins_left[56] ,
    \ces_4_1_io_ins_left[55] ,
    \ces_4_1_io_ins_left[54] ,
    \ces_4_1_io_ins_left[53] ,
    \ces_4_1_io_ins_left[52] ,
    \ces_4_1_io_ins_left[51] ,
    \ces_4_1_io_ins_left[50] ,
    \ces_4_1_io_ins_left[49] ,
    \ces_4_1_io_ins_left[48] ,
    \ces_4_1_io_ins_left[47] ,
    \ces_4_1_io_ins_left[46] ,
    \ces_4_1_io_ins_left[45] ,
    \ces_4_1_io_ins_left[44] ,
    \ces_4_1_io_ins_left[43] ,
    \ces_4_1_io_ins_left[42] ,
    \ces_4_1_io_ins_left[41] ,
    \ces_4_1_io_ins_left[40] ,
    \ces_4_1_io_ins_left[39] ,
    \ces_4_1_io_ins_left[38] ,
    \ces_4_1_io_ins_left[37] ,
    \ces_4_1_io_ins_left[36] ,
    \ces_4_1_io_ins_left[35] ,
    \ces_4_1_io_ins_left[34] ,
    \ces_4_1_io_ins_left[33] ,
    \ces_4_1_io_ins_left[32] ,
    \ces_4_1_io_ins_left[31] ,
    \ces_4_1_io_ins_left[30] ,
    \ces_4_1_io_ins_left[29] ,
    \ces_4_1_io_ins_left[28] ,
    \ces_4_1_io_ins_left[27] ,
    \ces_4_1_io_ins_left[26] ,
    \ces_4_1_io_ins_left[25] ,
    \ces_4_1_io_ins_left[24] ,
    \ces_4_1_io_ins_left[23] ,
    \ces_4_1_io_ins_left[22] ,
    \ces_4_1_io_ins_left[21] ,
    \ces_4_1_io_ins_left[20] ,
    \ces_4_1_io_ins_left[19] ,
    \ces_4_1_io_ins_left[18] ,
    \ces_4_1_io_ins_left[17] ,
    \ces_4_1_io_ins_left[16] ,
    \ces_4_1_io_ins_left[15] ,
    \ces_4_1_io_ins_left[14] ,
    \ces_4_1_io_ins_left[13] ,
    \ces_4_1_io_ins_left[12] ,
    \ces_4_1_io_ins_left[11] ,
    \ces_4_1_io_ins_left[10] ,
    \ces_4_1_io_ins_left[9] ,
    \ces_4_1_io_ins_left[8] ,
    \ces_4_1_io_ins_left[7] ,
    \ces_4_1_io_ins_left[6] ,
    \ces_4_1_io_ins_left[5] ,
    \ces_4_1_io_ins_left[4] ,
    \ces_4_1_io_ins_left[3] ,
    \ces_4_1_io_ins_left[2] ,
    \ces_4_1_io_ins_left[1] ,
    \ces_4_1_io_ins_left[0] }),
    .io_ins_right({\ces_4_0_io_outs_right[63] ,
    \ces_4_0_io_outs_right[62] ,
    \ces_4_0_io_outs_right[61] ,
    \ces_4_0_io_outs_right[60] ,
    \ces_4_0_io_outs_right[59] ,
    \ces_4_0_io_outs_right[58] ,
    \ces_4_0_io_outs_right[57] ,
    \ces_4_0_io_outs_right[56] ,
    \ces_4_0_io_outs_right[55] ,
    \ces_4_0_io_outs_right[54] ,
    \ces_4_0_io_outs_right[53] ,
    \ces_4_0_io_outs_right[52] ,
    \ces_4_0_io_outs_right[51] ,
    \ces_4_0_io_outs_right[50] ,
    \ces_4_0_io_outs_right[49] ,
    \ces_4_0_io_outs_right[48] ,
    \ces_4_0_io_outs_right[47] ,
    \ces_4_0_io_outs_right[46] ,
    \ces_4_0_io_outs_right[45] ,
    \ces_4_0_io_outs_right[44] ,
    \ces_4_0_io_outs_right[43] ,
    \ces_4_0_io_outs_right[42] ,
    \ces_4_0_io_outs_right[41] ,
    \ces_4_0_io_outs_right[40] ,
    \ces_4_0_io_outs_right[39] ,
    \ces_4_0_io_outs_right[38] ,
    \ces_4_0_io_outs_right[37] ,
    \ces_4_0_io_outs_right[36] ,
    \ces_4_0_io_outs_right[35] ,
    \ces_4_0_io_outs_right[34] ,
    \ces_4_0_io_outs_right[33] ,
    \ces_4_0_io_outs_right[32] ,
    \ces_4_0_io_outs_right[31] ,
    \ces_4_0_io_outs_right[30] ,
    \ces_4_0_io_outs_right[29] ,
    \ces_4_0_io_outs_right[28] ,
    \ces_4_0_io_outs_right[27] ,
    \ces_4_0_io_outs_right[26] ,
    \ces_4_0_io_outs_right[25] ,
    \ces_4_0_io_outs_right[24] ,
    \ces_4_0_io_outs_right[23] ,
    \ces_4_0_io_outs_right[22] ,
    \ces_4_0_io_outs_right[21] ,
    \ces_4_0_io_outs_right[20] ,
    \ces_4_0_io_outs_right[19] ,
    \ces_4_0_io_outs_right[18] ,
    \ces_4_0_io_outs_right[17] ,
    \ces_4_0_io_outs_right[16] ,
    \ces_4_0_io_outs_right[15] ,
    \ces_4_0_io_outs_right[14] ,
    \ces_4_0_io_outs_right[13] ,
    \ces_4_0_io_outs_right[12] ,
    \ces_4_0_io_outs_right[11] ,
    \ces_4_0_io_outs_right[10] ,
    \ces_4_0_io_outs_right[9] ,
    \ces_4_0_io_outs_right[8] ,
    \ces_4_0_io_outs_right[7] ,
    \ces_4_0_io_outs_right[6] ,
    \ces_4_0_io_outs_right[5] ,
    \ces_4_0_io_outs_right[4] ,
    \ces_4_0_io_outs_right[3] ,
    \ces_4_0_io_outs_right[2] ,
    \ces_4_0_io_outs_right[1] ,
    \ces_4_0_io_outs_right[0] }),
    .io_ins_up({\ces_3_1_io_outs_up[63] ,
    \ces_3_1_io_outs_up[62] ,
    \ces_3_1_io_outs_up[61] ,
    \ces_3_1_io_outs_up[60] ,
    \ces_3_1_io_outs_up[59] ,
    \ces_3_1_io_outs_up[58] ,
    \ces_3_1_io_outs_up[57] ,
    \ces_3_1_io_outs_up[56] ,
    \ces_3_1_io_outs_up[55] ,
    \ces_3_1_io_outs_up[54] ,
    \ces_3_1_io_outs_up[53] ,
    \ces_3_1_io_outs_up[52] ,
    \ces_3_1_io_outs_up[51] ,
    \ces_3_1_io_outs_up[50] ,
    \ces_3_1_io_outs_up[49] ,
    \ces_3_1_io_outs_up[48] ,
    \ces_3_1_io_outs_up[47] ,
    \ces_3_1_io_outs_up[46] ,
    \ces_3_1_io_outs_up[45] ,
    \ces_3_1_io_outs_up[44] ,
    \ces_3_1_io_outs_up[43] ,
    \ces_3_1_io_outs_up[42] ,
    \ces_3_1_io_outs_up[41] ,
    \ces_3_1_io_outs_up[40] ,
    \ces_3_1_io_outs_up[39] ,
    \ces_3_1_io_outs_up[38] ,
    \ces_3_1_io_outs_up[37] ,
    \ces_3_1_io_outs_up[36] ,
    \ces_3_1_io_outs_up[35] ,
    \ces_3_1_io_outs_up[34] ,
    \ces_3_1_io_outs_up[33] ,
    \ces_3_1_io_outs_up[32] ,
    \ces_3_1_io_outs_up[31] ,
    \ces_3_1_io_outs_up[30] ,
    \ces_3_1_io_outs_up[29] ,
    \ces_3_1_io_outs_up[28] ,
    \ces_3_1_io_outs_up[27] ,
    \ces_3_1_io_outs_up[26] ,
    \ces_3_1_io_outs_up[25] ,
    \ces_3_1_io_outs_up[24] ,
    \ces_3_1_io_outs_up[23] ,
    \ces_3_1_io_outs_up[22] ,
    \ces_3_1_io_outs_up[21] ,
    \ces_3_1_io_outs_up[20] ,
    \ces_3_1_io_outs_up[19] ,
    \ces_3_1_io_outs_up[18] ,
    \ces_3_1_io_outs_up[17] ,
    \ces_3_1_io_outs_up[16] ,
    \ces_3_1_io_outs_up[15] ,
    \ces_3_1_io_outs_up[14] ,
    \ces_3_1_io_outs_up[13] ,
    \ces_3_1_io_outs_up[12] ,
    \ces_3_1_io_outs_up[11] ,
    \ces_3_1_io_outs_up[10] ,
    \ces_3_1_io_outs_up[9] ,
    \ces_3_1_io_outs_up[8] ,
    \ces_3_1_io_outs_up[7] ,
    \ces_3_1_io_outs_up[6] ,
    \ces_3_1_io_outs_up[5] ,
    \ces_3_1_io_outs_up[4] ,
    \ces_3_1_io_outs_up[3] ,
    \ces_3_1_io_outs_up[2] ,
    \ces_3_1_io_outs_up[1] ,
    \ces_3_1_io_outs_up[0] }),
    .io_outs_down({\ces_3_1_io_ins_down[63] ,
    \ces_3_1_io_ins_down[62] ,
    \ces_3_1_io_ins_down[61] ,
    \ces_3_1_io_ins_down[60] ,
    \ces_3_1_io_ins_down[59] ,
    \ces_3_1_io_ins_down[58] ,
    \ces_3_1_io_ins_down[57] ,
    \ces_3_1_io_ins_down[56] ,
    \ces_3_1_io_ins_down[55] ,
    \ces_3_1_io_ins_down[54] ,
    \ces_3_1_io_ins_down[53] ,
    \ces_3_1_io_ins_down[52] ,
    \ces_3_1_io_ins_down[51] ,
    \ces_3_1_io_ins_down[50] ,
    \ces_3_1_io_ins_down[49] ,
    \ces_3_1_io_ins_down[48] ,
    \ces_3_1_io_ins_down[47] ,
    \ces_3_1_io_ins_down[46] ,
    \ces_3_1_io_ins_down[45] ,
    \ces_3_1_io_ins_down[44] ,
    \ces_3_1_io_ins_down[43] ,
    \ces_3_1_io_ins_down[42] ,
    \ces_3_1_io_ins_down[41] ,
    \ces_3_1_io_ins_down[40] ,
    \ces_3_1_io_ins_down[39] ,
    \ces_3_1_io_ins_down[38] ,
    \ces_3_1_io_ins_down[37] ,
    \ces_3_1_io_ins_down[36] ,
    \ces_3_1_io_ins_down[35] ,
    \ces_3_1_io_ins_down[34] ,
    \ces_3_1_io_ins_down[33] ,
    \ces_3_1_io_ins_down[32] ,
    \ces_3_1_io_ins_down[31] ,
    \ces_3_1_io_ins_down[30] ,
    \ces_3_1_io_ins_down[29] ,
    \ces_3_1_io_ins_down[28] ,
    \ces_3_1_io_ins_down[27] ,
    \ces_3_1_io_ins_down[26] ,
    \ces_3_1_io_ins_down[25] ,
    \ces_3_1_io_ins_down[24] ,
    \ces_3_1_io_ins_down[23] ,
    \ces_3_1_io_ins_down[22] ,
    \ces_3_1_io_ins_down[21] ,
    \ces_3_1_io_ins_down[20] ,
    \ces_3_1_io_ins_down[19] ,
    \ces_3_1_io_ins_down[18] ,
    \ces_3_1_io_ins_down[17] ,
    \ces_3_1_io_ins_down[16] ,
    \ces_3_1_io_ins_down[15] ,
    \ces_3_1_io_ins_down[14] ,
    \ces_3_1_io_ins_down[13] ,
    \ces_3_1_io_ins_down[12] ,
    \ces_3_1_io_ins_down[11] ,
    \ces_3_1_io_ins_down[10] ,
    \ces_3_1_io_ins_down[9] ,
    \ces_3_1_io_ins_down[8] ,
    \ces_3_1_io_ins_down[7] ,
    \ces_3_1_io_ins_down[6] ,
    \ces_3_1_io_ins_down[5] ,
    \ces_3_1_io_ins_down[4] ,
    \ces_3_1_io_ins_down[3] ,
    \ces_3_1_io_ins_down[2] ,
    \ces_3_1_io_ins_down[1] ,
    \ces_3_1_io_ins_down[0] }),
    .io_outs_left({\ces_4_0_io_ins_left[63] ,
    \ces_4_0_io_ins_left[62] ,
    \ces_4_0_io_ins_left[61] ,
    \ces_4_0_io_ins_left[60] ,
    \ces_4_0_io_ins_left[59] ,
    \ces_4_0_io_ins_left[58] ,
    \ces_4_0_io_ins_left[57] ,
    \ces_4_0_io_ins_left[56] ,
    \ces_4_0_io_ins_left[55] ,
    \ces_4_0_io_ins_left[54] ,
    \ces_4_0_io_ins_left[53] ,
    \ces_4_0_io_ins_left[52] ,
    \ces_4_0_io_ins_left[51] ,
    \ces_4_0_io_ins_left[50] ,
    \ces_4_0_io_ins_left[49] ,
    \ces_4_0_io_ins_left[48] ,
    \ces_4_0_io_ins_left[47] ,
    \ces_4_0_io_ins_left[46] ,
    \ces_4_0_io_ins_left[45] ,
    \ces_4_0_io_ins_left[44] ,
    \ces_4_0_io_ins_left[43] ,
    \ces_4_0_io_ins_left[42] ,
    \ces_4_0_io_ins_left[41] ,
    \ces_4_0_io_ins_left[40] ,
    \ces_4_0_io_ins_left[39] ,
    \ces_4_0_io_ins_left[38] ,
    \ces_4_0_io_ins_left[37] ,
    \ces_4_0_io_ins_left[36] ,
    \ces_4_0_io_ins_left[35] ,
    \ces_4_0_io_ins_left[34] ,
    \ces_4_0_io_ins_left[33] ,
    \ces_4_0_io_ins_left[32] ,
    \ces_4_0_io_ins_left[31] ,
    \ces_4_0_io_ins_left[30] ,
    \ces_4_0_io_ins_left[29] ,
    \ces_4_0_io_ins_left[28] ,
    \ces_4_0_io_ins_left[27] ,
    \ces_4_0_io_ins_left[26] ,
    \ces_4_0_io_ins_left[25] ,
    \ces_4_0_io_ins_left[24] ,
    \ces_4_0_io_ins_left[23] ,
    \ces_4_0_io_ins_left[22] ,
    \ces_4_0_io_ins_left[21] ,
    \ces_4_0_io_ins_left[20] ,
    \ces_4_0_io_ins_left[19] ,
    \ces_4_0_io_ins_left[18] ,
    \ces_4_0_io_ins_left[17] ,
    \ces_4_0_io_ins_left[16] ,
    \ces_4_0_io_ins_left[15] ,
    \ces_4_0_io_ins_left[14] ,
    \ces_4_0_io_ins_left[13] ,
    \ces_4_0_io_ins_left[12] ,
    \ces_4_0_io_ins_left[11] ,
    \ces_4_0_io_ins_left[10] ,
    \ces_4_0_io_ins_left[9] ,
    \ces_4_0_io_ins_left[8] ,
    \ces_4_0_io_ins_left[7] ,
    \ces_4_0_io_ins_left[6] ,
    \ces_4_0_io_ins_left[5] ,
    \ces_4_0_io_ins_left[4] ,
    \ces_4_0_io_ins_left[3] ,
    \ces_4_0_io_ins_left[2] ,
    \ces_4_0_io_ins_left[1] ,
    \ces_4_0_io_ins_left[0] }),
    .io_outs_right({\ces_4_1_io_outs_right[63] ,
    \ces_4_1_io_outs_right[62] ,
    \ces_4_1_io_outs_right[61] ,
    \ces_4_1_io_outs_right[60] ,
    \ces_4_1_io_outs_right[59] ,
    \ces_4_1_io_outs_right[58] ,
    \ces_4_1_io_outs_right[57] ,
    \ces_4_1_io_outs_right[56] ,
    \ces_4_1_io_outs_right[55] ,
    \ces_4_1_io_outs_right[54] ,
    \ces_4_1_io_outs_right[53] ,
    \ces_4_1_io_outs_right[52] ,
    \ces_4_1_io_outs_right[51] ,
    \ces_4_1_io_outs_right[50] ,
    \ces_4_1_io_outs_right[49] ,
    \ces_4_1_io_outs_right[48] ,
    \ces_4_1_io_outs_right[47] ,
    \ces_4_1_io_outs_right[46] ,
    \ces_4_1_io_outs_right[45] ,
    \ces_4_1_io_outs_right[44] ,
    \ces_4_1_io_outs_right[43] ,
    \ces_4_1_io_outs_right[42] ,
    \ces_4_1_io_outs_right[41] ,
    \ces_4_1_io_outs_right[40] ,
    \ces_4_1_io_outs_right[39] ,
    \ces_4_1_io_outs_right[38] ,
    \ces_4_1_io_outs_right[37] ,
    \ces_4_1_io_outs_right[36] ,
    \ces_4_1_io_outs_right[35] ,
    \ces_4_1_io_outs_right[34] ,
    \ces_4_1_io_outs_right[33] ,
    \ces_4_1_io_outs_right[32] ,
    \ces_4_1_io_outs_right[31] ,
    \ces_4_1_io_outs_right[30] ,
    \ces_4_1_io_outs_right[29] ,
    \ces_4_1_io_outs_right[28] ,
    \ces_4_1_io_outs_right[27] ,
    \ces_4_1_io_outs_right[26] ,
    \ces_4_1_io_outs_right[25] ,
    \ces_4_1_io_outs_right[24] ,
    \ces_4_1_io_outs_right[23] ,
    \ces_4_1_io_outs_right[22] ,
    \ces_4_1_io_outs_right[21] ,
    \ces_4_1_io_outs_right[20] ,
    \ces_4_1_io_outs_right[19] ,
    \ces_4_1_io_outs_right[18] ,
    \ces_4_1_io_outs_right[17] ,
    \ces_4_1_io_outs_right[16] ,
    \ces_4_1_io_outs_right[15] ,
    \ces_4_1_io_outs_right[14] ,
    \ces_4_1_io_outs_right[13] ,
    \ces_4_1_io_outs_right[12] ,
    \ces_4_1_io_outs_right[11] ,
    \ces_4_1_io_outs_right[10] ,
    \ces_4_1_io_outs_right[9] ,
    \ces_4_1_io_outs_right[8] ,
    \ces_4_1_io_outs_right[7] ,
    \ces_4_1_io_outs_right[6] ,
    \ces_4_1_io_outs_right[5] ,
    \ces_4_1_io_outs_right[4] ,
    \ces_4_1_io_outs_right[3] ,
    \ces_4_1_io_outs_right[2] ,
    \ces_4_1_io_outs_right[1] ,
    \ces_4_1_io_outs_right[0] }),
    .io_outs_up({\ces_4_1_io_outs_up[63] ,
    \ces_4_1_io_outs_up[62] ,
    \ces_4_1_io_outs_up[61] ,
    \ces_4_1_io_outs_up[60] ,
    \ces_4_1_io_outs_up[59] ,
    \ces_4_1_io_outs_up[58] ,
    \ces_4_1_io_outs_up[57] ,
    \ces_4_1_io_outs_up[56] ,
    \ces_4_1_io_outs_up[55] ,
    \ces_4_1_io_outs_up[54] ,
    \ces_4_1_io_outs_up[53] ,
    \ces_4_1_io_outs_up[52] ,
    \ces_4_1_io_outs_up[51] ,
    \ces_4_1_io_outs_up[50] ,
    \ces_4_1_io_outs_up[49] ,
    \ces_4_1_io_outs_up[48] ,
    \ces_4_1_io_outs_up[47] ,
    \ces_4_1_io_outs_up[46] ,
    \ces_4_1_io_outs_up[45] ,
    \ces_4_1_io_outs_up[44] ,
    \ces_4_1_io_outs_up[43] ,
    \ces_4_1_io_outs_up[42] ,
    \ces_4_1_io_outs_up[41] ,
    \ces_4_1_io_outs_up[40] ,
    \ces_4_1_io_outs_up[39] ,
    \ces_4_1_io_outs_up[38] ,
    \ces_4_1_io_outs_up[37] ,
    \ces_4_1_io_outs_up[36] ,
    \ces_4_1_io_outs_up[35] ,
    \ces_4_1_io_outs_up[34] ,
    \ces_4_1_io_outs_up[33] ,
    \ces_4_1_io_outs_up[32] ,
    \ces_4_1_io_outs_up[31] ,
    \ces_4_1_io_outs_up[30] ,
    \ces_4_1_io_outs_up[29] ,
    \ces_4_1_io_outs_up[28] ,
    \ces_4_1_io_outs_up[27] ,
    \ces_4_1_io_outs_up[26] ,
    \ces_4_1_io_outs_up[25] ,
    \ces_4_1_io_outs_up[24] ,
    \ces_4_1_io_outs_up[23] ,
    \ces_4_1_io_outs_up[22] ,
    \ces_4_1_io_outs_up[21] ,
    \ces_4_1_io_outs_up[20] ,
    \ces_4_1_io_outs_up[19] ,
    \ces_4_1_io_outs_up[18] ,
    \ces_4_1_io_outs_up[17] ,
    \ces_4_1_io_outs_up[16] ,
    \ces_4_1_io_outs_up[15] ,
    \ces_4_1_io_outs_up[14] ,
    \ces_4_1_io_outs_up[13] ,
    \ces_4_1_io_outs_up[12] ,
    \ces_4_1_io_outs_up[11] ,
    \ces_4_1_io_outs_up[10] ,
    \ces_4_1_io_outs_up[9] ,
    \ces_4_1_io_outs_up[8] ,
    \ces_4_1_io_outs_up[7] ,
    \ces_4_1_io_outs_up[6] ,
    \ces_4_1_io_outs_up[5] ,
    \ces_4_1_io_outs_up[4] ,
    \ces_4_1_io_outs_up[3] ,
    \ces_4_1_io_outs_up[2] ,
    \ces_4_1_io_outs_up[1] ,
    \ces_4_1_io_outs_up[0] }));
 Element ces_4_2 (.clock(clknet_3_4_0_clock),
    .io_lsbIns_1(ces_4_1_io_lsbOuts_1),
    .io_lsbIns_2(ces_4_1_io_lsbOuts_2),
    .io_lsbIns_3(ces_4_1_io_lsbOuts_3),
    .io_lsbIns_4(ces_4_1_io_lsbOuts_4),
    .io_lsbIns_5(ces_4_1_io_lsbOuts_5),
    .io_lsbIns_6(ces_4_1_io_lsbOuts_6),
    .io_lsbIns_7(ces_4_1_io_lsbOuts_7),
    .io_lsbOuts_0(ces_4_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_2_io_lsbOuts_7),
    .io_ins_down({\ces_4_2_io_ins_down[63] ,
    \ces_4_2_io_ins_down[62] ,
    \ces_4_2_io_ins_down[61] ,
    \ces_4_2_io_ins_down[60] ,
    \ces_4_2_io_ins_down[59] ,
    \ces_4_2_io_ins_down[58] ,
    \ces_4_2_io_ins_down[57] ,
    \ces_4_2_io_ins_down[56] ,
    \ces_4_2_io_ins_down[55] ,
    \ces_4_2_io_ins_down[54] ,
    \ces_4_2_io_ins_down[53] ,
    \ces_4_2_io_ins_down[52] ,
    \ces_4_2_io_ins_down[51] ,
    \ces_4_2_io_ins_down[50] ,
    \ces_4_2_io_ins_down[49] ,
    \ces_4_2_io_ins_down[48] ,
    \ces_4_2_io_ins_down[47] ,
    \ces_4_2_io_ins_down[46] ,
    \ces_4_2_io_ins_down[45] ,
    \ces_4_2_io_ins_down[44] ,
    \ces_4_2_io_ins_down[43] ,
    \ces_4_2_io_ins_down[42] ,
    \ces_4_2_io_ins_down[41] ,
    \ces_4_2_io_ins_down[40] ,
    \ces_4_2_io_ins_down[39] ,
    \ces_4_2_io_ins_down[38] ,
    \ces_4_2_io_ins_down[37] ,
    \ces_4_2_io_ins_down[36] ,
    \ces_4_2_io_ins_down[35] ,
    \ces_4_2_io_ins_down[34] ,
    \ces_4_2_io_ins_down[33] ,
    \ces_4_2_io_ins_down[32] ,
    \ces_4_2_io_ins_down[31] ,
    \ces_4_2_io_ins_down[30] ,
    \ces_4_2_io_ins_down[29] ,
    \ces_4_2_io_ins_down[28] ,
    \ces_4_2_io_ins_down[27] ,
    \ces_4_2_io_ins_down[26] ,
    \ces_4_2_io_ins_down[25] ,
    \ces_4_2_io_ins_down[24] ,
    \ces_4_2_io_ins_down[23] ,
    \ces_4_2_io_ins_down[22] ,
    \ces_4_2_io_ins_down[21] ,
    \ces_4_2_io_ins_down[20] ,
    \ces_4_2_io_ins_down[19] ,
    \ces_4_2_io_ins_down[18] ,
    \ces_4_2_io_ins_down[17] ,
    \ces_4_2_io_ins_down[16] ,
    \ces_4_2_io_ins_down[15] ,
    \ces_4_2_io_ins_down[14] ,
    \ces_4_2_io_ins_down[13] ,
    \ces_4_2_io_ins_down[12] ,
    \ces_4_2_io_ins_down[11] ,
    \ces_4_2_io_ins_down[10] ,
    \ces_4_2_io_ins_down[9] ,
    \ces_4_2_io_ins_down[8] ,
    \ces_4_2_io_ins_down[7] ,
    \ces_4_2_io_ins_down[6] ,
    \ces_4_2_io_ins_down[5] ,
    \ces_4_2_io_ins_down[4] ,
    \ces_4_2_io_ins_down[3] ,
    \ces_4_2_io_ins_down[2] ,
    \ces_4_2_io_ins_down[1] ,
    \ces_4_2_io_ins_down[0] }),
    .io_ins_left({\ces_4_2_io_ins_left[63] ,
    \ces_4_2_io_ins_left[62] ,
    \ces_4_2_io_ins_left[61] ,
    \ces_4_2_io_ins_left[60] ,
    \ces_4_2_io_ins_left[59] ,
    \ces_4_2_io_ins_left[58] ,
    \ces_4_2_io_ins_left[57] ,
    \ces_4_2_io_ins_left[56] ,
    \ces_4_2_io_ins_left[55] ,
    \ces_4_2_io_ins_left[54] ,
    \ces_4_2_io_ins_left[53] ,
    \ces_4_2_io_ins_left[52] ,
    \ces_4_2_io_ins_left[51] ,
    \ces_4_2_io_ins_left[50] ,
    \ces_4_2_io_ins_left[49] ,
    \ces_4_2_io_ins_left[48] ,
    \ces_4_2_io_ins_left[47] ,
    \ces_4_2_io_ins_left[46] ,
    \ces_4_2_io_ins_left[45] ,
    \ces_4_2_io_ins_left[44] ,
    \ces_4_2_io_ins_left[43] ,
    \ces_4_2_io_ins_left[42] ,
    \ces_4_2_io_ins_left[41] ,
    \ces_4_2_io_ins_left[40] ,
    \ces_4_2_io_ins_left[39] ,
    \ces_4_2_io_ins_left[38] ,
    \ces_4_2_io_ins_left[37] ,
    \ces_4_2_io_ins_left[36] ,
    \ces_4_2_io_ins_left[35] ,
    \ces_4_2_io_ins_left[34] ,
    \ces_4_2_io_ins_left[33] ,
    \ces_4_2_io_ins_left[32] ,
    \ces_4_2_io_ins_left[31] ,
    \ces_4_2_io_ins_left[30] ,
    \ces_4_2_io_ins_left[29] ,
    \ces_4_2_io_ins_left[28] ,
    \ces_4_2_io_ins_left[27] ,
    \ces_4_2_io_ins_left[26] ,
    \ces_4_2_io_ins_left[25] ,
    \ces_4_2_io_ins_left[24] ,
    \ces_4_2_io_ins_left[23] ,
    \ces_4_2_io_ins_left[22] ,
    \ces_4_2_io_ins_left[21] ,
    \ces_4_2_io_ins_left[20] ,
    \ces_4_2_io_ins_left[19] ,
    \ces_4_2_io_ins_left[18] ,
    \ces_4_2_io_ins_left[17] ,
    \ces_4_2_io_ins_left[16] ,
    \ces_4_2_io_ins_left[15] ,
    \ces_4_2_io_ins_left[14] ,
    \ces_4_2_io_ins_left[13] ,
    \ces_4_2_io_ins_left[12] ,
    \ces_4_2_io_ins_left[11] ,
    \ces_4_2_io_ins_left[10] ,
    \ces_4_2_io_ins_left[9] ,
    \ces_4_2_io_ins_left[8] ,
    \ces_4_2_io_ins_left[7] ,
    \ces_4_2_io_ins_left[6] ,
    \ces_4_2_io_ins_left[5] ,
    \ces_4_2_io_ins_left[4] ,
    \ces_4_2_io_ins_left[3] ,
    \ces_4_2_io_ins_left[2] ,
    \ces_4_2_io_ins_left[1] ,
    \ces_4_2_io_ins_left[0] }),
    .io_ins_right({\ces_4_1_io_outs_right[63] ,
    \ces_4_1_io_outs_right[62] ,
    \ces_4_1_io_outs_right[61] ,
    \ces_4_1_io_outs_right[60] ,
    \ces_4_1_io_outs_right[59] ,
    \ces_4_1_io_outs_right[58] ,
    \ces_4_1_io_outs_right[57] ,
    \ces_4_1_io_outs_right[56] ,
    \ces_4_1_io_outs_right[55] ,
    \ces_4_1_io_outs_right[54] ,
    \ces_4_1_io_outs_right[53] ,
    \ces_4_1_io_outs_right[52] ,
    \ces_4_1_io_outs_right[51] ,
    \ces_4_1_io_outs_right[50] ,
    \ces_4_1_io_outs_right[49] ,
    \ces_4_1_io_outs_right[48] ,
    \ces_4_1_io_outs_right[47] ,
    \ces_4_1_io_outs_right[46] ,
    \ces_4_1_io_outs_right[45] ,
    \ces_4_1_io_outs_right[44] ,
    \ces_4_1_io_outs_right[43] ,
    \ces_4_1_io_outs_right[42] ,
    \ces_4_1_io_outs_right[41] ,
    \ces_4_1_io_outs_right[40] ,
    \ces_4_1_io_outs_right[39] ,
    \ces_4_1_io_outs_right[38] ,
    \ces_4_1_io_outs_right[37] ,
    \ces_4_1_io_outs_right[36] ,
    \ces_4_1_io_outs_right[35] ,
    \ces_4_1_io_outs_right[34] ,
    \ces_4_1_io_outs_right[33] ,
    \ces_4_1_io_outs_right[32] ,
    \ces_4_1_io_outs_right[31] ,
    \ces_4_1_io_outs_right[30] ,
    \ces_4_1_io_outs_right[29] ,
    \ces_4_1_io_outs_right[28] ,
    \ces_4_1_io_outs_right[27] ,
    \ces_4_1_io_outs_right[26] ,
    \ces_4_1_io_outs_right[25] ,
    \ces_4_1_io_outs_right[24] ,
    \ces_4_1_io_outs_right[23] ,
    \ces_4_1_io_outs_right[22] ,
    \ces_4_1_io_outs_right[21] ,
    \ces_4_1_io_outs_right[20] ,
    \ces_4_1_io_outs_right[19] ,
    \ces_4_1_io_outs_right[18] ,
    \ces_4_1_io_outs_right[17] ,
    \ces_4_1_io_outs_right[16] ,
    \ces_4_1_io_outs_right[15] ,
    \ces_4_1_io_outs_right[14] ,
    \ces_4_1_io_outs_right[13] ,
    \ces_4_1_io_outs_right[12] ,
    \ces_4_1_io_outs_right[11] ,
    \ces_4_1_io_outs_right[10] ,
    \ces_4_1_io_outs_right[9] ,
    \ces_4_1_io_outs_right[8] ,
    \ces_4_1_io_outs_right[7] ,
    \ces_4_1_io_outs_right[6] ,
    \ces_4_1_io_outs_right[5] ,
    \ces_4_1_io_outs_right[4] ,
    \ces_4_1_io_outs_right[3] ,
    \ces_4_1_io_outs_right[2] ,
    \ces_4_1_io_outs_right[1] ,
    \ces_4_1_io_outs_right[0] }),
    .io_ins_up({\ces_3_2_io_outs_up[63] ,
    \ces_3_2_io_outs_up[62] ,
    \ces_3_2_io_outs_up[61] ,
    \ces_3_2_io_outs_up[60] ,
    \ces_3_2_io_outs_up[59] ,
    \ces_3_2_io_outs_up[58] ,
    \ces_3_2_io_outs_up[57] ,
    \ces_3_2_io_outs_up[56] ,
    \ces_3_2_io_outs_up[55] ,
    \ces_3_2_io_outs_up[54] ,
    \ces_3_2_io_outs_up[53] ,
    \ces_3_2_io_outs_up[52] ,
    \ces_3_2_io_outs_up[51] ,
    \ces_3_2_io_outs_up[50] ,
    \ces_3_2_io_outs_up[49] ,
    \ces_3_2_io_outs_up[48] ,
    \ces_3_2_io_outs_up[47] ,
    \ces_3_2_io_outs_up[46] ,
    \ces_3_2_io_outs_up[45] ,
    \ces_3_2_io_outs_up[44] ,
    \ces_3_2_io_outs_up[43] ,
    \ces_3_2_io_outs_up[42] ,
    \ces_3_2_io_outs_up[41] ,
    \ces_3_2_io_outs_up[40] ,
    \ces_3_2_io_outs_up[39] ,
    \ces_3_2_io_outs_up[38] ,
    \ces_3_2_io_outs_up[37] ,
    \ces_3_2_io_outs_up[36] ,
    \ces_3_2_io_outs_up[35] ,
    \ces_3_2_io_outs_up[34] ,
    \ces_3_2_io_outs_up[33] ,
    \ces_3_2_io_outs_up[32] ,
    \ces_3_2_io_outs_up[31] ,
    \ces_3_2_io_outs_up[30] ,
    \ces_3_2_io_outs_up[29] ,
    \ces_3_2_io_outs_up[28] ,
    \ces_3_2_io_outs_up[27] ,
    \ces_3_2_io_outs_up[26] ,
    \ces_3_2_io_outs_up[25] ,
    \ces_3_2_io_outs_up[24] ,
    \ces_3_2_io_outs_up[23] ,
    \ces_3_2_io_outs_up[22] ,
    \ces_3_2_io_outs_up[21] ,
    \ces_3_2_io_outs_up[20] ,
    \ces_3_2_io_outs_up[19] ,
    \ces_3_2_io_outs_up[18] ,
    \ces_3_2_io_outs_up[17] ,
    \ces_3_2_io_outs_up[16] ,
    \ces_3_2_io_outs_up[15] ,
    \ces_3_2_io_outs_up[14] ,
    \ces_3_2_io_outs_up[13] ,
    \ces_3_2_io_outs_up[12] ,
    \ces_3_2_io_outs_up[11] ,
    \ces_3_2_io_outs_up[10] ,
    \ces_3_2_io_outs_up[9] ,
    \ces_3_2_io_outs_up[8] ,
    \ces_3_2_io_outs_up[7] ,
    \ces_3_2_io_outs_up[6] ,
    \ces_3_2_io_outs_up[5] ,
    \ces_3_2_io_outs_up[4] ,
    \ces_3_2_io_outs_up[3] ,
    \ces_3_2_io_outs_up[2] ,
    \ces_3_2_io_outs_up[1] ,
    \ces_3_2_io_outs_up[0] }),
    .io_outs_down({\ces_3_2_io_ins_down[63] ,
    \ces_3_2_io_ins_down[62] ,
    \ces_3_2_io_ins_down[61] ,
    \ces_3_2_io_ins_down[60] ,
    \ces_3_2_io_ins_down[59] ,
    \ces_3_2_io_ins_down[58] ,
    \ces_3_2_io_ins_down[57] ,
    \ces_3_2_io_ins_down[56] ,
    \ces_3_2_io_ins_down[55] ,
    \ces_3_2_io_ins_down[54] ,
    \ces_3_2_io_ins_down[53] ,
    \ces_3_2_io_ins_down[52] ,
    \ces_3_2_io_ins_down[51] ,
    \ces_3_2_io_ins_down[50] ,
    \ces_3_2_io_ins_down[49] ,
    \ces_3_2_io_ins_down[48] ,
    \ces_3_2_io_ins_down[47] ,
    \ces_3_2_io_ins_down[46] ,
    \ces_3_2_io_ins_down[45] ,
    \ces_3_2_io_ins_down[44] ,
    \ces_3_2_io_ins_down[43] ,
    \ces_3_2_io_ins_down[42] ,
    \ces_3_2_io_ins_down[41] ,
    \ces_3_2_io_ins_down[40] ,
    \ces_3_2_io_ins_down[39] ,
    \ces_3_2_io_ins_down[38] ,
    \ces_3_2_io_ins_down[37] ,
    \ces_3_2_io_ins_down[36] ,
    \ces_3_2_io_ins_down[35] ,
    \ces_3_2_io_ins_down[34] ,
    \ces_3_2_io_ins_down[33] ,
    \ces_3_2_io_ins_down[32] ,
    \ces_3_2_io_ins_down[31] ,
    \ces_3_2_io_ins_down[30] ,
    \ces_3_2_io_ins_down[29] ,
    \ces_3_2_io_ins_down[28] ,
    \ces_3_2_io_ins_down[27] ,
    \ces_3_2_io_ins_down[26] ,
    \ces_3_2_io_ins_down[25] ,
    \ces_3_2_io_ins_down[24] ,
    \ces_3_2_io_ins_down[23] ,
    \ces_3_2_io_ins_down[22] ,
    \ces_3_2_io_ins_down[21] ,
    \ces_3_2_io_ins_down[20] ,
    \ces_3_2_io_ins_down[19] ,
    \ces_3_2_io_ins_down[18] ,
    \ces_3_2_io_ins_down[17] ,
    \ces_3_2_io_ins_down[16] ,
    \ces_3_2_io_ins_down[15] ,
    \ces_3_2_io_ins_down[14] ,
    \ces_3_2_io_ins_down[13] ,
    \ces_3_2_io_ins_down[12] ,
    \ces_3_2_io_ins_down[11] ,
    \ces_3_2_io_ins_down[10] ,
    \ces_3_2_io_ins_down[9] ,
    \ces_3_2_io_ins_down[8] ,
    \ces_3_2_io_ins_down[7] ,
    \ces_3_2_io_ins_down[6] ,
    \ces_3_2_io_ins_down[5] ,
    \ces_3_2_io_ins_down[4] ,
    \ces_3_2_io_ins_down[3] ,
    \ces_3_2_io_ins_down[2] ,
    \ces_3_2_io_ins_down[1] ,
    \ces_3_2_io_ins_down[0] }),
    .io_outs_left({\ces_4_1_io_ins_left[63] ,
    \ces_4_1_io_ins_left[62] ,
    \ces_4_1_io_ins_left[61] ,
    \ces_4_1_io_ins_left[60] ,
    \ces_4_1_io_ins_left[59] ,
    \ces_4_1_io_ins_left[58] ,
    \ces_4_1_io_ins_left[57] ,
    \ces_4_1_io_ins_left[56] ,
    \ces_4_1_io_ins_left[55] ,
    \ces_4_1_io_ins_left[54] ,
    \ces_4_1_io_ins_left[53] ,
    \ces_4_1_io_ins_left[52] ,
    \ces_4_1_io_ins_left[51] ,
    \ces_4_1_io_ins_left[50] ,
    \ces_4_1_io_ins_left[49] ,
    \ces_4_1_io_ins_left[48] ,
    \ces_4_1_io_ins_left[47] ,
    \ces_4_1_io_ins_left[46] ,
    \ces_4_1_io_ins_left[45] ,
    \ces_4_1_io_ins_left[44] ,
    \ces_4_1_io_ins_left[43] ,
    \ces_4_1_io_ins_left[42] ,
    \ces_4_1_io_ins_left[41] ,
    \ces_4_1_io_ins_left[40] ,
    \ces_4_1_io_ins_left[39] ,
    \ces_4_1_io_ins_left[38] ,
    \ces_4_1_io_ins_left[37] ,
    \ces_4_1_io_ins_left[36] ,
    \ces_4_1_io_ins_left[35] ,
    \ces_4_1_io_ins_left[34] ,
    \ces_4_1_io_ins_left[33] ,
    \ces_4_1_io_ins_left[32] ,
    \ces_4_1_io_ins_left[31] ,
    \ces_4_1_io_ins_left[30] ,
    \ces_4_1_io_ins_left[29] ,
    \ces_4_1_io_ins_left[28] ,
    \ces_4_1_io_ins_left[27] ,
    \ces_4_1_io_ins_left[26] ,
    \ces_4_1_io_ins_left[25] ,
    \ces_4_1_io_ins_left[24] ,
    \ces_4_1_io_ins_left[23] ,
    \ces_4_1_io_ins_left[22] ,
    \ces_4_1_io_ins_left[21] ,
    \ces_4_1_io_ins_left[20] ,
    \ces_4_1_io_ins_left[19] ,
    \ces_4_1_io_ins_left[18] ,
    \ces_4_1_io_ins_left[17] ,
    \ces_4_1_io_ins_left[16] ,
    \ces_4_1_io_ins_left[15] ,
    \ces_4_1_io_ins_left[14] ,
    \ces_4_1_io_ins_left[13] ,
    \ces_4_1_io_ins_left[12] ,
    \ces_4_1_io_ins_left[11] ,
    \ces_4_1_io_ins_left[10] ,
    \ces_4_1_io_ins_left[9] ,
    \ces_4_1_io_ins_left[8] ,
    \ces_4_1_io_ins_left[7] ,
    \ces_4_1_io_ins_left[6] ,
    \ces_4_1_io_ins_left[5] ,
    \ces_4_1_io_ins_left[4] ,
    \ces_4_1_io_ins_left[3] ,
    \ces_4_1_io_ins_left[2] ,
    \ces_4_1_io_ins_left[1] ,
    \ces_4_1_io_ins_left[0] }),
    .io_outs_right({\ces_4_2_io_outs_right[63] ,
    \ces_4_2_io_outs_right[62] ,
    \ces_4_2_io_outs_right[61] ,
    \ces_4_2_io_outs_right[60] ,
    \ces_4_2_io_outs_right[59] ,
    \ces_4_2_io_outs_right[58] ,
    \ces_4_2_io_outs_right[57] ,
    \ces_4_2_io_outs_right[56] ,
    \ces_4_2_io_outs_right[55] ,
    \ces_4_2_io_outs_right[54] ,
    \ces_4_2_io_outs_right[53] ,
    \ces_4_2_io_outs_right[52] ,
    \ces_4_2_io_outs_right[51] ,
    \ces_4_2_io_outs_right[50] ,
    \ces_4_2_io_outs_right[49] ,
    \ces_4_2_io_outs_right[48] ,
    \ces_4_2_io_outs_right[47] ,
    \ces_4_2_io_outs_right[46] ,
    \ces_4_2_io_outs_right[45] ,
    \ces_4_2_io_outs_right[44] ,
    \ces_4_2_io_outs_right[43] ,
    \ces_4_2_io_outs_right[42] ,
    \ces_4_2_io_outs_right[41] ,
    \ces_4_2_io_outs_right[40] ,
    \ces_4_2_io_outs_right[39] ,
    \ces_4_2_io_outs_right[38] ,
    \ces_4_2_io_outs_right[37] ,
    \ces_4_2_io_outs_right[36] ,
    \ces_4_2_io_outs_right[35] ,
    \ces_4_2_io_outs_right[34] ,
    \ces_4_2_io_outs_right[33] ,
    \ces_4_2_io_outs_right[32] ,
    \ces_4_2_io_outs_right[31] ,
    \ces_4_2_io_outs_right[30] ,
    \ces_4_2_io_outs_right[29] ,
    \ces_4_2_io_outs_right[28] ,
    \ces_4_2_io_outs_right[27] ,
    \ces_4_2_io_outs_right[26] ,
    \ces_4_2_io_outs_right[25] ,
    \ces_4_2_io_outs_right[24] ,
    \ces_4_2_io_outs_right[23] ,
    \ces_4_2_io_outs_right[22] ,
    \ces_4_2_io_outs_right[21] ,
    \ces_4_2_io_outs_right[20] ,
    \ces_4_2_io_outs_right[19] ,
    \ces_4_2_io_outs_right[18] ,
    \ces_4_2_io_outs_right[17] ,
    \ces_4_2_io_outs_right[16] ,
    \ces_4_2_io_outs_right[15] ,
    \ces_4_2_io_outs_right[14] ,
    \ces_4_2_io_outs_right[13] ,
    \ces_4_2_io_outs_right[12] ,
    \ces_4_2_io_outs_right[11] ,
    \ces_4_2_io_outs_right[10] ,
    \ces_4_2_io_outs_right[9] ,
    \ces_4_2_io_outs_right[8] ,
    \ces_4_2_io_outs_right[7] ,
    \ces_4_2_io_outs_right[6] ,
    \ces_4_2_io_outs_right[5] ,
    \ces_4_2_io_outs_right[4] ,
    \ces_4_2_io_outs_right[3] ,
    \ces_4_2_io_outs_right[2] ,
    \ces_4_2_io_outs_right[1] ,
    \ces_4_2_io_outs_right[0] }),
    .io_outs_up({\ces_4_2_io_outs_up[63] ,
    \ces_4_2_io_outs_up[62] ,
    \ces_4_2_io_outs_up[61] ,
    \ces_4_2_io_outs_up[60] ,
    \ces_4_2_io_outs_up[59] ,
    \ces_4_2_io_outs_up[58] ,
    \ces_4_2_io_outs_up[57] ,
    \ces_4_2_io_outs_up[56] ,
    \ces_4_2_io_outs_up[55] ,
    \ces_4_2_io_outs_up[54] ,
    \ces_4_2_io_outs_up[53] ,
    \ces_4_2_io_outs_up[52] ,
    \ces_4_2_io_outs_up[51] ,
    \ces_4_2_io_outs_up[50] ,
    \ces_4_2_io_outs_up[49] ,
    \ces_4_2_io_outs_up[48] ,
    \ces_4_2_io_outs_up[47] ,
    \ces_4_2_io_outs_up[46] ,
    \ces_4_2_io_outs_up[45] ,
    \ces_4_2_io_outs_up[44] ,
    \ces_4_2_io_outs_up[43] ,
    \ces_4_2_io_outs_up[42] ,
    \ces_4_2_io_outs_up[41] ,
    \ces_4_2_io_outs_up[40] ,
    \ces_4_2_io_outs_up[39] ,
    \ces_4_2_io_outs_up[38] ,
    \ces_4_2_io_outs_up[37] ,
    \ces_4_2_io_outs_up[36] ,
    \ces_4_2_io_outs_up[35] ,
    \ces_4_2_io_outs_up[34] ,
    \ces_4_2_io_outs_up[33] ,
    \ces_4_2_io_outs_up[32] ,
    \ces_4_2_io_outs_up[31] ,
    \ces_4_2_io_outs_up[30] ,
    \ces_4_2_io_outs_up[29] ,
    \ces_4_2_io_outs_up[28] ,
    \ces_4_2_io_outs_up[27] ,
    \ces_4_2_io_outs_up[26] ,
    \ces_4_2_io_outs_up[25] ,
    \ces_4_2_io_outs_up[24] ,
    \ces_4_2_io_outs_up[23] ,
    \ces_4_2_io_outs_up[22] ,
    \ces_4_2_io_outs_up[21] ,
    \ces_4_2_io_outs_up[20] ,
    \ces_4_2_io_outs_up[19] ,
    \ces_4_2_io_outs_up[18] ,
    \ces_4_2_io_outs_up[17] ,
    \ces_4_2_io_outs_up[16] ,
    \ces_4_2_io_outs_up[15] ,
    \ces_4_2_io_outs_up[14] ,
    \ces_4_2_io_outs_up[13] ,
    \ces_4_2_io_outs_up[12] ,
    \ces_4_2_io_outs_up[11] ,
    \ces_4_2_io_outs_up[10] ,
    \ces_4_2_io_outs_up[9] ,
    \ces_4_2_io_outs_up[8] ,
    \ces_4_2_io_outs_up[7] ,
    \ces_4_2_io_outs_up[6] ,
    \ces_4_2_io_outs_up[5] ,
    \ces_4_2_io_outs_up[4] ,
    \ces_4_2_io_outs_up[3] ,
    \ces_4_2_io_outs_up[2] ,
    \ces_4_2_io_outs_up[1] ,
    \ces_4_2_io_outs_up[0] }));
 Element ces_4_3 (.clock(clknet_3_4_0_clock),
    .io_lsbIns_1(ces_4_2_io_lsbOuts_1),
    .io_lsbIns_2(ces_4_2_io_lsbOuts_2),
    .io_lsbIns_3(ces_4_2_io_lsbOuts_3),
    .io_lsbIns_4(ces_4_2_io_lsbOuts_4),
    .io_lsbIns_5(ces_4_2_io_lsbOuts_5),
    .io_lsbIns_6(ces_4_2_io_lsbOuts_6),
    .io_lsbIns_7(ces_4_2_io_lsbOuts_7),
    .io_lsbOuts_0(ces_4_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_3_io_lsbOuts_7),
    .io_ins_down({\ces_4_3_io_ins_down[63] ,
    \ces_4_3_io_ins_down[62] ,
    \ces_4_3_io_ins_down[61] ,
    \ces_4_3_io_ins_down[60] ,
    \ces_4_3_io_ins_down[59] ,
    \ces_4_3_io_ins_down[58] ,
    \ces_4_3_io_ins_down[57] ,
    \ces_4_3_io_ins_down[56] ,
    \ces_4_3_io_ins_down[55] ,
    \ces_4_3_io_ins_down[54] ,
    \ces_4_3_io_ins_down[53] ,
    \ces_4_3_io_ins_down[52] ,
    \ces_4_3_io_ins_down[51] ,
    \ces_4_3_io_ins_down[50] ,
    \ces_4_3_io_ins_down[49] ,
    \ces_4_3_io_ins_down[48] ,
    \ces_4_3_io_ins_down[47] ,
    \ces_4_3_io_ins_down[46] ,
    \ces_4_3_io_ins_down[45] ,
    \ces_4_3_io_ins_down[44] ,
    \ces_4_3_io_ins_down[43] ,
    \ces_4_3_io_ins_down[42] ,
    \ces_4_3_io_ins_down[41] ,
    \ces_4_3_io_ins_down[40] ,
    \ces_4_3_io_ins_down[39] ,
    \ces_4_3_io_ins_down[38] ,
    \ces_4_3_io_ins_down[37] ,
    \ces_4_3_io_ins_down[36] ,
    \ces_4_3_io_ins_down[35] ,
    \ces_4_3_io_ins_down[34] ,
    \ces_4_3_io_ins_down[33] ,
    \ces_4_3_io_ins_down[32] ,
    \ces_4_3_io_ins_down[31] ,
    \ces_4_3_io_ins_down[30] ,
    \ces_4_3_io_ins_down[29] ,
    \ces_4_3_io_ins_down[28] ,
    \ces_4_3_io_ins_down[27] ,
    \ces_4_3_io_ins_down[26] ,
    \ces_4_3_io_ins_down[25] ,
    \ces_4_3_io_ins_down[24] ,
    \ces_4_3_io_ins_down[23] ,
    \ces_4_3_io_ins_down[22] ,
    \ces_4_3_io_ins_down[21] ,
    \ces_4_3_io_ins_down[20] ,
    \ces_4_3_io_ins_down[19] ,
    \ces_4_3_io_ins_down[18] ,
    \ces_4_3_io_ins_down[17] ,
    \ces_4_3_io_ins_down[16] ,
    \ces_4_3_io_ins_down[15] ,
    \ces_4_3_io_ins_down[14] ,
    \ces_4_3_io_ins_down[13] ,
    \ces_4_3_io_ins_down[12] ,
    \ces_4_3_io_ins_down[11] ,
    \ces_4_3_io_ins_down[10] ,
    \ces_4_3_io_ins_down[9] ,
    \ces_4_3_io_ins_down[8] ,
    \ces_4_3_io_ins_down[7] ,
    \ces_4_3_io_ins_down[6] ,
    \ces_4_3_io_ins_down[5] ,
    \ces_4_3_io_ins_down[4] ,
    \ces_4_3_io_ins_down[3] ,
    \ces_4_3_io_ins_down[2] ,
    \ces_4_3_io_ins_down[1] ,
    \ces_4_3_io_ins_down[0] }),
    .io_ins_left({\ces_4_3_io_ins_left[63] ,
    \ces_4_3_io_ins_left[62] ,
    \ces_4_3_io_ins_left[61] ,
    \ces_4_3_io_ins_left[60] ,
    \ces_4_3_io_ins_left[59] ,
    \ces_4_3_io_ins_left[58] ,
    \ces_4_3_io_ins_left[57] ,
    \ces_4_3_io_ins_left[56] ,
    \ces_4_3_io_ins_left[55] ,
    \ces_4_3_io_ins_left[54] ,
    \ces_4_3_io_ins_left[53] ,
    \ces_4_3_io_ins_left[52] ,
    \ces_4_3_io_ins_left[51] ,
    \ces_4_3_io_ins_left[50] ,
    \ces_4_3_io_ins_left[49] ,
    \ces_4_3_io_ins_left[48] ,
    \ces_4_3_io_ins_left[47] ,
    \ces_4_3_io_ins_left[46] ,
    \ces_4_3_io_ins_left[45] ,
    \ces_4_3_io_ins_left[44] ,
    \ces_4_3_io_ins_left[43] ,
    \ces_4_3_io_ins_left[42] ,
    \ces_4_3_io_ins_left[41] ,
    \ces_4_3_io_ins_left[40] ,
    \ces_4_3_io_ins_left[39] ,
    \ces_4_3_io_ins_left[38] ,
    \ces_4_3_io_ins_left[37] ,
    \ces_4_3_io_ins_left[36] ,
    \ces_4_3_io_ins_left[35] ,
    \ces_4_3_io_ins_left[34] ,
    \ces_4_3_io_ins_left[33] ,
    \ces_4_3_io_ins_left[32] ,
    \ces_4_3_io_ins_left[31] ,
    \ces_4_3_io_ins_left[30] ,
    \ces_4_3_io_ins_left[29] ,
    \ces_4_3_io_ins_left[28] ,
    \ces_4_3_io_ins_left[27] ,
    \ces_4_3_io_ins_left[26] ,
    \ces_4_3_io_ins_left[25] ,
    \ces_4_3_io_ins_left[24] ,
    \ces_4_3_io_ins_left[23] ,
    \ces_4_3_io_ins_left[22] ,
    \ces_4_3_io_ins_left[21] ,
    \ces_4_3_io_ins_left[20] ,
    \ces_4_3_io_ins_left[19] ,
    \ces_4_3_io_ins_left[18] ,
    \ces_4_3_io_ins_left[17] ,
    \ces_4_3_io_ins_left[16] ,
    \ces_4_3_io_ins_left[15] ,
    \ces_4_3_io_ins_left[14] ,
    \ces_4_3_io_ins_left[13] ,
    \ces_4_3_io_ins_left[12] ,
    \ces_4_3_io_ins_left[11] ,
    \ces_4_3_io_ins_left[10] ,
    \ces_4_3_io_ins_left[9] ,
    \ces_4_3_io_ins_left[8] ,
    \ces_4_3_io_ins_left[7] ,
    \ces_4_3_io_ins_left[6] ,
    \ces_4_3_io_ins_left[5] ,
    \ces_4_3_io_ins_left[4] ,
    \ces_4_3_io_ins_left[3] ,
    \ces_4_3_io_ins_left[2] ,
    \ces_4_3_io_ins_left[1] ,
    \ces_4_3_io_ins_left[0] }),
    .io_ins_right({\ces_4_2_io_outs_right[63] ,
    \ces_4_2_io_outs_right[62] ,
    \ces_4_2_io_outs_right[61] ,
    \ces_4_2_io_outs_right[60] ,
    \ces_4_2_io_outs_right[59] ,
    \ces_4_2_io_outs_right[58] ,
    \ces_4_2_io_outs_right[57] ,
    \ces_4_2_io_outs_right[56] ,
    \ces_4_2_io_outs_right[55] ,
    \ces_4_2_io_outs_right[54] ,
    \ces_4_2_io_outs_right[53] ,
    \ces_4_2_io_outs_right[52] ,
    \ces_4_2_io_outs_right[51] ,
    \ces_4_2_io_outs_right[50] ,
    \ces_4_2_io_outs_right[49] ,
    \ces_4_2_io_outs_right[48] ,
    \ces_4_2_io_outs_right[47] ,
    \ces_4_2_io_outs_right[46] ,
    \ces_4_2_io_outs_right[45] ,
    \ces_4_2_io_outs_right[44] ,
    \ces_4_2_io_outs_right[43] ,
    \ces_4_2_io_outs_right[42] ,
    \ces_4_2_io_outs_right[41] ,
    \ces_4_2_io_outs_right[40] ,
    \ces_4_2_io_outs_right[39] ,
    \ces_4_2_io_outs_right[38] ,
    \ces_4_2_io_outs_right[37] ,
    \ces_4_2_io_outs_right[36] ,
    \ces_4_2_io_outs_right[35] ,
    \ces_4_2_io_outs_right[34] ,
    \ces_4_2_io_outs_right[33] ,
    \ces_4_2_io_outs_right[32] ,
    \ces_4_2_io_outs_right[31] ,
    \ces_4_2_io_outs_right[30] ,
    \ces_4_2_io_outs_right[29] ,
    \ces_4_2_io_outs_right[28] ,
    \ces_4_2_io_outs_right[27] ,
    \ces_4_2_io_outs_right[26] ,
    \ces_4_2_io_outs_right[25] ,
    \ces_4_2_io_outs_right[24] ,
    \ces_4_2_io_outs_right[23] ,
    \ces_4_2_io_outs_right[22] ,
    \ces_4_2_io_outs_right[21] ,
    \ces_4_2_io_outs_right[20] ,
    \ces_4_2_io_outs_right[19] ,
    \ces_4_2_io_outs_right[18] ,
    \ces_4_2_io_outs_right[17] ,
    \ces_4_2_io_outs_right[16] ,
    \ces_4_2_io_outs_right[15] ,
    \ces_4_2_io_outs_right[14] ,
    \ces_4_2_io_outs_right[13] ,
    \ces_4_2_io_outs_right[12] ,
    \ces_4_2_io_outs_right[11] ,
    \ces_4_2_io_outs_right[10] ,
    \ces_4_2_io_outs_right[9] ,
    \ces_4_2_io_outs_right[8] ,
    \ces_4_2_io_outs_right[7] ,
    \ces_4_2_io_outs_right[6] ,
    \ces_4_2_io_outs_right[5] ,
    \ces_4_2_io_outs_right[4] ,
    \ces_4_2_io_outs_right[3] ,
    \ces_4_2_io_outs_right[2] ,
    \ces_4_2_io_outs_right[1] ,
    \ces_4_2_io_outs_right[0] }),
    .io_ins_up({\ces_3_3_io_outs_up[63] ,
    \ces_3_3_io_outs_up[62] ,
    \ces_3_3_io_outs_up[61] ,
    \ces_3_3_io_outs_up[60] ,
    \ces_3_3_io_outs_up[59] ,
    \ces_3_3_io_outs_up[58] ,
    \ces_3_3_io_outs_up[57] ,
    \ces_3_3_io_outs_up[56] ,
    \ces_3_3_io_outs_up[55] ,
    \ces_3_3_io_outs_up[54] ,
    \ces_3_3_io_outs_up[53] ,
    \ces_3_3_io_outs_up[52] ,
    \ces_3_3_io_outs_up[51] ,
    \ces_3_3_io_outs_up[50] ,
    \ces_3_3_io_outs_up[49] ,
    \ces_3_3_io_outs_up[48] ,
    \ces_3_3_io_outs_up[47] ,
    \ces_3_3_io_outs_up[46] ,
    \ces_3_3_io_outs_up[45] ,
    \ces_3_3_io_outs_up[44] ,
    \ces_3_3_io_outs_up[43] ,
    \ces_3_3_io_outs_up[42] ,
    \ces_3_3_io_outs_up[41] ,
    \ces_3_3_io_outs_up[40] ,
    \ces_3_3_io_outs_up[39] ,
    \ces_3_3_io_outs_up[38] ,
    \ces_3_3_io_outs_up[37] ,
    \ces_3_3_io_outs_up[36] ,
    \ces_3_3_io_outs_up[35] ,
    \ces_3_3_io_outs_up[34] ,
    \ces_3_3_io_outs_up[33] ,
    \ces_3_3_io_outs_up[32] ,
    \ces_3_3_io_outs_up[31] ,
    \ces_3_3_io_outs_up[30] ,
    \ces_3_3_io_outs_up[29] ,
    \ces_3_3_io_outs_up[28] ,
    \ces_3_3_io_outs_up[27] ,
    \ces_3_3_io_outs_up[26] ,
    \ces_3_3_io_outs_up[25] ,
    \ces_3_3_io_outs_up[24] ,
    \ces_3_3_io_outs_up[23] ,
    \ces_3_3_io_outs_up[22] ,
    \ces_3_3_io_outs_up[21] ,
    \ces_3_3_io_outs_up[20] ,
    \ces_3_3_io_outs_up[19] ,
    \ces_3_3_io_outs_up[18] ,
    \ces_3_3_io_outs_up[17] ,
    \ces_3_3_io_outs_up[16] ,
    \ces_3_3_io_outs_up[15] ,
    \ces_3_3_io_outs_up[14] ,
    \ces_3_3_io_outs_up[13] ,
    \ces_3_3_io_outs_up[12] ,
    \ces_3_3_io_outs_up[11] ,
    \ces_3_3_io_outs_up[10] ,
    \ces_3_3_io_outs_up[9] ,
    \ces_3_3_io_outs_up[8] ,
    \ces_3_3_io_outs_up[7] ,
    \ces_3_3_io_outs_up[6] ,
    \ces_3_3_io_outs_up[5] ,
    \ces_3_3_io_outs_up[4] ,
    \ces_3_3_io_outs_up[3] ,
    \ces_3_3_io_outs_up[2] ,
    \ces_3_3_io_outs_up[1] ,
    \ces_3_3_io_outs_up[0] }),
    .io_outs_down({\ces_3_3_io_ins_down[63] ,
    \ces_3_3_io_ins_down[62] ,
    \ces_3_3_io_ins_down[61] ,
    \ces_3_3_io_ins_down[60] ,
    \ces_3_3_io_ins_down[59] ,
    \ces_3_3_io_ins_down[58] ,
    \ces_3_3_io_ins_down[57] ,
    \ces_3_3_io_ins_down[56] ,
    \ces_3_3_io_ins_down[55] ,
    \ces_3_3_io_ins_down[54] ,
    \ces_3_3_io_ins_down[53] ,
    \ces_3_3_io_ins_down[52] ,
    \ces_3_3_io_ins_down[51] ,
    \ces_3_3_io_ins_down[50] ,
    \ces_3_3_io_ins_down[49] ,
    \ces_3_3_io_ins_down[48] ,
    \ces_3_3_io_ins_down[47] ,
    \ces_3_3_io_ins_down[46] ,
    \ces_3_3_io_ins_down[45] ,
    \ces_3_3_io_ins_down[44] ,
    \ces_3_3_io_ins_down[43] ,
    \ces_3_3_io_ins_down[42] ,
    \ces_3_3_io_ins_down[41] ,
    \ces_3_3_io_ins_down[40] ,
    \ces_3_3_io_ins_down[39] ,
    \ces_3_3_io_ins_down[38] ,
    \ces_3_3_io_ins_down[37] ,
    \ces_3_3_io_ins_down[36] ,
    \ces_3_3_io_ins_down[35] ,
    \ces_3_3_io_ins_down[34] ,
    \ces_3_3_io_ins_down[33] ,
    \ces_3_3_io_ins_down[32] ,
    \ces_3_3_io_ins_down[31] ,
    \ces_3_3_io_ins_down[30] ,
    \ces_3_3_io_ins_down[29] ,
    \ces_3_3_io_ins_down[28] ,
    \ces_3_3_io_ins_down[27] ,
    \ces_3_3_io_ins_down[26] ,
    \ces_3_3_io_ins_down[25] ,
    \ces_3_3_io_ins_down[24] ,
    \ces_3_3_io_ins_down[23] ,
    \ces_3_3_io_ins_down[22] ,
    \ces_3_3_io_ins_down[21] ,
    \ces_3_3_io_ins_down[20] ,
    \ces_3_3_io_ins_down[19] ,
    \ces_3_3_io_ins_down[18] ,
    \ces_3_3_io_ins_down[17] ,
    \ces_3_3_io_ins_down[16] ,
    \ces_3_3_io_ins_down[15] ,
    \ces_3_3_io_ins_down[14] ,
    \ces_3_3_io_ins_down[13] ,
    \ces_3_3_io_ins_down[12] ,
    \ces_3_3_io_ins_down[11] ,
    \ces_3_3_io_ins_down[10] ,
    \ces_3_3_io_ins_down[9] ,
    \ces_3_3_io_ins_down[8] ,
    \ces_3_3_io_ins_down[7] ,
    \ces_3_3_io_ins_down[6] ,
    \ces_3_3_io_ins_down[5] ,
    \ces_3_3_io_ins_down[4] ,
    \ces_3_3_io_ins_down[3] ,
    \ces_3_3_io_ins_down[2] ,
    \ces_3_3_io_ins_down[1] ,
    \ces_3_3_io_ins_down[0] }),
    .io_outs_left({\ces_4_2_io_ins_left[63] ,
    \ces_4_2_io_ins_left[62] ,
    \ces_4_2_io_ins_left[61] ,
    \ces_4_2_io_ins_left[60] ,
    \ces_4_2_io_ins_left[59] ,
    \ces_4_2_io_ins_left[58] ,
    \ces_4_2_io_ins_left[57] ,
    \ces_4_2_io_ins_left[56] ,
    \ces_4_2_io_ins_left[55] ,
    \ces_4_2_io_ins_left[54] ,
    \ces_4_2_io_ins_left[53] ,
    \ces_4_2_io_ins_left[52] ,
    \ces_4_2_io_ins_left[51] ,
    \ces_4_2_io_ins_left[50] ,
    \ces_4_2_io_ins_left[49] ,
    \ces_4_2_io_ins_left[48] ,
    \ces_4_2_io_ins_left[47] ,
    \ces_4_2_io_ins_left[46] ,
    \ces_4_2_io_ins_left[45] ,
    \ces_4_2_io_ins_left[44] ,
    \ces_4_2_io_ins_left[43] ,
    \ces_4_2_io_ins_left[42] ,
    \ces_4_2_io_ins_left[41] ,
    \ces_4_2_io_ins_left[40] ,
    \ces_4_2_io_ins_left[39] ,
    \ces_4_2_io_ins_left[38] ,
    \ces_4_2_io_ins_left[37] ,
    \ces_4_2_io_ins_left[36] ,
    \ces_4_2_io_ins_left[35] ,
    \ces_4_2_io_ins_left[34] ,
    \ces_4_2_io_ins_left[33] ,
    \ces_4_2_io_ins_left[32] ,
    \ces_4_2_io_ins_left[31] ,
    \ces_4_2_io_ins_left[30] ,
    \ces_4_2_io_ins_left[29] ,
    \ces_4_2_io_ins_left[28] ,
    \ces_4_2_io_ins_left[27] ,
    \ces_4_2_io_ins_left[26] ,
    \ces_4_2_io_ins_left[25] ,
    \ces_4_2_io_ins_left[24] ,
    \ces_4_2_io_ins_left[23] ,
    \ces_4_2_io_ins_left[22] ,
    \ces_4_2_io_ins_left[21] ,
    \ces_4_2_io_ins_left[20] ,
    \ces_4_2_io_ins_left[19] ,
    \ces_4_2_io_ins_left[18] ,
    \ces_4_2_io_ins_left[17] ,
    \ces_4_2_io_ins_left[16] ,
    \ces_4_2_io_ins_left[15] ,
    \ces_4_2_io_ins_left[14] ,
    \ces_4_2_io_ins_left[13] ,
    \ces_4_2_io_ins_left[12] ,
    \ces_4_2_io_ins_left[11] ,
    \ces_4_2_io_ins_left[10] ,
    \ces_4_2_io_ins_left[9] ,
    \ces_4_2_io_ins_left[8] ,
    \ces_4_2_io_ins_left[7] ,
    \ces_4_2_io_ins_left[6] ,
    \ces_4_2_io_ins_left[5] ,
    \ces_4_2_io_ins_left[4] ,
    \ces_4_2_io_ins_left[3] ,
    \ces_4_2_io_ins_left[2] ,
    \ces_4_2_io_ins_left[1] ,
    \ces_4_2_io_ins_left[0] }),
    .io_outs_right({\ces_4_3_io_outs_right[63] ,
    \ces_4_3_io_outs_right[62] ,
    \ces_4_3_io_outs_right[61] ,
    \ces_4_3_io_outs_right[60] ,
    \ces_4_3_io_outs_right[59] ,
    \ces_4_3_io_outs_right[58] ,
    \ces_4_3_io_outs_right[57] ,
    \ces_4_3_io_outs_right[56] ,
    \ces_4_3_io_outs_right[55] ,
    \ces_4_3_io_outs_right[54] ,
    \ces_4_3_io_outs_right[53] ,
    \ces_4_3_io_outs_right[52] ,
    \ces_4_3_io_outs_right[51] ,
    \ces_4_3_io_outs_right[50] ,
    \ces_4_3_io_outs_right[49] ,
    \ces_4_3_io_outs_right[48] ,
    \ces_4_3_io_outs_right[47] ,
    \ces_4_3_io_outs_right[46] ,
    \ces_4_3_io_outs_right[45] ,
    \ces_4_3_io_outs_right[44] ,
    \ces_4_3_io_outs_right[43] ,
    \ces_4_3_io_outs_right[42] ,
    \ces_4_3_io_outs_right[41] ,
    \ces_4_3_io_outs_right[40] ,
    \ces_4_3_io_outs_right[39] ,
    \ces_4_3_io_outs_right[38] ,
    \ces_4_3_io_outs_right[37] ,
    \ces_4_3_io_outs_right[36] ,
    \ces_4_3_io_outs_right[35] ,
    \ces_4_3_io_outs_right[34] ,
    \ces_4_3_io_outs_right[33] ,
    \ces_4_3_io_outs_right[32] ,
    \ces_4_3_io_outs_right[31] ,
    \ces_4_3_io_outs_right[30] ,
    \ces_4_3_io_outs_right[29] ,
    \ces_4_3_io_outs_right[28] ,
    \ces_4_3_io_outs_right[27] ,
    \ces_4_3_io_outs_right[26] ,
    \ces_4_3_io_outs_right[25] ,
    \ces_4_3_io_outs_right[24] ,
    \ces_4_3_io_outs_right[23] ,
    \ces_4_3_io_outs_right[22] ,
    \ces_4_3_io_outs_right[21] ,
    \ces_4_3_io_outs_right[20] ,
    \ces_4_3_io_outs_right[19] ,
    \ces_4_3_io_outs_right[18] ,
    \ces_4_3_io_outs_right[17] ,
    \ces_4_3_io_outs_right[16] ,
    \ces_4_3_io_outs_right[15] ,
    \ces_4_3_io_outs_right[14] ,
    \ces_4_3_io_outs_right[13] ,
    \ces_4_3_io_outs_right[12] ,
    \ces_4_3_io_outs_right[11] ,
    \ces_4_3_io_outs_right[10] ,
    \ces_4_3_io_outs_right[9] ,
    \ces_4_3_io_outs_right[8] ,
    \ces_4_3_io_outs_right[7] ,
    \ces_4_3_io_outs_right[6] ,
    \ces_4_3_io_outs_right[5] ,
    \ces_4_3_io_outs_right[4] ,
    \ces_4_3_io_outs_right[3] ,
    \ces_4_3_io_outs_right[2] ,
    \ces_4_3_io_outs_right[1] ,
    \ces_4_3_io_outs_right[0] }),
    .io_outs_up({\ces_4_3_io_outs_up[63] ,
    \ces_4_3_io_outs_up[62] ,
    \ces_4_3_io_outs_up[61] ,
    \ces_4_3_io_outs_up[60] ,
    \ces_4_3_io_outs_up[59] ,
    \ces_4_3_io_outs_up[58] ,
    \ces_4_3_io_outs_up[57] ,
    \ces_4_3_io_outs_up[56] ,
    \ces_4_3_io_outs_up[55] ,
    \ces_4_3_io_outs_up[54] ,
    \ces_4_3_io_outs_up[53] ,
    \ces_4_3_io_outs_up[52] ,
    \ces_4_3_io_outs_up[51] ,
    \ces_4_3_io_outs_up[50] ,
    \ces_4_3_io_outs_up[49] ,
    \ces_4_3_io_outs_up[48] ,
    \ces_4_3_io_outs_up[47] ,
    \ces_4_3_io_outs_up[46] ,
    \ces_4_3_io_outs_up[45] ,
    \ces_4_3_io_outs_up[44] ,
    \ces_4_3_io_outs_up[43] ,
    \ces_4_3_io_outs_up[42] ,
    \ces_4_3_io_outs_up[41] ,
    \ces_4_3_io_outs_up[40] ,
    \ces_4_3_io_outs_up[39] ,
    \ces_4_3_io_outs_up[38] ,
    \ces_4_3_io_outs_up[37] ,
    \ces_4_3_io_outs_up[36] ,
    \ces_4_3_io_outs_up[35] ,
    \ces_4_3_io_outs_up[34] ,
    \ces_4_3_io_outs_up[33] ,
    \ces_4_3_io_outs_up[32] ,
    \ces_4_3_io_outs_up[31] ,
    \ces_4_3_io_outs_up[30] ,
    \ces_4_3_io_outs_up[29] ,
    \ces_4_3_io_outs_up[28] ,
    \ces_4_3_io_outs_up[27] ,
    \ces_4_3_io_outs_up[26] ,
    \ces_4_3_io_outs_up[25] ,
    \ces_4_3_io_outs_up[24] ,
    \ces_4_3_io_outs_up[23] ,
    \ces_4_3_io_outs_up[22] ,
    \ces_4_3_io_outs_up[21] ,
    \ces_4_3_io_outs_up[20] ,
    \ces_4_3_io_outs_up[19] ,
    \ces_4_3_io_outs_up[18] ,
    \ces_4_3_io_outs_up[17] ,
    \ces_4_3_io_outs_up[16] ,
    \ces_4_3_io_outs_up[15] ,
    \ces_4_3_io_outs_up[14] ,
    \ces_4_3_io_outs_up[13] ,
    \ces_4_3_io_outs_up[12] ,
    \ces_4_3_io_outs_up[11] ,
    \ces_4_3_io_outs_up[10] ,
    \ces_4_3_io_outs_up[9] ,
    \ces_4_3_io_outs_up[8] ,
    \ces_4_3_io_outs_up[7] ,
    \ces_4_3_io_outs_up[6] ,
    \ces_4_3_io_outs_up[5] ,
    \ces_4_3_io_outs_up[4] ,
    \ces_4_3_io_outs_up[3] ,
    \ces_4_3_io_outs_up[2] ,
    \ces_4_3_io_outs_up[1] ,
    \ces_4_3_io_outs_up[0] }));
 Element ces_4_4 (.clock(clknet_3_6_0_clock),
    .io_lsbIns_1(ces_4_3_io_lsbOuts_1),
    .io_lsbIns_2(ces_4_3_io_lsbOuts_2),
    .io_lsbIns_3(ces_4_3_io_lsbOuts_3),
    .io_lsbIns_4(ces_4_3_io_lsbOuts_4),
    .io_lsbIns_5(ces_4_3_io_lsbOuts_5),
    .io_lsbIns_6(ces_4_3_io_lsbOuts_6),
    .io_lsbIns_7(ces_4_3_io_lsbOuts_7),
    .io_lsbOuts_0(ces_4_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_4_io_lsbOuts_7),
    .io_ins_down({\ces_4_4_io_ins_down[63] ,
    \ces_4_4_io_ins_down[62] ,
    \ces_4_4_io_ins_down[61] ,
    \ces_4_4_io_ins_down[60] ,
    \ces_4_4_io_ins_down[59] ,
    \ces_4_4_io_ins_down[58] ,
    \ces_4_4_io_ins_down[57] ,
    \ces_4_4_io_ins_down[56] ,
    \ces_4_4_io_ins_down[55] ,
    \ces_4_4_io_ins_down[54] ,
    \ces_4_4_io_ins_down[53] ,
    \ces_4_4_io_ins_down[52] ,
    \ces_4_4_io_ins_down[51] ,
    \ces_4_4_io_ins_down[50] ,
    \ces_4_4_io_ins_down[49] ,
    \ces_4_4_io_ins_down[48] ,
    \ces_4_4_io_ins_down[47] ,
    \ces_4_4_io_ins_down[46] ,
    \ces_4_4_io_ins_down[45] ,
    \ces_4_4_io_ins_down[44] ,
    \ces_4_4_io_ins_down[43] ,
    \ces_4_4_io_ins_down[42] ,
    \ces_4_4_io_ins_down[41] ,
    \ces_4_4_io_ins_down[40] ,
    \ces_4_4_io_ins_down[39] ,
    \ces_4_4_io_ins_down[38] ,
    \ces_4_4_io_ins_down[37] ,
    \ces_4_4_io_ins_down[36] ,
    \ces_4_4_io_ins_down[35] ,
    \ces_4_4_io_ins_down[34] ,
    \ces_4_4_io_ins_down[33] ,
    \ces_4_4_io_ins_down[32] ,
    \ces_4_4_io_ins_down[31] ,
    \ces_4_4_io_ins_down[30] ,
    \ces_4_4_io_ins_down[29] ,
    \ces_4_4_io_ins_down[28] ,
    \ces_4_4_io_ins_down[27] ,
    \ces_4_4_io_ins_down[26] ,
    \ces_4_4_io_ins_down[25] ,
    \ces_4_4_io_ins_down[24] ,
    \ces_4_4_io_ins_down[23] ,
    \ces_4_4_io_ins_down[22] ,
    \ces_4_4_io_ins_down[21] ,
    \ces_4_4_io_ins_down[20] ,
    \ces_4_4_io_ins_down[19] ,
    \ces_4_4_io_ins_down[18] ,
    \ces_4_4_io_ins_down[17] ,
    \ces_4_4_io_ins_down[16] ,
    \ces_4_4_io_ins_down[15] ,
    \ces_4_4_io_ins_down[14] ,
    \ces_4_4_io_ins_down[13] ,
    \ces_4_4_io_ins_down[12] ,
    \ces_4_4_io_ins_down[11] ,
    \ces_4_4_io_ins_down[10] ,
    \ces_4_4_io_ins_down[9] ,
    \ces_4_4_io_ins_down[8] ,
    \ces_4_4_io_ins_down[7] ,
    \ces_4_4_io_ins_down[6] ,
    \ces_4_4_io_ins_down[5] ,
    \ces_4_4_io_ins_down[4] ,
    \ces_4_4_io_ins_down[3] ,
    \ces_4_4_io_ins_down[2] ,
    \ces_4_4_io_ins_down[1] ,
    \ces_4_4_io_ins_down[0] }),
    .io_ins_left({\ces_4_4_io_ins_left[63] ,
    \ces_4_4_io_ins_left[62] ,
    \ces_4_4_io_ins_left[61] ,
    \ces_4_4_io_ins_left[60] ,
    \ces_4_4_io_ins_left[59] ,
    \ces_4_4_io_ins_left[58] ,
    \ces_4_4_io_ins_left[57] ,
    \ces_4_4_io_ins_left[56] ,
    \ces_4_4_io_ins_left[55] ,
    \ces_4_4_io_ins_left[54] ,
    \ces_4_4_io_ins_left[53] ,
    \ces_4_4_io_ins_left[52] ,
    \ces_4_4_io_ins_left[51] ,
    \ces_4_4_io_ins_left[50] ,
    \ces_4_4_io_ins_left[49] ,
    \ces_4_4_io_ins_left[48] ,
    \ces_4_4_io_ins_left[47] ,
    \ces_4_4_io_ins_left[46] ,
    \ces_4_4_io_ins_left[45] ,
    \ces_4_4_io_ins_left[44] ,
    \ces_4_4_io_ins_left[43] ,
    \ces_4_4_io_ins_left[42] ,
    \ces_4_4_io_ins_left[41] ,
    \ces_4_4_io_ins_left[40] ,
    \ces_4_4_io_ins_left[39] ,
    \ces_4_4_io_ins_left[38] ,
    \ces_4_4_io_ins_left[37] ,
    \ces_4_4_io_ins_left[36] ,
    \ces_4_4_io_ins_left[35] ,
    \ces_4_4_io_ins_left[34] ,
    \ces_4_4_io_ins_left[33] ,
    \ces_4_4_io_ins_left[32] ,
    \ces_4_4_io_ins_left[31] ,
    \ces_4_4_io_ins_left[30] ,
    \ces_4_4_io_ins_left[29] ,
    \ces_4_4_io_ins_left[28] ,
    \ces_4_4_io_ins_left[27] ,
    \ces_4_4_io_ins_left[26] ,
    \ces_4_4_io_ins_left[25] ,
    \ces_4_4_io_ins_left[24] ,
    \ces_4_4_io_ins_left[23] ,
    \ces_4_4_io_ins_left[22] ,
    \ces_4_4_io_ins_left[21] ,
    \ces_4_4_io_ins_left[20] ,
    \ces_4_4_io_ins_left[19] ,
    \ces_4_4_io_ins_left[18] ,
    \ces_4_4_io_ins_left[17] ,
    \ces_4_4_io_ins_left[16] ,
    \ces_4_4_io_ins_left[15] ,
    \ces_4_4_io_ins_left[14] ,
    \ces_4_4_io_ins_left[13] ,
    \ces_4_4_io_ins_left[12] ,
    \ces_4_4_io_ins_left[11] ,
    \ces_4_4_io_ins_left[10] ,
    \ces_4_4_io_ins_left[9] ,
    \ces_4_4_io_ins_left[8] ,
    \ces_4_4_io_ins_left[7] ,
    \ces_4_4_io_ins_left[6] ,
    \ces_4_4_io_ins_left[5] ,
    \ces_4_4_io_ins_left[4] ,
    \ces_4_4_io_ins_left[3] ,
    \ces_4_4_io_ins_left[2] ,
    \ces_4_4_io_ins_left[1] ,
    \ces_4_4_io_ins_left[0] }),
    .io_ins_right({\ces_4_3_io_outs_right[63] ,
    \ces_4_3_io_outs_right[62] ,
    \ces_4_3_io_outs_right[61] ,
    \ces_4_3_io_outs_right[60] ,
    \ces_4_3_io_outs_right[59] ,
    \ces_4_3_io_outs_right[58] ,
    \ces_4_3_io_outs_right[57] ,
    \ces_4_3_io_outs_right[56] ,
    \ces_4_3_io_outs_right[55] ,
    \ces_4_3_io_outs_right[54] ,
    \ces_4_3_io_outs_right[53] ,
    \ces_4_3_io_outs_right[52] ,
    \ces_4_3_io_outs_right[51] ,
    \ces_4_3_io_outs_right[50] ,
    \ces_4_3_io_outs_right[49] ,
    \ces_4_3_io_outs_right[48] ,
    \ces_4_3_io_outs_right[47] ,
    \ces_4_3_io_outs_right[46] ,
    \ces_4_3_io_outs_right[45] ,
    \ces_4_3_io_outs_right[44] ,
    \ces_4_3_io_outs_right[43] ,
    \ces_4_3_io_outs_right[42] ,
    \ces_4_3_io_outs_right[41] ,
    \ces_4_3_io_outs_right[40] ,
    \ces_4_3_io_outs_right[39] ,
    \ces_4_3_io_outs_right[38] ,
    \ces_4_3_io_outs_right[37] ,
    \ces_4_3_io_outs_right[36] ,
    \ces_4_3_io_outs_right[35] ,
    \ces_4_3_io_outs_right[34] ,
    \ces_4_3_io_outs_right[33] ,
    \ces_4_3_io_outs_right[32] ,
    \ces_4_3_io_outs_right[31] ,
    \ces_4_3_io_outs_right[30] ,
    \ces_4_3_io_outs_right[29] ,
    \ces_4_3_io_outs_right[28] ,
    \ces_4_3_io_outs_right[27] ,
    \ces_4_3_io_outs_right[26] ,
    \ces_4_3_io_outs_right[25] ,
    \ces_4_3_io_outs_right[24] ,
    \ces_4_3_io_outs_right[23] ,
    \ces_4_3_io_outs_right[22] ,
    \ces_4_3_io_outs_right[21] ,
    \ces_4_3_io_outs_right[20] ,
    \ces_4_3_io_outs_right[19] ,
    \ces_4_3_io_outs_right[18] ,
    \ces_4_3_io_outs_right[17] ,
    \ces_4_3_io_outs_right[16] ,
    \ces_4_3_io_outs_right[15] ,
    \ces_4_3_io_outs_right[14] ,
    \ces_4_3_io_outs_right[13] ,
    \ces_4_3_io_outs_right[12] ,
    \ces_4_3_io_outs_right[11] ,
    \ces_4_3_io_outs_right[10] ,
    \ces_4_3_io_outs_right[9] ,
    \ces_4_3_io_outs_right[8] ,
    \ces_4_3_io_outs_right[7] ,
    \ces_4_3_io_outs_right[6] ,
    \ces_4_3_io_outs_right[5] ,
    \ces_4_3_io_outs_right[4] ,
    \ces_4_3_io_outs_right[3] ,
    \ces_4_3_io_outs_right[2] ,
    \ces_4_3_io_outs_right[1] ,
    \ces_4_3_io_outs_right[0] }),
    .io_ins_up({\ces_3_4_io_outs_up[63] ,
    \ces_3_4_io_outs_up[62] ,
    \ces_3_4_io_outs_up[61] ,
    \ces_3_4_io_outs_up[60] ,
    \ces_3_4_io_outs_up[59] ,
    \ces_3_4_io_outs_up[58] ,
    \ces_3_4_io_outs_up[57] ,
    \ces_3_4_io_outs_up[56] ,
    \ces_3_4_io_outs_up[55] ,
    \ces_3_4_io_outs_up[54] ,
    \ces_3_4_io_outs_up[53] ,
    \ces_3_4_io_outs_up[52] ,
    \ces_3_4_io_outs_up[51] ,
    \ces_3_4_io_outs_up[50] ,
    \ces_3_4_io_outs_up[49] ,
    \ces_3_4_io_outs_up[48] ,
    \ces_3_4_io_outs_up[47] ,
    \ces_3_4_io_outs_up[46] ,
    \ces_3_4_io_outs_up[45] ,
    \ces_3_4_io_outs_up[44] ,
    \ces_3_4_io_outs_up[43] ,
    \ces_3_4_io_outs_up[42] ,
    \ces_3_4_io_outs_up[41] ,
    \ces_3_4_io_outs_up[40] ,
    \ces_3_4_io_outs_up[39] ,
    \ces_3_4_io_outs_up[38] ,
    \ces_3_4_io_outs_up[37] ,
    \ces_3_4_io_outs_up[36] ,
    \ces_3_4_io_outs_up[35] ,
    \ces_3_4_io_outs_up[34] ,
    \ces_3_4_io_outs_up[33] ,
    \ces_3_4_io_outs_up[32] ,
    \ces_3_4_io_outs_up[31] ,
    \ces_3_4_io_outs_up[30] ,
    \ces_3_4_io_outs_up[29] ,
    \ces_3_4_io_outs_up[28] ,
    \ces_3_4_io_outs_up[27] ,
    \ces_3_4_io_outs_up[26] ,
    \ces_3_4_io_outs_up[25] ,
    \ces_3_4_io_outs_up[24] ,
    \ces_3_4_io_outs_up[23] ,
    \ces_3_4_io_outs_up[22] ,
    \ces_3_4_io_outs_up[21] ,
    \ces_3_4_io_outs_up[20] ,
    \ces_3_4_io_outs_up[19] ,
    \ces_3_4_io_outs_up[18] ,
    \ces_3_4_io_outs_up[17] ,
    \ces_3_4_io_outs_up[16] ,
    \ces_3_4_io_outs_up[15] ,
    \ces_3_4_io_outs_up[14] ,
    \ces_3_4_io_outs_up[13] ,
    \ces_3_4_io_outs_up[12] ,
    \ces_3_4_io_outs_up[11] ,
    \ces_3_4_io_outs_up[10] ,
    \ces_3_4_io_outs_up[9] ,
    \ces_3_4_io_outs_up[8] ,
    \ces_3_4_io_outs_up[7] ,
    \ces_3_4_io_outs_up[6] ,
    \ces_3_4_io_outs_up[5] ,
    \ces_3_4_io_outs_up[4] ,
    \ces_3_4_io_outs_up[3] ,
    \ces_3_4_io_outs_up[2] ,
    \ces_3_4_io_outs_up[1] ,
    \ces_3_4_io_outs_up[0] }),
    .io_outs_down({\ces_3_4_io_ins_down[63] ,
    \ces_3_4_io_ins_down[62] ,
    \ces_3_4_io_ins_down[61] ,
    \ces_3_4_io_ins_down[60] ,
    \ces_3_4_io_ins_down[59] ,
    \ces_3_4_io_ins_down[58] ,
    \ces_3_4_io_ins_down[57] ,
    \ces_3_4_io_ins_down[56] ,
    \ces_3_4_io_ins_down[55] ,
    \ces_3_4_io_ins_down[54] ,
    \ces_3_4_io_ins_down[53] ,
    \ces_3_4_io_ins_down[52] ,
    \ces_3_4_io_ins_down[51] ,
    \ces_3_4_io_ins_down[50] ,
    \ces_3_4_io_ins_down[49] ,
    \ces_3_4_io_ins_down[48] ,
    \ces_3_4_io_ins_down[47] ,
    \ces_3_4_io_ins_down[46] ,
    \ces_3_4_io_ins_down[45] ,
    \ces_3_4_io_ins_down[44] ,
    \ces_3_4_io_ins_down[43] ,
    \ces_3_4_io_ins_down[42] ,
    \ces_3_4_io_ins_down[41] ,
    \ces_3_4_io_ins_down[40] ,
    \ces_3_4_io_ins_down[39] ,
    \ces_3_4_io_ins_down[38] ,
    \ces_3_4_io_ins_down[37] ,
    \ces_3_4_io_ins_down[36] ,
    \ces_3_4_io_ins_down[35] ,
    \ces_3_4_io_ins_down[34] ,
    \ces_3_4_io_ins_down[33] ,
    \ces_3_4_io_ins_down[32] ,
    \ces_3_4_io_ins_down[31] ,
    \ces_3_4_io_ins_down[30] ,
    \ces_3_4_io_ins_down[29] ,
    \ces_3_4_io_ins_down[28] ,
    \ces_3_4_io_ins_down[27] ,
    \ces_3_4_io_ins_down[26] ,
    \ces_3_4_io_ins_down[25] ,
    \ces_3_4_io_ins_down[24] ,
    \ces_3_4_io_ins_down[23] ,
    \ces_3_4_io_ins_down[22] ,
    \ces_3_4_io_ins_down[21] ,
    \ces_3_4_io_ins_down[20] ,
    \ces_3_4_io_ins_down[19] ,
    \ces_3_4_io_ins_down[18] ,
    \ces_3_4_io_ins_down[17] ,
    \ces_3_4_io_ins_down[16] ,
    \ces_3_4_io_ins_down[15] ,
    \ces_3_4_io_ins_down[14] ,
    \ces_3_4_io_ins_down[13] ,
    \ces_3_4_io_ins_down[12] ,
    \ces_3_4_io_ins_down[11] ,
    \ces_3_4_io_ins_down[10] ,
    \ces_3_4_io_ins_down[9] ,
    \ces_3_4_io_ins_down[8] ,
    \ces_3_4_io_ins_down[7] ,
    \ces_3_4_io_ins_down[6] ,
    \ces_3_4_io_ins_down[5] ,
    \ces_3_4_io_ins_down[4] ,
    \ces_3_4_io_ins_down[3] ,
    \ces_3_4_io_ins_down[2] ,
    \ces_3_4_io_ins_down[1] ,
    \ces_3_4_io_ins_down[0] }),
    .io_outs_left({\ces_4_3_io_ins_left[63] ,
    \ces_4_3_io_ins_left[62] ,
    \ces_4_3_io_ins_left[61] ,
    \ces_4_3_io_ins_left[60] ,
    \ces_4_3_io_ins_left[59] ,
    \ces_4_3_io_ins_left[58] ,
    \ces_4_3_io_ins_left[57] ,
    \ces_4_3_io_ins_left[56] ,
    \ces_4_3_io_ins_left[55] ,
    \ces_4_3_io_ins_left[54] ,
    \ces_4_3_io_ins_left[53] ,
    \ces_4_3_io_ins_left[52] ,
    \ces_4_3_io_ins_left[51] ,
    \ces_4_3_io_ins_left[50] ,
    \ces_4_3_io_ins_left[49] ,
    \ces_4_3_io_ins_left[48] ,
    \ces_4_3_io_ins_left[47] ,
    \ces_4_3_io_ins_left[46] ,
    \ces_4_3_io_ins_left[45] ,
    \ces_4_3_io_ins_left[44] ,
    \ces_4_3_io_ins_left[43] ,
    \ces_4_3_io_ins_left[42] ,
    \ces_4_3_io_ins_left[41] ,
    \ces_4_3_io_ins_left[40] ,
    \ces_4_3_io_ins_left[39] ,
    \ces_4_3_io_ins_left[38] ,
    \ces_4_3_io_ins_left[37] ,
    \ces_4_3_io_ins_left[36] ,
    \ces_4_3_io_ins_left[35] ,
    \ces_4_3_io_ins_left[34] ,
    \ces_4_3_io_ins_left[33] ,
    \ces_4_3_io_ins_left[32] ,
    \ces_4_3_io_ins_left[31] ,
    \ces_4_3_io_ins_left[30] ,
    \ces_4_3_io_ins_left[29] ,
    \ces_4_3_io_ins_left[28] ,
    \ces_4_3_io_ins_left[27] ,
    \ces_4_3_io_ins_left[26] ,
    \ces_4_3_io_ins_left[25] ,
    \ces_4_3_io_ins_left[24] ,
    \ces_4_3_io_ins_left[23] ,
    \ces_4_3_io_ins_left[22] ,
    \ces_4_3_io_ins_left[21] ,
    \ces_4_3_io_ins_left[20] ,
    \ces_4_3_io_ins_left[19] ,
    \ces_4_3_io_ins_left[18] ,
    \ces_4_3_io_ins_left[17] ,
    \ces_4_3_io_ins_left[16] ,
    \ces_4_3_io_ins_left[15] ,
    \ces_4_3_io_ins_left[14] ,
    \ces_4_3_io_ins_left[13] ,
    \ces_4_3_io_ins_left[12] ,
    \ces_4_3_io_ins_left[11] ,
    \ces_4_3_io_ins_left[10] ,
    \ces_4_3_io_ins_left[9] ,
    \ces_4_3_io_ins_left[8] ,
    \ces_4_3_io_ins_left[7] ,
    \ces_4_3_io_ins_left[6] ,
    \ces_4_3_io_ins_left[5] ,
    \ces_4_3_io_ins_left[4] ,
    \ces_4_3_io_ins_left[3] ,
    \ces_4_3_io_ins_left[2] ,
    \ces_4_3_io_ins_left[1] ,
    \ces_4_3_io_ins_left[0] }),
    .io_outs_right({\ces_4_4_io_outs_right[63] ,
    \ces_4_4_io_outs_right[62] ,
    \ces_4_4_io_outs_right[61] ,
    \ces_4_4_io_outs_right[60] ,
    \ces_4_4_io_outs_right[59] ,
    \ces_4_4_io_outs_right[58] ,
    \ces_4_4_io_outs_right[57] ,
    \ces_4_4_io_outs_right[56] ,
    \ces_4_4_io_outs_right[55] ,
    \ces_4_4_io_outs_right[54] ,
    \ces_4_4_io_outs_right[53] ,
    \ces_4_4_io_outs_right[52] ,
    \ces_4_4_io_outs_right[51] ,
    \ces_4_4_io_outs_right[50] ,
    \ces_4_4_io_outs_right[49] ,
    \ces_4_4_io_outs_right[48] ,
    \ces_4_4_io_outs_right[47] ,
    \ces_4_4_io_outs_right[46] ,
    \ces_4_4_io_outs_right[45] ,
    \ces_4_4_io_outs_right[44] ,
    \ces_4_4_io_outs_right[43] ,
    \ces_4_4_io_outs_right[42] ,
    \ces_4_4_io_outs_right[41] ,
    \ces_4_4_io_outs_right[40] ,
    \ces_4_4_io_outs_right[39] ,
    \ces_4_4_io_outs_right[38] ,
    \ces_4_4_io_outs_right[37] ,
    \ces_4_4_io_outs_right[36] ,
    \ces_4_4_io_outs_right[35] ,
    \ces_4_4_io_outs_right[34] ,
    \ces_4_4_io_outs_right[33] ,
    \ces_4_4_io_outs_right[32] ,
    \ces_4_4_io_outs_right[31] ,
    \ces_4_4_io_outs_right[30] ,
    \ces_4_4_io_outs_right[29] ,
    \ces_4_4_io_outs_right[28] ,
    \ces_4_4_io_outs_right[27] ,
    \ces_4_4_io_outs_right[26] ,
    \ces_4_4_io_outs_right[25] ,
    \ces_4_4_io_outs_right[24] ,
    \ces_4_4_io_outs_right[23] ,
    \ces_4_4_io_outs_right[22] ,
    \ces_4_4_io_outs_right[21] ,
    \ces_4_4_io_outs_right[20] ,
    \ces_4_4_io_outs_right[19] ,
    \ces_4_4_io_outs_right[18] ,
    \ces_4_4_io_outs_right[17] ,
    \ces_4_4_io_outs_right[16] ,
    \ces_4_4_io_outs_right[15] ,
    \ces_4_4_io_outs_right[14] ,
    \ces_4_4_io_outs_right[13] ,
    \ces_4_4_io_outs_right[12] ,
    \ces_4_4_io_outs_right[11] ,
    \ces_4_4_io_outs_right[10] ,
    \ces_4_4_io_outs_right[9] ,
    \ces_4_4_io_outs_right[8] ,
    \ces_4_4_io_outs_right[7] ,
    \ces_4_4_io_outs_right[6] ,
    \ces_4_4_io_outs_right[5] ,
    \ces_4_4_io_outs_right[4] ,
    \ces_4_4_io_outs_right[3] ,
    \ces_4_4_io_outs_right[2] ,
    \ces_4_4_io_outs_right[1] ,
    \ces_4_4_io_outs_right[0] }),
    .io_outs_up({\ces_4_4_io_outs_up[63] ,
    \ces_4_4_io_outs_up[62] ,
    \ces_4_4_io_outs_up[61] ,
    \ces_4_4_io_outs_up[60] ,
    \ces_4_4_io_outs_up[59] ,
    \ces_4_4_io_outs_up[58] ,
    \ces_4_4_io_outs_up[57] ,
    \ces_4_4_io_outs_up[56] ,
    \ces_4_4_io_outs_up[55] ,
    \ces_4_4_io_outs_up[54] ,
    \ces_4_4_io_outs_up[53] ,
    \ces_4_4_io_outs_up[52] ,
    \ces_4_4_io_outs_up[51] ,
    \ces_4_4_io_outs_up[50] ,
    \ces_4_4_io_outs_up[49] ,
    \ces_4_4_io_outs_up[48] ,
    \ces_4_4_io_outs_up[47] ,
    \ces_4_4_io_outs_up[46] ,
    \ces_4_4_io_outs_up[45] ,
    \ces_4_4_io_outs_up[44] ,
    \ces_4_4_io_outs_up[43] ,
    \ces_4_4_io_outs_up[42] ,
    \ces_4_4_io_outs_up[41] ,
    \ces_4_4_io_outs_up[40] ,
    \ces_4_4_io_outs_up[39] ,
    \ces_4_4_io_outs_up[38] ,
    \ces_4_4_io_outs_up[37] ,
    \ces_4_4_io_outs_up[36] ,
    \ces_4_4_io_outs_up[35] ,
    \ces_4_4_io_outs_up[34] ,
    \ces_4_4_io_outs_up[33] ,
    \ces_4_4_io_outs_up[32] ,
    \ces_4_4_io_outs_up[31] ,
    \ces_4_4_io_outs_up[30] ,
    \ces_4_4_io_outs_up[29] ,
    \ces_4_4_io_outs_up[28] ,
    \ces_4_4_io_outs_up[27] ,
    \ces_4_4_io_outs_up[26] ,
    \ces_4_4_io_outs_up[25] ,
    \ces_4_4_io_outs_up[24] ,
    \ces_4_4_io_outs_up[23] ,
    \ces_4_4_io_outs_up[22] ,
    \ces_4_4_io_outs_up[21] ,
    \ces_4_4_io_outs_up[20] ,
    \ces_4_4_io_outs_up[19] ,
    \ces_4_4_io_outs_up[18] ,
    \ces_4_4_io_outs_up[17] ,
    \ces_4_4_io_outs_up[16] ,
    \ces_4_4_io_outs_up[15] ,
    \ces_4_4_io_outs_up[14] ,
    \ces_4_4_io_outs_up[13] ,
    \ces_4_4_io_outs_up[12] ,
    \ces_4_4_io_outs_up[11] ,
    \ces_4_4_io_outs_up[10] ,
    \ces_4_4_io_outs_up[9] ,
    \ces_4_4_io_outs_up[8] ,
    \ces_4_4_io_outs_up[7] ,
    \ces_4_4_io_outs_up[6] ,
    \ces_4_4_io_outs_up[5] ,
    \ces_4_4_io_outs_up[4] ,
    \ces_4_4_io_outs_up[3] ,
    \ces_4_4_io_outs_up[2] ,
    \ces_4_4_io_outs_up[1] ,
    \ces_4_4_io_outs_up[0] }));
 Element ces_4_5 (.clock(clknet_3_6_0_clock),
    .io_lsbIns_1(ces_4_4_io_lsbOuts_1),
    .io_lsbIns_2(ces_4_4_io_lsbOuts_2),
    .io_lsbIns_3(ces_4_4_io_lsbOuts_3),
    .io_lsbIns_4(ces_4_4_io_lsbOuts_4),
    .io_lsbIns_5(ces_4_4_io_lsbOuts_5),
    .io_lsbIns_6(ces_4_4_io_lsbOuts_6),
    .io_lsbIns_7(ces_4_4_io_lsbOuts_7),
    .io_lsbOuts_0(ces_4_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_5_io_lsbOuts_7),
    .io_ins_down({\ces_4_5_io_ins_down[63] ,
    \ces_4_5_io_ins_down[62] ,
    \ces_4_5_io_ins_down[61] ,
    \ces_4_5_io_ins_down[60] ,
    \ces_4_5_io_ins_down[59] ,
    \ces_4_5_io_ins_down[58] ,
    \ces_4_5_io_ins_down[57] ,
    \ces_4_5_io_ins_down[56] ,
    \ces_4_5_io_ins_down[55] ,
    \ces_4_5_io_ins_down[54] ,
    \ces_4_5_io_ins_down[53] ,
    \ces_4_5_io_ins_down[52] ,
    \ces_4_5_io_ins_down[51] ,
    \ces_4_5_io_ins_down[50] ,
    \ces_4_5_io_ins_down[49] ,
    \ces_4_5_io_ins_down[48] ,
    \ces_4_5_io_ins_down[47] ,
    \ces_4_5_io_ins_down[46] ,
    \ces_4_5_io_ins_down[45] ,
    \ces_4_5_io_ins_down[44] ,
    \ces_4_5_io_ins_down[43] ,
    \ces_4_5_io_ins_down[42] ,
    \ces_4_5_io_ins_down[41] ,
    \ces_4_5_io_ins_down[40] ,
    \ces_4_5_io_ins_down[39] ,
    \ces_4_5_io_ins_down[38] ,
    \ces_4_5_io_ins_down[37] ,
    \ces_4_5_io_ins_down[36] ,
    \ces_4_5_io_ins_down[35] ,
    \ces_4_5_io_ins_down[34] ,
    \ces_4_5_io_ins_down[33] ,
    \ces_4_5_io_ins_down[32] ,
    \ces_4_5_io_ins_down[31] ,
    \ces_4_5_io_ins_down[30] ,
    \ces_4_5_io_ins_down[29] ,
    \ces_4_5_io_ins_down[28] ,
    \ces_4_5_io_ins_down[27] ,
    \ces_4_5_io_ins_down[26] ,
    \ces_4_5_io_ins_down[25] ,
    \ces_4_5_io_ins_down[24] ,
    \ces_4_5_io_ins_down[23] ,
    \ces_4_5_io_ins_down[22] ,
    \ces_4_5_io_ins_down[21] ,
    \ces_4_5_io_ins_down[20] ,
    \ces_4_5_io_ins_down[19] ,
    \ces_4_5_io_ins_down[18] ,
    \ces_4_5_io_ins_down[17] ,
    \ces_4_5_io_ins_down[16] ,
    \ces_4_5_io_ins_down[15] ,
    \ces_4_5_io_ins_down[14] ,
    \ces_4_5_io_ins_down[13] ,
    \ces_4_5_io_ins_down[12] ,
    \ces_4_5_io_ins_down[11] ,
    \ces_4_5_io_ins_down[10] ,
    \ces_4_5_io_ins_down[9] ,
    \ces_4_5_io_ins_down[8] ,
    \ces_4_5_io_ins_down[7] ,
    \ces_4_5_io_ins_down[6] ,
    \ces_4_5_io_ins_down[5] ,
    \ces_4_5_io_ins_down[4] ,
    \ces_4_5_io_ins_down[3] ,
    \ces_4_5_io_ins_down[2] ,
    \ces_4_5_io_ins_down[1] ,
    \ces_4_5_io_ins_down[0] }),
    .io_ins_left({\ces_4_5_io_ins_left[63] ,
    \ces_4_5_io_ins_left[62] ,
    \ces_4_5_io_ins_left[61] ,
    \ces_4_5_io_ins_left[60] ,
    \ces_4_5_io_ins_left[59] ,
    \ces_4_5_io_ins_left[58] ,
    \ces_4_5_io_ins_left[57] ,
    \ces_4_5_io_ins_left[56] ,
    \ces_4_5_io_ins_left[55] ,
    \ces_4_5_io_ins_left[54] ,
    \ces_4_5_io_ins_left[53] ,
    \ces_4_5_io_ins_left[52] ,
    \ces_4_5_io_ins_left[51] ,
    \ces_4_5_io_ins_left[50] ,
    \ces_4_5_io_ins_left[49] ,
    \ces_4_5_io_ins_left[48] ,
    \ces_4_5_io_ins_left[47] ,
    \ces_4_5_io_ins_left[46] ,
    \ces_4_5_io_ins_left[45] ,
    \ces_4_5_io_ins_left[44] ,
    \ces_4_5_io_ins_left[43] ,
    \ces_4_5_io_ins_left[42] ,
    \ces_4_5_io_ins_left[41] ,
    \ces_4_5_io_ins_left[40] ,
    \ces_4_5_io_ins_left[39] ,
    \ces_4_5_io_ins_left[38] ,
    \ces_4_5_io_ins_left[37] ,
    \ces_4_5_io_ins_left[36] ,
    \ces_4_5_io_ins_left[35] ,
    \ces_4_5_io_ins_left[34] ,
    \ces_4_5_io_ins_left[33] ,
    \ces_4_5_io_ins_left[32] ,
    \ces_4_5_io_ins_left[31] ,
    \ces_4_5_io_ins_left[30] ,
    \ces_4_5_io_ins_left[29] ,
    \ces_4_5_io_ins_left[28] ,
    \ces_4_5_io_ins_left[27] ,
    \ces_4_5_io_ins_left[26] ,
    \ces_4_5_io_ins_left[25] ,
    \ces_4_5_io_ins_left[24] ,
    \ces_4_5_io_ins_left[23] ,
    \ces_4_5_io_ins_left[22] ,
    \ces_4_5_io_ins_left[21] ,
    \ces_4_5_io_ins_left[20] ,
    \ces_4_5_io_ins_left[19] ,
    \ces_4_5_io_ins_left[18] ,
    \ces_4_5_io_ins_left[17] ,
    \ces_4_5_io_ins_left[16] ,
    \ces_4_5_io_ins_left[15] ,
    \ces_4_5_io_ins_left[14] ,
    \ces_4_5_io_ins_left[13] ,
    \ces_4_5_io_ins_left[12] ,
    \ces_4_5_io_ins_left[11] ,
    \ces_4_5_io_ins_left[10] ,
    \ces_4_5_io_ins_left[9] ,
    \ces_4_5_io_ins_left[8] ,
    \ces_4_5_io_ins_left[7] ,
    \ces_4_5_io_ins_left[6] ,
    \ces_4_5_io_ins_left[5] ,
    \ces_4_5_io_ins_left[4] ,
    \ces_4_5_io_ins_left[3] ,
    \ces_4_5_io_ins_left[2] ,
    \ces_4_5_io_ins_left[1] ,
    \ces_4_5_io_ins_left[0] }),
    .io_ins_right({\ces_4_4_io_outs_right[63] ,
    \ces_4_4_io_outs_right[62] ,
    \ces_4_4_io_outs_right[61] ,
    \ces_4_4_io_outs_right[60] ,
    \ces_4_4_io_outs_right[59] ,
    \ces_4_4_io_outs_right[58] ,
    \ces_4_4_io_outs_right[57] ,
    \ces_4_4_io_outs_right[56] ,
    \ces_4_4_io_outs_right[55] ,
    \ces_4_4_io_outs_right[54] ,
    \ces_4_4_io_outs_right[53] ,
    \ces_4_4_io_outs_right[52] ,
    \ces_4_4_io_outs_right[51] ,
    \ces_4_4_io_outs_right[50] ,
    \ces_4_4_io_outs_right[49] ,
    \ces_4_4_io_outs_right[48] ,
    \ces_4_4_io_outs_right[47] ,
    \ces_4_4_io_outs_right[46] ,
    \ces_4_4_io_outs_right[45] ,
    \ces_4_4_io_outs_right[44] ,
    \ces_4_4_io_outs_right[43] ,
    \ces_4_4_io_outs_right[42] ,
    \ces_4_4_io_outs_right[41] ,
    \ces_4_4_io_outs_right[40] ,
    \ces_4_4_io_outs_right[39] ,
    \ces_4_4_io_outs_right[38] ,
    \ces_4_4_io_outs_right[37] ,
    \ces_4_4_io_outs_right[36] ,
    \ces_4_4_io_outs_right[35] ,
    \ces_4_4_io_outs_right[34] ,
    \ces_4_4_io_outs_right[33] ,
    \ces_4_4_io_outs_right[32] ,
    \ces_4_4_io_outs_right[31] ,
    \ces_4_4_io_outs_right[30] ,
    \ces_4_4_io_outs_right[29] ,
    \ces_4_4_io_outs_right[28] ,
    \ces_4_4_io_outs_right[27] ,
    \ces_4_4_io_outs_right[26] ,
    \ces_4_4_io_outs_right[25] ,
    \ces_4_4_io_outs_right[24] ,
    \ces_4_4_io_outs_right[23] ,
    \ces_4_4_io_outs_right[22] ,
    \ces_4_4_io_outs_right[21] ,
    \ces_4_4_io_outs_right[20] ,
    \ces_4_4_io_outs_right[19] ,
    \ces_4_4_io_outs_right[18] ,
    \ces_4_4_io_outs_right[17] ,
    \ces_4_4_io_outs_right[16] ,
    \ces_4_4_io_outs_right[15] ,
    \ces_4_4_io_outs_right[14] ,
    \ces_4_4_io_outs_right[13] ,
    \ces_4_4_io_outs_right[12] ,
    \ces_4_4_io_outs_right[11] ,
    \ces_4_4_io_outs_right[10] ,
    \ces_4_4_io_outs_right[9] ,
    \ces_4_4_io_outs_right[8] ,
    \ces_4_4_io_outs_right[7] ,
    \ces_4_4_io_outs_right[6] ,
    \ces_4_4_io_outs_right[5] ,
    \ces_4_4_io_outs_right[4] ,
    \ces_4_4_io_outs_right[3] ,
    \ces_4_4_io_outs_right[2] ,
    \ces_4_4_io_outs_right[1] ,
    \ces_4_4_io_outs_right[0] }),
    .io_ins_up({\ces_3_5_io_outs_up[63] ,
    \ces_3_5_io_outs_up[62] ,
    \ces_3_5_io_outs_up[61] ,
    \ces_3_5_io_outs_up[60] ,
    \ces_3_5_io_outs_up[59] ,
    \ces_3_5_io_outs_up[58] ,
    \ces_3_5_io_outs_up[57] ,
    \ces_3_5_io_outs_up[56] ,
    \ces_3_5_io_outs_up[55] ,
    \ces_3_5_io_outs_up[54] ,
    \ces_3_5_io_outs_up[53] ,
    \ces_3_5_io_outs_up[52] ,
    \ces_3_5_io_outs_up[51] ,
    \ces_3_5_io_outs_up[50] ,
    \ces_3_5_io_outs_up[49] ,
    \ces_3_5_io_outs_up[48] ,
    \ces_3_5_io_outs_up[47] ,
    \ces_3_5_io_outs_up[46] ,
    \ces_3_5_io_outs_up[45] ,
    \ces_3_5_io_outs_up[44] ,
    \ces_3_5_io_outs_up[43] ,
    \ces_3_5_io_outs_up[42] ,
    \ces_3_5_io_outs_up[41] ,
    \ces_3_5_io_outs_up[40] ,
    \ces_3_5_io_outs_up[39] ,
    \ces_3_5_io_outs_up[38] ,
    \ces_3_5_io_outs_up[37] ,
    \ces_3_5_io_outs_up[36] ,
    \ces_3_5_io_outs_up[35] ,
    \ces_3_5_io_outs_up[34] ,
    \ces_3_5_io_outs_up[33] ,
    \ces_3_5_io_outs_up[32] ,
    \ces_3_5_io_outs_up[31] ,
    \ces_3_5_io_outs_up[30] ,
    \ces_3_5_io_outs_up[29] ,
    \ces_3_5_io_outs_up[28] ,
    \ces_3_5_io_outs_up[27] ,
    \ces_3_5_io_outs_up[26] ,
    \ces_3_5_io_outs_up[25] ,
    \ces_3_5_io_outs_up[24] ,
    \ces_3_5_io_outs_up[23] ,
    \ces_3_5_io_outs_up[22] ,
    \ces_3_5_io_outs_up[21] ,
    \ces_3_5_io_outs_up[20] ,
    \ces_3_5_io_outs_up[19] ,
    \ces_3_5_io_outs_up[18] ,
    \ces_3_5_io_outs_up[17] ,
    \ces_3_5_io_outs_up[16] ,
    \ces_3_5_io_outs_up[15] ,
    \ces_3_5_io_outs_up[14] ,
    \ces_3_5_io_outs_up[13] ,
    \ces_3_5_io_outs_up[12] ,
    \ces_3_5_io_outs_up[11] ,
    \ces_3_5_io_outs_up[10] ,
    \ces_3_5_io_outs_up[9] ,
    \ces_3_5_io_outs_up[8] ,
    \ces_3_5_io_outs_up[7] ,
    \ces_3_5_io_outs_up[6] ,
    \ces_3_5_io_outs_up[5] ,
    \ces_3_5_io_outs_up[4] ,
    \ces_3_5_io_outs_up[3] ,
    \ces_3_5_io_outs_up[2] ,
    \ces_3_5_io_outs_up[1] ,
    \ces_3_5_io_outs_up[0] }),
    .io_outs_down({\ces_3_5_io_ins_down[63] ,
    \ces_3_5_io_ins_down[62] ,
    \ces_3_5_io_ins_down[61] ,
    \ces_3_5_io_ins_down[60] ,
    \ces_3_5_io_ins_down[59] ,
    \ces_3_5_io_ins_down[58] ,
    \ces_3_5_io_ins_down[57] ,
    \ces_3_5_io_ins_down[56] ,
    \ces_3_5_io_ins_down[55] ,
    \ces_3_5_io_ins_down[54] ,
    \ces_3_5_io_ins_down[53] ,
    \ces_3_5_io_ins_down[52] ,
    \ces_3_5_io_ins_down[51] ,
    \ces_3_5_io_ins_down[50] ,
    \ces_3_5_io_ins_down[49] ,
    \ces_3_5_io_ins_down[48] ,
    \ces_3_5_io_ins_down[47] ,
    \ces_3_5_io_ins_down[46] ,
    \ces_3_5_io_ins_down[45] ,
    \ces_3_5_io_ins_down[44] ,
    \ces_3_5_io_ins_down[43] ,
    \ces_3_5_io_ins_down[42] ,
    \ces_3_5_io_ins_down[41] ,
    \ces_3_5_io_ins_down[40] ,
    \ces_3_5_io_ins_down[39] ,
    \ces_3_5_io_ins_down[38] ,
    \ces_3_5_io_ins_down[37] ,
    \ces_3_5_io_ins_down[36] ,
    \ces_3_5_io_ins_down[35] ,
    \ces_3_5_io_ins_down[34] ,
    \ces_3_5_io_ins_down[33] ,
    \ces_3_5_io_ins_down[32] ,
    \ces_3_5_io_ins_down[31] ,
    \ces_3_5_io_ins_down[30] ,
    \ces_3_5_io_ins_down[29] ,
    \ces_3_5_io_ins_down[28] ,
    \ces_3_5_io_ins_down[27] ,
    \ces_3_5_io_ins_down[26] ,
    \ces_3_5_io_ins_down[25] ,
    \ces_3_5_io_ins_down[24] ,
    \ces_3_5_io_ins_down[23] ,
    \ces_3_5_io_ins_down[22] ,
    \ces_3_5_io_ins_down[21] ,
    \ces_3_5_io_ins_down[20] ,
    \ces_3_5_io_ins_down[19] ,
    \ces_3_5_io_ins_down[18] ,
    \ces_3_5_io_ins_down[17] ,
    \ces_3_5_io_ins_down[16] ,
    \ces_3_5_io_ins_down[15] ,
    \ces_3_5_io_ins_down[14] ,
    \ces_3_5_io_ins_down[13] ,
    \ces_3_5_io_ins_down[12] ,
    \ces_3_5_io_ins_down[11] ,
    \ces_3_5_io_ins_down[10] ,
    \ces_3_5_io_ins_down[9] ,
    \ces_3_5_io_ins_down[8] ,
    \ces_3_5_io_ins_down[7] ,
    \ces_3_5_io_ins_down[6] ,
    \ces_3_5_io_ins_down[5] ,
    \ces_3_5_io_ins_down[4] ,
    \ces_3_5_io_ins_down[3] ,
    \ces_3_5_io_ins_down[2] ,
    \ces_3_5_io_ins_down[1] ,
    \ces_3_5_io_ins_down[0] }),
    .io_outs_left({\ces_4_4_io_ins_left[63] ,
    \ces_4_4_io_ins_left[62] ,
    \ces_4_4_io_ins_left[61] ,
    \ces_4_4_io_ins_left[60] ,
    \ces_4_4_io_ins_left[59] ,
    \ces_4_4_io_ins_left[58] ,
    \ces_4_4_io_ins_left[57] ,
    \ces_4_4_io_ins_left[56] ,
    \ces_4_4_io_ins_left[55] ,
    \ces_4_4_io_ins_left[54] ,
    \ces_4_4_io_ins_left[53] ,
    \ces_4_4_io_ins_left[52] ,
    \ces_4_4_io_ins_left[51] ,
    \ces_4_4_io_ins_left[50] ,
    \ces_4_4_io_ins_left[49] ,
    \ces_4_4_io_ins_left[48] ,
    \ces_4_4_io_ins_left[47] ,
    \ces_4_4_io_ins_left[46] ,
    \ces_4_4_io_ins_left[45] ,
    \ces_4_4_io_ins_left[44] ,
    \ces_4_4_io_ins_left[43] ,
    \ces_4_4_io_ins_left[42] ,
    \ces_4_4_io_ins_left[41] ,
    \ces_4_4_io_ins_left[40] ,
    \ces_4_4_io_ins_left[39] ,
    \ces_4_4_io_ins_left[38] ,
    \ces_4_4_io_ins_left[37] ,
    \ces_4_4_io_ins_left[36] ,
    \ces_4_4_io_ins_left[35] ,
    \ces_4_4_io_ins_left[34] ,
    \ces_4_4_io_ins_left[33] ,
    \ces_4_4_io_ins_left[32] ,
    \ces_4_4_io_ins_left[31] ,
    \ces_4_4_io_ins_left[30] ,
    \ces_4_4_io_ins_left[29] ,
    \ces_4_4_io_ins_left[28] ,
    \ces_4_4_io_ins_left[27] ,
    \ces_4_4_io_ins_left[26] ,
    \ces_4_4_io_ins_left[25] ,
    \ces_4_4_io_ins_left[24] ,
    \ces_4_4_io_ins_left[23] ,
    \ces_4_4_io_ins_left[22] ,
    \ces_4_4_io_ins_left[21] ,
    \ces_4_4_io_ins_left[20] ,
    \ces_4_4_io_ins_left[19] ,
    \ces_4_4_io_ins_left[18] ,
    \ces_4_4_io_ins_left[17] ,
    \ces_4_4_io_ins_left[16] ,
    \ces_4_4_io_ins_left[15] ,
    \ces_4_4_io_ins_left[14] ,
    \ces_4_4_io_ins_left[13] ,
    \ces_4_4_io_ins_left[12] ,
    \ces_4_4_io_ins_left[11] ,
    \ces_4_4_io_ins_left[10] ,
    \ces_4_4_io_ins_left[9] ,
    \ces_4_4_io_ins_left[8] ,
    \ces_4_4_io_ins_left[7] ,
    \ces_4_4_io_ins_left[6] ,
    \ces_4_4_io_ins_left[5] ,
    \ces_4_4_io_ins_left[4] ,
    \ces_4_4_io_ins_left[3] ,
    \ces_4_4_io_ins_left[2] ,
    \ces_4_4_io_ins_left[1] ,
    \ces_4_4_io_ins_left[0] }),
    .io_outs_right({\ces_4_5_io_outs_right[63] ,
    \ces_4_5_io_outs_right[62] ,
    \ces_4_5_io_outs_right[61] ,
    \ces_4_5_io_outs_right[60] ,
    \ces_4_5_io_outs_right[59] ,
    \ces_4_5_io_outs_right[58] ,
    \ces_4_5_io_outs_right[57] ,
    \ces_4_5_io_outs_right[56] ,
    \ces_4_5_io_outs_right[55] ,
    \ces_4_5_io_outs_right[54] ,
    \ces_4_5_io_outs_right[53] ,
    \ces_4_5_io_outs_right[52] ,
    \ces_4_5_io_outs_right[51] ,
    \ces_4_5_io_outs_right[50] ,
    \ces_4_5_io_outs_right[49] ,
    \ces_4_5_io_outs_right[48] ,
    \ces_4_5_io_outs_right[47] ,
    \ces_4_5_io_outs_right[46] ,
    \ces_4_5_io_outs_right[45] ,
    \ces_4_5_io_outs_right[44] ,
    \ces_4_5_io_outs_right[43] ,
    \ces_4_5_io_outs_right[42] ,
    \ces_4_5_io_outs_right[41] ,
    \ces_4_5_io_outs_right[40] ,
    \ces_4_5_io_outs_right[39] ,
    \ces_4_5_io_outs_right[38] ,
    \ces_4_5_io_outs_right[37] ,
    \ces_4_5_io_outs_right[36] ,
    \ces_4_5_io_outs_right[35] ,
    \ces_4_5_io_outs_right[34] ,
    \ces_4_5_io_outs_right[33] ,
    \ces_4_5_io_outs_right[32] ,
    \ces_4_5_io_outs_right[31] ,
    \ces_4_5_io_outs_right[30] ,
    \ces_4_5_io_outs_right[29] ,
    \ces_4_5_io_outs_right[28] ,
    \ces_4_5_io_outs_right[27] ,
    \ces_4_5_io_outs_right[26] ,
    \ces_4_5_io_outs_right[25] ,
    \ces_4_5_io_outs_right[24] ,
    \ces_4_5_io_outs_right[23] ,
    \ces_4_5_io_outs_right[22] ,
    \ces_4_5_io_outs_right[21] ,
    \ces_4_5_io_outs_right[20] ,
    \ces_4_5_io_outs_right[19] ,
    \ces_4_5_io_outs_right[18] ,
    \ces_4_5_io_outs_right[17] ,
    \ces_4_5_io_outs_right[16] ,
    \ces_4_5_io_outs_right[15] ,
    \ces_4_5_io_outs_right[14] ,
    \ces_4_5_io_outs_right[13] ,
    \ces_4_5_io_outs_right[12] ,
    \ces_4_5_io_outs_right[11] ,
    \ces_4_5_io_outs_right[10] ,
    \ces_4_5_io_outs_right[9] ,
    \ces_4_5_io_outs_right[8] ,
    \ces_4_5_io_outs_right[7] ,
    \ces_4_5_io_outs_right[6] ,
    \ces_4_5_io_outs_right[5] ,
    \ces_4_5_io_outs_right[4] ,
    \ces_4_5_io_outs_right[3] ,
    \ces_4_5_io_outs_right[2] ,
    \ces_4_5_io_outs_right[1] ,
    \ces_4_5_io_outs_right[0] }),
    .io_outs_up({\ces_4_5_io_outs_up[63] ,
    \ces_4_5_io_outs_up[62] ,
    \ces_4_5_io_outs_up[61] ,
    \ces_4_5_io_outs_up[60] ,
    \ces_4_5_io_outs_up[59] ,
    \ces_4_5_io_outs_up[58] ,
    \ces_4_5_io_outs_up[57] ,
    \ces_4_5_io_outs_up[56] ,
    \ces_4_5_io_outs_up[55] ,
    \ces_4_5_io_outs_up[54] ,
    \ces_4_5_io_outs_up[53] ,
    \ces_4_5_io_outs_up[52] ,
    \ces_4_5_io_outs_up[51] ,
    \ces_4_5_io_outs_up[50] ,
    \ces_4_5_io_outs_up[49] ,
    \ces_4_5_io_outs_up[48] ,
    \ces_4_5_io_outs_up[47] ,
    \ces_4_5_io_outs_up[46] ,
    \ces_4_5_io_outs_up[45] ,
    \ces_4_5_io_outs_up[44] ,
    \ces_4_5_io_outs_up[43] ,
    \ces_4_5_io_outs_up[42] ,
    \ces_4_5_io_outs_up[41] ,
    \ces_4_5_io_outs_up[40] ,
    \ces_4_5_io_outs_up[39] ,
    \ces_4_5_io_outs_up[38] ,
    \ces_4_5_io_outs_up[37] ,
    \ces_4_5_io_outs_up[36] ,
    \ces_4_5_io_outs_up[35] ,
    \ces_4_5_io_outs_up[34] ,
    \ces_4_5_io_outs_up[33] ,
    \ces_4_5_io_outs_up[32] ,
    \ces_4_5_io_outs_up[31] ,
    \ces_4_5_io_outs_up[30] ,
    \ces_4_5_io_outs_up[29] ,
    \ces_4_5_io_outs_up[28] ,
    \ces_4_5_io_outs_up[27] ,
    \ces_4_5_io_outs_up[26] ,
    \ces_4_5_io_outs_up[25] ,
    \ces_4_5_io_outs_up[24] ,
    \ces_4_5_io_outs_up[23] ,
    \ces_4_5_io_outs_up[22] ,
    \ces_4_5_io_outs_up[21] ,
    \ces_4_5_io_outs_up[20] ,
    \ces_4_5_io_outs_up[19] ,
    \ces_4_5_io_outs_up[18] ,
    \ces_4_5_io_outs_up[17] ,
    \ces_4_5_io_outs_up[16] ,
    \ces_4_5_io_outs_up[15] ,
    \ces_4_5_io_outs_up[14] ,
    \ces_4_5_io_outs_up[13] ,
    \ces_4_5_io_outs_up[12] ,
    \ces_4_5_io_outs_up[11] ,
    \ces_4_5_io_outs_up[10] ,
    \ces_4_5_io_outs_up[9] ,
    \ces_4_5_io_outs_up[8] ,
    \ces_4_5_io_outs_up[7] ,
    \ces_4_5_io_outs_up[6] ,
    \ces_4_5_io_outs_up[5] ,
    \ces_4_5_io_outs_up[4] ,
    \ces_4_5_io_outs_up[3] ,
    \ces_4_5_io_outs_up[2] ,
    \ces_4_5_io_outs_up[1] ,
    \ces_4_5_io_outs_up[0] }));
 Element ces_4_6 (.clock(clknet_3_6_0_clock),
    .io_lsbIns_1(ces_4_5_io_lsbOuts_1),
    .io_lsbIns_2(ces_4_5_io_lsbOuts_2),
    .io_lsbIns_3(ces_4_5_io_lsbOuts_3),
    .io_lsbIns_4(ces_4_5_io_lsbOuts_4),
    .io_lsbIns_5(ces_4_5_io_lsbOuts_5),
    .io_lsbIns_6(ces_4_5_io_lsbOuts_6),
    .io_lsbIns_7(ces_4_5_io_lsbOuts_7),
    .io_lsbOuts_0(ces_4_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_6_io_lsbOuts_7),
    .io_ins_down({\ces_4_6_io_ins_down[63] ,
    \ces_4_6_io_ins_down[62] ,
    \ces_4_6_io_ins_down[61] ,
    \ces_4_6_io_ins_down[60] ,
    \ces_4_6_io_ins_down[59] ,
    \ces_4_6_io_ins_down[58] ,
    \ces_4_6_io_ins_down[57] ,
    \ces_4_6_io_ins_down[56] ,
    \ces_4_6_io_ins_down[55] ,
    \ces_4_6_io_ins_down[54] ,
    \ces_4_6_io_ins_down[53] ,
    \ces_4_6_io_ins_down[52] ,
    \ces_4_6_io_ins_down[51] ,
    \ces_4_6_io_ins_down[50] ,
    \ces_4_6_io_ins_down[49] ,
    \ces_4_6_io_ins_down[48] ,
    \ces_4_6_io_ins_down[47] ,
    \ces_4_6_io_ins_down[46] ,
    \ces_4_6_io_ins_down[45] ,
    \ces_4_6_io_ins_down[44] ,
    \ces_4_6_io_ins_down[43] ,
    \ces_4_6_io_ins_down[42] ,
    \ces_4_6_io_ins_down[41] ,
    \ces_4_6_io_ins_down[40] ,
    \ces_4_6_io_ins_down[39] ,
    \ces_4_6_io_ins_down[38] ,
    \ces_4_6_io_ins_down[37] ,
    \ces_4_6_io_ins_down[36] ,
    \ces_4_6_io_ins_down[35] ,
    \ces_4_6_io_ins_down[34] ,
    \ces_4_6_io_ins_down[33] ,
    \ces_4_6_io_ins_down[32] ,
    \ces_4_6_io_ins_down[31] ,
    \ces_4_6_io_ins_down[30] ,
    \ces_4_6_io_ins_down[29] ,
    \ces_4_6_io_ins_down[28] ,
    \ces_4_6_io_ins_down[27] ,
    \ces_4_6_io_ins_down[26] ,
    \ces_4_6_io_ins_down[25] ,
    \ces_4_6_io_ins_down[24] ,
    \ces_4_6_io_ins_down[23] ,
    \ces_4_6_io_ins_down[22] ,
    \ces_4_6_io_ins_down[21] ,
    \ces_4_6_io_ins_down[20] ,
    \ces_4_6_io_ins_down[19] ,
    \ces_4_6_io_ins_down[18] ,
    \ces_4_6_io_ins_down[17] ,
    \ces_4_6_io_ins_down[16] ,
    \ces_4_6_io_ins_down[15] ,
    \ces_4_6_io_ins_down[14] ,
    \ces_4_6_io_ins_down[13] ,
    \ces_4_6_io_ins_down[12] ,
    \ces_4_6_io_ins_down[11] ,
    \ces_4_6_io_ins_down[10] ,
    \ces_4_6_io_ins_down[9] ,
    \ces_4_6_io_ins_down[8] ,
    \ces_4_6_io_ins_down[7] ,
    \ces_4_6_io_ins_down[6] ,
    \ces_4_6_io_ins_down[5] ,
    \ces_4_6_io_ins_down[4] ,
    \ces_4_6_io_ins_down[3] ,
    \ces_4_6_io_ins_down[2] ,
    \ces_4_6_io_ins_down[1] ,
    \ces_4_6_io_ins_down[0] }),
    .io_ins_left({\ces_4_6_io_ins_left[63] ,
    \ces_4_6_io_ins_left[62] ,
    \ces_4_6_io_ins_left[61] ,
    \ces_4_6_io_ins_left[60] ,
    \ces_4_6_io_ins_left[59] ,
    \ces_4_6_io_ins_left[58] ,
    \ces_4_6_io_ins_left[57] ,
    \ces_4_6_io_ins_left[56] ,
    \ces_4_6_io_ins_left[55] ,
    \ces_4_6_io_ins_left[54] ,
    \ces_4_6_io_ins_left[53] ,
    \ces_4_6_io_ins_left[52] ,
    \ces_4_6_io_ins_left[51] ,
    \ces_4_6_io_ins_left[50] ,
    \ces_4_6_io_ins_left[49] ,
    \ces_4_6_io_ins_left[48] ,
    \ces_4_6_io_ins_left[47] ,
    \ces_4_6_io_ins_left[46] ,
    \ces_4_6_io_ins_left[45] ,
    \ces_4_6_io_ins_left[44] ,
    \ces_4_6_io_ins_left[43] ,
    \ces_4_6_io_ins_left[42] ,
    \ces_4_6_io_ins_left[41] ,
    \ces_4_6_io_ins_left[40] ,
    \ces_4_6_io_ins_left[39] ,
    \ces_4_6_io_ins_left[38] ,
    \ces_4_6_io_ins_left[37] ,
    \ces_4_6_io_ins_left[36] ,
    \ces_4_6_io_ins_left[35] ,
    \ces_4_6_io_ins_left[34] ,
    \ces_4_6_io_ins_left[33] ,
    \ces_4_6_io_ins_left[32] ,
    \ces_4_6_io_ins_left[31] ,
    \ces_4_6_io_ins_left[30] ,
    \ces_4_6_io_ins_left[29] ,
    \ces_4_6_io_ins_left[28] ,
    \ces_4_6_io_ins_left[27] ,
    \ces_4_6_io_ins_left[26] ,
    \ces_4_6_io_ins_left[25] ,
    \ces_4_6_io_ins_left[24] ,
    \ces_4_6_io_ins_left[23] ,
    \ces_4_6_io_ins_left[22] ,
    \ces_4_6_io_ins_left[21] ,
    \ces_4_6_io_ins_left[20] ,
    \ces_4_6_io_ins_left[19] ,
    \ces_4_6_io_ins_left[18] ,
    \ces_4_6_io_ins_left[17] ,
    \ces_4_6_io_ins_left[16] ,
    \ces_4_6_io_ins_left[15] ,
    \ces_4_6_io_ins_left[14] ,
    \ces_4_6_io_ins_left[13] ,
    \ces_4_6_io_ins_left[12] ,
    \ces_4_6_io_ins_left[11] ,
    \ces_4_6_io_ins_left[10] ,
    \ces_4_6_io_ins_left[9] ,
    \ces_4_6_io_ins_left[8] ,
    \ces_4_6_io_ins_left[7] ,
    \ces_4_6_io_ins_left[6] ,
    \ces_4_6_io_ins_left[5] ,
    \ces_4_6_io_ins_left[4] ,
    \ces_4_6_io_ins_left[3] ,
    \ces_4_6_io_ins_left[2] ,
    \ces_4_6_io_ins_left[1] ,
    \ces_4_6_io_ins_left[0] }),
    .io_ins_right({\ces_4_5_io_outs_right[63] ,
    \ces_4_5_io_outs_right[62] ,
    \ces_4_5_io_outs_right[61] ,
    \ces_4_5_io_outs_right[60] ,
    \ces_4_5_io_outs_right[59] ,
    \ces_4_5_io_outs_right[58] ,
    \ces_4_5_io_outs_right[57] ,
    \ces_4_5_io_outs_right[56] ,
    \ces_4_5_io_outs_right[55] ,
    \ces_4_5_io_outs_right[54] ,
    \ces_4_5_io_outs_right[53] ,
    \ces_4_5_io_outs_right[52] ,
    \ces_4_5_io_outs_right[51] ,
    \ces_4_5_io_outs_right[50] ,
    \ces_4_5_io_outs_right[49] ,
    \ces_4_5_io_outs_right[48] ,
    \ces_4_5_io_outs_right[47] ,
    \ces_4_5_io_outs_right[46] ,
    \ces_4_5_io_outs_right[45] ,
    \ces_4_5_io_outs_right[44] ,
    \ces_4_5_io_outs_right[43] ,
    \ces_4_5_io_outs_right[42] ,
    \ces_4_5_io_outs_right[41] ,
    \ces_4_5_io_outs_right[40] ,
    \ces_4_5_io_outs_right[39] ,
    \ces_4_5_io_outs_right[38] ,
    \ces_4_5_io_outs_right[37] ,
    \ces_4_5_io_outs_right[36] ,
    \ces_4_5_io_outs_right[35] ,
    \ces_4_5_io_outs_right[34] ,
    \ces_4_5_io_outs_right[33] ,
    \ces_4_5_io_outs_right[32] ,
    \ces_4_5_io_outs_right[31] ,
    \ces_4_5_io_outs_right[30] ,
    \ces_4_5_io_outs_right[29] ,
    \ces_4_5_io_outs_right[28] ,
    \ces_4_5_io_outs_right[27] ,
    \ces_4_5_io_outs_right[26] ,
    \ces_4_5_io_outs_right[25] ,
    \ces_4_5_io_outs_right[24] ,
    \ces_4_5_io_outs_right[23] ,
    \ces_4_5_io_outs_right[22] ,
    \ces_4_5_io_outs_right[21] ,
    \ces_4_5_io_outs_right[20] ,
    \ces_4_5_io_outs_right[19] ,
    \ces_4_5_io_outs_right[18] ,
    \ces_4_5_io_outs_right[17] ,
    \ces_4_5_io_outs_right[16] ,
    \ces_4_5_io_outs_right[15] ,
    \ces_4_5_io_outs_right[14] ,
    \ces_4_5_io_outs_right[13] ,
    \ces_4_5_io_outs_right[12] ,
    \ces_4_5_io_outs_right[11] ,
    \ces_4_5_io_outs_right[10] ,
    \ces_4_5_io_outs_right[9] ,
    \ces_4_5_io_outs_right[8] ,
    \ces_4_5_io_outs_right[7] ,
    \ces_4_5_io_outs_right[6] ,
    \ces_4_5_io_outs_right[5] ,
    \ces_4_5_io_outs_right[4] ,
    \ces_4_5_io_outs_right[3] ,
    \ces_4_5_io_outs_right[2] ,
    \ces_4_5_io_outs_right[1] ,
    \ces_4_5_io_outs_right[0] }),
    .io_ins_up({\ces_3_6_io_outs_up[63] ,
    \ces_3_6_io_outs_up[62] ,
    \ces_3_6_io_outs_up[61] ,
    \ces_3_6_io_outs_up[60] ,
    \ces_3_6_io_outs_up[59] ,
    \ces_3_6_io_outs_up[58] ,
    \ces_3_6_io_outs_up[57] ,
    \ces_3_6_io_outs_up[56] ,
    \ces_3_6_io_outs_up[55] ,
    \ces_3_6_io_outs_up[54] ,
    \ces_3_6_io_outs_up[53] ,
    \ces_3_6_io_outs_up[52] ,
    \ces_3_6_io_outs_up[51] ,
    \ces_3_6_io_outs_up[50] ,
    \ces_3_6_io_outs_up[49] ,
    \ces_3_6_io_outs_up[48] ,
    \ces_3_6_io_outs_up[47] ,
    \ces_3_6_io_outs_up[46] ,
    \ces_3_6_io_outs_up[45] ,
    \ces_3_6_io_outs_up[44] ,
    \ces_3_6_io_outs_up[43] ,
    \ces_3_6_io_outs_up[42] ,
    \ces_3_6_io_outs_up[41] ,
    \ces_3_6_io_outs_up[40] ,
    \ces_3_6_io_outs_up[39] ,
    \ces_3_6_io_outs_up[38] ,
    \ces_3_6_io_outs_up[37] ,
    \ces_3_6_io_outs_up[36] ,
    \ces_3_6_io_outs_up[35] ,
    \ces_3_6_io_outs_up[34] ,
    \ces_3_6_io_outs_up[33] ,
    \ces_3_6_io_outs_up[32] ,
    \ces_3_6_io_outs_up[31] ,
    \ces_3_6_io_outs_up[30] ,
    \ces_3_6_io_outs_up[29] ,
    \ces_3_6_io_outs_up[28] ,
    \ces_3_6_io_outs_up[27] ,
    \ces_3_6_io_outs_up[26] ,
    \ces_3_6_io_outs_up[25] ,
    \ces_3_6_io_outs_up[24] ,
    \ces_3_6_io_outs_up[23] ,
    \ces_3_6_io_outs_up[22] ,
    \ces_3_6_io_outs_up[21] ,
    \ces_3_6_io_outs_up[20] ,
    \ces_3_6_io_outs_up[19] ,
    \ces_3_6_io_outs_up[18] ,
    \ces_3_6_io_outs_up[17] ,
    \ces_3_6_io_outs_up[16] ,
    \ces_3_6_io_outs_up[15] ,
    \ces_3_6_io_outs_up[14] ,
    \ces_3_6_io_outs_up[13] ,
    \ces_3_6_io_outs_up[12] ,
    \ces_3_6_io_outs_up[11] ,
    \ces_3_6_io_outs_up[10] ,
    \ces_3_6_io_outs_up[9] ,
    \ces_3_6_io_outs_up[8] ,
    \ces_3_6_io_outs_up[7] ,
    \ces_3_6_io_outs_up[6] ,
    \ces_3_6_io_outs_up[5] ,
    \ces_3_6_io_outs_up[4] ,
    \ces_3_6_io_outs_up[3] ,
    \ces_3_6_io_outs_up[2] ,
    \ces_3_6_io_outs_up[1] ,
    \ces_3_6_io_outs_up[0] }),
    .io_outs_down({\ces_3_6_io_ins_down[63] ,
    \ces_3_6_io_ins_down[62] ,
    \ces_3_6_io_ins_down[61] ,
    \ces_3_6_io_ins_down[60] ,
    \ces_3_6_io_ins_down[59] ,
    \ces_3_6_io_ins_down[58] ,
    \ces_3_6_io_ins_down[57] ,
    \ces_3_6_io_ins_down[56] ,
    \ces_3_6_io_ins_down[55] ,
    \ces_3_6_io_ins_down[54] ,
    \ces_3_6_io_ins_down[53] ,
    \ces_3_6_io_ins_down[52] ,
    \ces_3_6_io_ins_down[51] ,
    \ces_3_6_io_ins_down[50] ,
    \ces_3_6_io_ins_down[49] ,
    \ces_3_6_io_ins_down[48] ,
    \ces_3_6_io_ins_down[47] ,
    \ces_3_6_io_ins_down[46] ,
    \ces_3_6_io_ins_down[45] ,
    \ces_3_6_io_ins_down[44] ,
    \ces_3_6_io_ins_down[43] ,
    \ces_3_6_io_ins_down[42] ,
    \ces_3_6_io_ins_down[41] ,
    \ces_3_6_io_ins_down[40] ,
    \ces_3_6_io_ins_down[39] ,
    \ces_3_6_io_ins_down[38] ,
    \ces_3_6_io_ins_down[37] ,
    \ces_3_6_io_ins_down[36] ,
    \ces_3_6_io_ins_down[35] ,
    \ces_3_6_io_ins_down[34] ,
    \ces_3_6_io_ins_down[33] ,
    \ces_3_6_io_ins_down[32] ,
    \ces_3_6_io_ins_down[31] ,
    \ces_3_6_io_ins_down[30] ,
    \ces_3_6_io_ins_down[29] ,
    \ces_3_6_io_ins_down[28] ,
    \ces_3_6_io_ins_down[27] ,
    \ces_3_6_io_ins_down[26] ,
    \ces_3_6_io_ins_down[25] ,
    \ces_3_6_io_ins_down[24] ,
    \ces_3_6_io_ins_down[23] ,
    \ces_3_6_io_ins_down[22] ,
    \ces_3_6_io_ins_down[21] ,
    \ces_3_6_io_ins_down[20] ,
    \ces_3_6_io_ins_down[19] ,
    \ces_3_6_io_ins_down[18] ,
    \ces_3_6_io_ins_down[17] ,
    \ces_3_6_io_ins_down[16] ,
    \ces_3_6_io_ins_down[15] ,
    \ces_3_6_io_ins_down[14] ,
    \ces_3_6_io_ins_down[13] ,
    \ces_3_6_io_ins_down[12] ,
    \ces_3_6_io_ins_down[11] ,
    \ces_3_6_io_ins_down[10] ,
    \ces_3_6_io_ins_down[9] ,
    \ces_3_6_io_ins_down[8] ,
    \ces_3_6_io_ins_down[7] ,
    \ces_3_6_io_ins_down[6] ,
    \ces_3_6_io_ins_down[5] ,
    \ces_3_6_io_ins_down[4] ,
    \ces_3_6_io_ins_down[3] ,
    \ces_3_6_io_ins_down[2] ,
    \ces_3_6_io_ins_down[1] ,
    \ces_3_6_io_ins_down[0] }),
    .io_outs_left({\ces_4_5_io_ins_left[63] ,
    \ces_4_5_io_ins_left[62] ,
    \ces_4_5_io_ins_left[61] ,
    \ces_4_5_io_ins_left[60] ,
    \ces_4_5_io_ins_left[59] ,
    \ces_4_5_io_ins_left[58] ,
    \ces_4_5_io_ins_left[57] ,
    \ces_4_5_io_ins_left[56] ,
    \ces_4_5_io_ins_left[55] ,
    \ces_4_5_io_ins_left[54] ,
    \ces_4_5_io_ins_left[53] ,
    \ces_4_5_io_ins_left[52] ,
    \ces_4_5_io_ins_left[51] ,
    \ces_4_5_io_ins_left[50] ,
    \ces_4_5_io_ins_left[49] ,
    \ces_4_5_io_ins_left[48] ,
    \ces_4_5_io_ins_left[47] ,
    \ces_4_5_io_ins_left[46] ,
    \ces_4_5_io_ins_left[45] ,
    \ces_4_5_io_ins_left[44] ,
    \ces_4_5_io_ins_left[43] ,
    \ces_4_5_io_ins_left[42] ,
    \ces_4_5_io_ins_left[41] ,
    \ces_4_5_io_ins_left[40] ,
    \ces_4_5_io_ins_left[39] ,
    \ces_4_5_io_ins_left[38] ,
    \ces_4_5_io_ins_left[37] ,
    \ces_4_5_io_ins_left[36] ,
    \ces_4_5_io_ins_left[35] ,
    \ces_4_5_io_ins_left[34] ,
    \ces_4_5_io_ins_left[33] ,
    \ces_4_5_io_ins_left[32] ,
    \ces_4_5_io_ins_left[31] ,
    \ces_4_5_io_ins_left[30] ,
    \ces_4_5_io_ins_left[29] ,
    \ces_4_5_io_ins_left[28] ,
    \ces_4_5_io_ins_left[27] ,
    \ces_4_5_io_ins_left[26] ,
    \ces_4_5_io_ins_left[25] ,
    \ces_4_5_io_ins_left[24] ,
    \ces_4_5_io_ins_left[23] ,
    \ces_4_5_io_ins_left[22] ,
    \ces_4_5_io_ins_left[21] ,
    \ces_4_5_io_ins_left[20] ,
    \ces_4_5_io_ins_left[19] ,
    \ces_4_5_io_ins_left[18] ,
    \ces_4_5_io_ins_left[17] ,
    \ces_4_5_io_ins_left[16] ,
    \ces_4_5_io_ins_left[15] ,
    \ces_4_5_io_ins_left[14] ,
    \ces_4_5_io_ins_left[13] ,
    \ces_4_5_io_ins_left[12] ,
    \ces_4_5_io_ins_left[11] ,
    \ces_4_5_io_ins_left[10] ,
    \ces_4_5_io_ins_left[9] ,
    \ces_4_5_io_ins_left[8] ,
    \ces_4_5_io_ins_left[7] ,
    \ces_4_5_io_ins_left[6] ,
    \ces_4_5_io_ins_left[5] ,
    \ces_4_5_io_ins_left[4] ,
    \ces_4_5_io_ins_left[3] ,
    \ces_4_5_io_ins_left[2] ,
    \ces_4_5_io_ins_left[1] ,
    \ces_4_5_io_ins_left[0] }),
    .io_outs_right({\ces_4_6_io_outs_right[63] ,
    \ces_4_6_io_outs_right[62] ,
    \ces_4_6_io_outs_right[61] ,
    \ces_4_6_io_outs_right[60] ,
    \ces_4_6_io_outs_right[59] ,
    \ces_4_6_io_outs_right[58] ,
    \ces_4_6_io_outs_right[57] ,
    \ces_4_6_io_outs_right[56] ,
    \ces_4_6_io_outs_right[55] ,
    \ces_4_6_io_outs_right[54] ,
    \ces_4_6_io_outs_right[53] ,
    \ces_4_6_io_outs_right[52] ,
    \ces_4_6_io_outs_right[51] ,
    \ces_4_6_io_outs_right[50] ,
    \ces_4_6_io_outs_right[49] ,
    \ces_4_6_io_outs_right[48] ,
    \ces_4_6_io_outs_right[47] ,
    \ces_4_6_io_outs_right[46] ,
    \ces_4_6_io_outs_right[45] ,
    \ces_4_6_io_outs_right[44] ,
    \ces_4_6_io_outs_right[43] ,
    \ces_4_6_io_outs_right[42] ,
    \ces_4_6_io_outs_right[41] ,
    \ces_4_6_io_outs_right[40] ,
    \ces_4_6_io_outs_right[39] ,
    \ces_4_6_io_outs_right[38] ,
    \ces_4_6_io_outs_right[37] ,
    \ces_4_6_io_outs_right[36] ,
    \ces_4_6_io_outs_right[35] ,
    \ces_4_6_io_outs_right[34] ,
    \ces_4_6_io_outs_right[33] ,
    \ces_4_6_io_outs_right[32] ,
    \ces_4_6_io_outs_right[31] ,
    \ces_4_6_io_outs_right[30] ,
    \ces_4_6_io_outs_right[29] ,
    \ces_4_6_io_outs_right[28] ,
    \ces_4_6_io_outs_right[27] ,
    \ces_4_6_io_outs_right[26] ,
    \ces_4_6_io_outs_right[25] ,
    \ces_4_6_io_outs_right[24] ,
    \ces_4_6_io_outs_right[23] ,
    \ces_4_6_io_outs_right[22] ,
    \ces_4_6_io_outs_right[21] ,
    \ces_4_6_io_outs_right[20] ,
    \ces_4_6_io_outs_right[19] ,
    \ces_4_6_io_outs_right[18] ,
    \ces_4_6_io_outs_right[17] ,
    \ces_4_6_io_outs_right[16] ,
    \ces_4_6_io_outs_right[15] ,
    \ces_4_6_io_outs_right[14] ,
    \ces_4_6_io_outs_right[13] ,
    \ces_4_6_io_outs_right[12] ,
    \ces_4_6_io_outs_right[11] ,
    \ces_4_6_io_outs_right[10] ,
    \ces_4_6_io_outs_right[9] ,
    \ces_4_6_io_outs_right[8] ,
    \ces_4_6_io_outs_right[7] ,
    \ces_4_6_io_outs_right[6] ,
    \ces_4_6_io_outs_right[5] ,
    \ces_4_6_io_outs_right[4] ,
    \ces_4_6_io_outs_right[3] ,
    \ces_4_6_io_outs_right[2] ,
    \ces_4_6_io_outs_right[1] ,
    \ces_4_6_io_outs_right[0] }),
    .io_outs_up({\ces_4_6_io_outs_up[63] ,
    \ces_4_6_io_outs_up[62] ,
    \ces_4_6_io_outs_up[61] ,
    \ces_4_6_io_outs_up[60] ,
    \ces_4_6_io_outs_up[59] ,
    \ces_4_6_io_outs_up[58] ,
    \ces_4_6_io_outs_up[57] ,
    \ces_4_6_io_outs_up[56] ,
    \ces_4_6_io_outs_up[55] ,
    \ces_4_6_io_outs_up[54] ,
    \ces_4_6_io_outs_up[53] ,
    \ces_4_6_io_outs_up[52] ,
    \ces_4_6_io_outs_up[51] ,
    \ces_4_6_io_outs_up[50] ,
    \ces_4_6_io_outs_up[49] ,
    \ces_4_6_io_outs_up[48] ,
    \ces_4_6_io_outs_up[47] ,
    \ces_4_6_io_outs_up[46] ,
    \ces_4_6_io_outs_up[45] ,
    \ces_4_6_io_outs_up[44] ,
    \ces_4_6_io_outs_up[43] ,
    \ces_4_6_io_outs_up[42] ,
    \ces_4_6_io_outs_up[41] ,
    \ces_4_6_io_outs_up[40] ,
    \ces_4_6_io_outs_up[39] ,
    \ces_4_6_io_outs_up[38] ,
    \ces_4_6_io_outs_up[37] ,
    \ces_4_6_io_outs_up[36] ,
    \ces_4_6_io_outs_up[35] ,
    \ces_4_6_io_outs_up[34] ,
    \ces_4_6_io_outs_up[33] ,
    \ces_4_6_io_outs_up[32] ,
    \ces_4_6_io_outs_up[31] ,
    \ces_4_6_io_outs_up[30] ,
    \ces_4_6_io_outs_up[29] ,
    \ces_4_6_io_outs_up[28] ,
    \ces_4_6_io_outs_up[27] ,
    \ces_4_6_io_outs_up[26] ,
    \ces_4_6_io_outs_up[25] ,
    \ces_4_6_io_outs_up[24] ,
    \ces_4_6_io_outs_up[23] ,
    \ces_4_6_io_outs_up[22] ,
    \ces_4_6_io_outs_up[21] ,
    \ces_4_6_io_outs_up[20] ,
    \ces_4_6_io_outs_up[19] ,
    \ces_4_6_io_outs_up[18] ,
    \ces_4_6_io_outs_up[17] ,
    \ces_4_6_io_outs_up[16] ,
    \ces_4_6_io_outs_up[15] ,
    \ces_4_6_io_outs_up[14] ,
    \ces_4_6_io_outs_up[13] ,
    \ces_4_6_io_outs_up[12] ,
    \ces_4_6_io_outs_up[11] ,
    \ces_4_6_io_outs_up[10] ,
    \ces_4_6_io_outs_up[9] ,
    \ces_4_6_io_outs_up[8] ,
    \ces_4_6_io_outs_up[7] ,
    \ces_4_6_io_outs_up[6] ,
    \ces_4_6_io_outs_up[5] ,
    \ces_4_6_io_outs_up[4] ,
    \ces_4_6_io_outs_up[3] ,
    \ces_4_6_io_outs_up[2] ,
    \ces_4_6_io_outs_up[1] ,
    \ces_4_6_io_outs_up[0] }));
 Element ces_4_7 (.clock(clknet_3_6_0_clock),
    .io_lsbIns_1(ces_4_6_io_lsbOuts_1),
    .io_lsbIns_2(ces_4_6_io_lsbOuts_2),
    .io_lsbIns_3(ces_4_6_io_lsbOuts_3),
    .io_lsbIns_4(ces_4_6_io_lsbOuts_4),
    .io_lsbIns_5(ces_4_6_io_lsbOuts_5),
    .io_lsbIns_6(ces_4_6_io_lsbOuts_6),
    .io_lsbIns_7(ces_4_6_io_lsbOuts_7),
    .io_lsbOuts_0(ces_4_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_4_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_4_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_4_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_4_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_4_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_4_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_4_7_io_lsbOuts_7),
    .io_ins_down({\ces_4_7_io_ins_down[63] ,
    \ces_4_7_io_ins_down[62] ,
    \ces_4_7_io_ins_down[61] ,
    \ces_4_7_io_ins_down[60] ,
    \ces_4_7_io_ins_down[59] ,
    \ces_4_7_io_ins_down[58] ,
    \ces_4_7_io_ins_down[57] ,
    \ces_4_7_io_ins_down[56] ,
    \ces_4_7_io_ins_down[55] ,
    \ces_4_7_io_ins_down[54] ,
    \ces_4_7_io_ins_down[53] ,
    \ces_4_7_io_ins_down[52] ,
    \ces_4_7_io_ins_down[51] ,
    \ces_4_7_io_ins_down[50] ,
    \ces_4_7_io_ins_down[49] ,
    \ces_4_7_io_ins_down[48] ,
    \ces_4_7_io_ins_down[47] ,
    \ces_4_7_io_ins_down[46] ,
    \ces_4_7_io_ins_down[45] ,
    \ces_4_7_io_ins_down[44] ,
    \ces_4_7_io_ins_down[43] ,
    \ces_4_7_io_ins_down[42] ,
    \ces_4_7_io_ins_down[41] ,
    \ces_4_7_io_ins_down[40] ,
    \ces_4_7_io_ins_down[39] ,
    \ces_4_7_io_ins_down[38] ,
    \ces_4_7_io_ins_down[37] ,
    \ces_4_7_io_ins_down[36] ,
    \ces_4_7_io_ins_down[35] ,
    \ces_4_7_io_ins_down[34] ,
    \ces_4_7_io_ins_down[33] ,
    \ces_4_7_io_ins_down[32] ,
    \ces_4_7_io_ins_down[31] ,
    \ces_4_7_io_ins_down[30] ,
    \ces_4_7_io_ins_down[29] ,
    \ces_4_7_io_ins_down[28] ,
    \ces_4_7_io_ins_down[27] ,
    \ces_4_7_io_ins_down[26] ,
    \ces_4_7_io_ins_down[25] ,
    \ces_4_7_io_ins_down[24] ,
    \ces_4_7_io_ins_down[23] ,
    \ces_4_7_io_ins_down[22] ,
    \ces_4_7_io_ins_down[21] ,
    \ces_4_7_io_ins_down[20] ,
    \ces_4_7_io_ins_down[19] ,
    \ces_4_7_io_ins_down[18] ,
    \ces_4_7_io_ins_down[17] ,
    \ces_4_7_io_ins_down[16] ,
    \ces_4_7_io_ins_down[15] ,
    \ces_4_7_io_ins_down[14] ,
    \ces_4_7_io_ins_down[13] ,
    \ces_4_7_io_ins_down[12] ,
    \ces_4_7_io_ins_down[11] ,
    \ces_4_7_io_ins_down[10] ,
    \ces_4_7_io_ins_down[9] ,
    \ces_4_7_io_ins_down[8] ,
    \ces_4_7_io_ins_down[7] ,
    \ces_4_7_io_ins_down[6] ,
    \ces_4_7_io_ins_down[5] ,
    \ces_4_7_io_ins_down[4] ,
    \ces_4_7_io_ins_down[3] ,
    \ces_4_7_io_ins_down[2] ,
    \ces_4_7_io_ins_down[1] ,
    \ces_4_7_io_ins_down[0] }),
    .io_ins_left({net828,
    net827,
    net826,
    net825,
    net823,
    net822,
    net821,
    net820,
    net819,
    net818,
    net817,
    net816,
    net815,
    net814,
    net812,
    net811,
    net810,
    net809,
    net808,
    net807,
    net806,
    net805,
    net804,
    net803,
    net801,
    net800,
    net799,
    net798,
    net797,
    net796,
    net795,
    net794,
    net793,
    net792,
    net790,
    net789,
    net788,
    net787,
    net786,
    net785,
    net784,
    net783,
    net782,
    net781,
    net779,
    net778,
    net777,
    net776,
    net775,
    net774,
    net773,
    net772,
    net771,
    net770,
    net832,
    net831,
    net830,
    net829,
    net824,
    net813,
    net802,
    net791,
    net780,
    net769}),
    .io_ins_right({\ces_4_6_io_outs_right[63] ,
    \ces_4_6_io_outs_right[62] ,
    \ces_4_6_io_outs_right[61] ,
    \ces_4_6_io_outs_right[60] ,
    \ces_4_6_io_outs_right[59] ,
    \ces_4_6_io_outs_right[58] ,
    \ces_4_6_io_outs_right[57] ,
    \ces_4_6_io_outs_right[56] ,
    \ces_4_6_io_outs_right[55] ,
    \ces_4_6_io_outs_right[54] ,
    \ces_4_6_io_outs_right[53] ,
    \ces_4_6_io_outs_right[52] ,
    \ces_4_6_io_outs_right[51] ,
    \ces_4_6_io_outs_right[50] ,
    \ces_4_6_io_outs_right[49] ,
    \ces_4_6_io_outs_right[48] ,
    \ces_4_6_io_outs_right[47] ,
    \ces_4_6_io_outs_right[46] ,
    \ces_4_6_io_outs_right[45] ,
    \ces_4_6_io_outs_right[44] ,
    \ces_4_6_io_outs_right[43] ,
    \ces_4_6_io_outs_right[42] ,
    \ces_4_6_io_outs_right[41] ,
    \ces_4_6_io_outs_right[40] ,
    \ces_4_6_io_outs_right[39] ,
    \ces_4_6_io_outs_right[38] ,
    \ces_4_6_io_outs_right[37] ,
    \ces_4_6_io_outs_right[36] ,
    \ces_4_6_io_outs_right[35] ,
    \ces_4_6_io_outs_right[34] ,
    \ces_4_6_io_outs_right[33] ,
    \ces_4_6_io_outs_right[32] ,
    \ces_4_6_io_outs_right[31] ,
    \ces_4_6_io_outs_right[30] ,
    \ces_4_6_io_outs_right[29] ,
    \ces_4_6_io_outs_right[28] ,
    \ces_4_6_io_outs_right[27] ,
    \ces_4_6_io_outs_right[26] ,
    \ces_4_6_io_outs_right[25] ,
    \ces_4_6_io_outs_right[24] ,
    \ces_4_6_io_outs_right[23] ,
    \ces_4_6_io_outs_right[22] ,
    \ces_4_6_io_outs_right[21] ,
    \ces_4_6_io_outs_right[20] ,
    \ces_4_6_io_outs_right[19] ,
    \ces_4_6_io_outs_right[18] ,
    \ces_4_6_io_outs_right[17] ,
    \ces_4_6_io_outs_right[16] ,
    \ces_4_6_io_outs_right[15] ,
    \ces_4_6_io_outs_right[14] ,
    \ces_4_6_io_outs_right[13] ,
    \ces_4_6_io_outs_right[12] ,
    \ces_4_6_io_outs_right[11] ,
    \ces_4_6_io_outs_right[10] ,
    \ces_4_6_io_outs_right[9] ,
    \ces_4_6_io_outs_right[8] ,
    \ces_4_6_io_outs_right[7] ,
    \ces_4_6_io_outs_right[6] ,
    \ces_4_6_io_outs_right[5] ,
    \ces_4_6_io_outs_right[4] ,
    \ces_4_6_io_outs_right[3] ,
    \ces_4_6_io_outs_right[2] ,
    \ces_4_6_io_outs_right[1] ,
    \ces_4_6_io_outs_right[0] }),
    .io_ins_up({\ces_3_7_io_outs_up[63] ,
    \ces_3_7_io_outs_up[62] ,
    \ces_3_7_io_outs_up[61] ,
    \ces_3_7_io_outs_up[60] ,
    \ces_3_7_io_outs_up[59] ,
    \ces_3_7_io_outs_up[58] ,
    \ces_3_7_io_outs_up[57] ,
    \ces_3_7_io_outs_up[56] ,
    \ces_3_7_io_outs_up[55] ,
    \ces_3_7_io_outs_up[54] ,
    \ces_3_7_io_outs_up[53] ,
    \ces_3_7_io_outs_up[52] ,
    \ces_3_7_io_outs_up[51] ,
    \ces_3_7_io_outs_up[50] ,
    \ces_3_7_io_outs_up[49] ,
    \ces_3_7_io_outs_up[48] ,
    \ces_3_7_io_outs_up[47] ,
    \ces_3_7_io_outs_up[46] ,
    \ces_3_7_io_outs_up[45] ,
    \ces_3_7_io_outs_up[44] ,
    \ces_3_7_io_outs_up[43] ,
    \ces_3_7_io_outs_up[42] ,
    \ces_3_7_io_outs_up[41] ,
    \ces_3_7_io_outs_up[40] ,
    \ces_3_7_io_outs_up[39] ,
    \ces_3_7_io_outs_up[38] ,
    \ces_3_7_io_outs_up[37] ,
    \ces_3_7_io_outs_up[36] ,
    \ces_3_7_io_outs_up[35] ,
    \ces_3_7_io_outs_up[34] ,
    \ces_3_7_io_outs_up[33] ,
    \ces_3_7_io_outs_up[32] ,
    \ces_3_7_io_outs_up[31] ,
    \ces_3_7_io_outs_up[30] ,
    \ces_3_7_io_outs_up[29] ,
    \ces_3_7_io_outs_up[28] ,
    \ces_3_7_io_outs_up[27] ,
    \ces_3_7_io_outs_up[26] ,
    \ces_3_7_io_outs_up[25] ,
    \ces_3_7_io_outs_up[24] ,
    \ces_3_7_io_outs_up[23] ,
    \ces_3_7_io_outs_up[22] ,
    \ces_3_7_io_outs_up[21] ,
    \ces_3_7_io_outs_up[20] ,
    \ces_3_7_io_outs_up[19] ,
    \ces_3_7_io_outs_up[18] ,
    \ces_3_7_io_outs_up[17] ,
    \ces_3_7_io_outs_up[16] ,
    \ces_3_7_io_outs_up[15] ,
    \ces_3_7_io_outs_up[14] ,
    \ces_3_7_io_outs_up[13] ,
    \ces_3_7_io_outs_up[12] ,
    \ces_3_7_io_outs_up[11] ,
    \ces_3_7_io_outs_up[10] ,
    \ces_3_7_io_outs_up[9] ,
    \ces_3_7_io_outs_up[8] ,
    \ces_3_7_io_outs_up[7] ,
    \ces_3_7_io_outs_up[6] ,
    \ces_3_7_io_outs_up[5] ,
    \ces_3_7_io_outs_up[4] ,
    \ces_3_7_io_outs_up[3] ,
    \ces_3_7_io_outs_up[2] ,
    \ces_3_7_io_outs_up[1] ,
    \ces_3_7_io_outs_up[0] }),
    .io_outs_down({\ces_3_7_io_ins_down[63] ,
    \ces_3_7_io_ins_down[62] ,
    \ces_3_7_io_ins_down[61] ,
    \ces_3_7_io_ins_down[60] ,
    \ces_3_7_io_ins_down[59] ,
    \ces_3_7_io_ins_down[58] ,
    \ces_3_7_io_ins_down[57] ,
    \ces_3_7_io_ins_down[56] ,
    \ces_3_7_io_ins_down[55] ,
    \ces_3_7_io_ins_down[54] ,
    \ces_3_7_io_ins_down[53] ,
    \ces_3_7_io_ins_down[52] ,
    \ces_3_7_io_ins_down[51] ,
    \ces_3_7_io_ins_down[50] ,
    \ces_3_7_io_ins_down[49] ,
    \ces_3_7_io_ins_down[48] ,
    \ces_3_7_io_ins_down[47] ,
    \ces_3_7_io_ins_down[46] ,
    \ces_3_7_io_ins_down[45] ,
    \ces_3_7_io_ins_down[44] ,
    \ces_3_7_io_ins_down[43] ,
    \ces_3_7_io_ins_down[42] ,
    \ces_3_7_io_ins_down[41] ,
    \ces_3_7_io_ins_down[40] ,
    \ces_3_7_io_ins_down[39] ,
    \ces_3_7_io_ins_down[38] ,
    \ces_3_7_io_ins_down[37] ,
    \ces_3_7_io_ins_down[36] ,
    \ces_3_7_io_ins_down[35] ,
    \ces_3_7_io_ins_down[34] ,
    \ces_3_7_io_ins_down[33] ,
    \ces_3_7_io_ins_down[32] ,
    \ces_3_7_io_ins_down[31] ,
    \ces_3_7_io_ins_down[30] ,
    \ces_3_7_io_ins_down[29] ,
    \ces_3_7_io_ins_down[28] ,
    \ces_3_7_io_ins_down[27] ,
    \ces_3_7_io_ins_down[26] ,
    \ces_3_7_io_ins_down[25] ,
    \ces_3_7_io_ins_down[24] ,
    \ces_3_7_io_ins_down[23] ,
    \ces_3_7_io_ins_down[22] ,
    \ces_3_7_io_ins_down[21] ,
    \ces_3_7_io_ins_down[20] ,
    \ces_3_7_io_ins_down[19] ,
    \ces_3_7_io_ins_down[18] ,
    \ces_3_7_io_ins_down[17] ,
    \ces_3_7_io_ins_down[16] ,
    \ces_3_7_io_ins_down[15] ,
    \ces_3_7_io_ins_down[14] ,
    \ces_3_7_io_ins_down[13] ,
    \ces_3_7_io_ins_down[12] ,
    \ces_3_7_io_ins_down[11] ,
    \ces_3_7_io_ins_down[10] ,
    \ces_3_7_io_ins_down[9] ,
    \ces_3_7_io_ins_down[8] ,
    \ces_3_7_io_ins_down[7] ,
    \ces_3_7_io_ins_down[6] ,
    \ces_3_7_io_ins_down[5] ,
    \ces_3_7_io_ins_down[4] ,
    \ces_3_7_io_ins_down[3] ,
    \ces_3_7_io_ins_down[2] ,
    \ces_3_7_io_ins_down[1] ,
    \ces_3_7_io_ins_down[0] }),
    .io_outs_left({\ces_4_6_io_ins_left[63] ,
    \ces_4_6_io_ins_left[62] ,
    \ces_4_6_io_ins_left[61] ,
    \ces_4_6_io_ins_left[60] ,
    \ces_4_6_io_ins_left[59] ,
    \ces_4_6_io_ins_left[58] ,
    \ces_4_6_io_ins_left[57] ,
    \ces_4_6_io_ins_left[56] ,
    \ces_4_6_io_ins_left[55] ,
    \ces_4_6_io_ins_left[54] ,
    \ces_4_6_io_ins_left[53] ,
    \ces_4_6_io_ins_left[52] ,
    \ces_4_6_io_ins_left[51] ,
    \ces_4_6_io_ins_left[50] ,
    \ces_4_6_io_ins_left[49] ,
    \ces_4_6_io_ins_left[48] ,
    \ces_4_6_io_ins_left[47] ,
    \ces_4_6_io_ins_left[46] ,
    \ces_4_6_io_ins_left[45] ,
    \ces_4_6_io_ins_left[44] ,
    \ces_4_6_io_ins_left[43] ,
    \ces_4_6_io_ins_left[42] ,
    \ces_4_6_io_ins_left[41] ,
    \ces_4_6_io_ins_left[40] ,
    \ces_4_6_io_ins_left[39] ,
    \ces_4_6_io_ins_left[38] ,
    \ces_4_6_io_ins_left[37] ,
    \ces_4_6_io_ins_left[36] ,
    \ces_4_6_io_ins_left[35] ,
    \ces_4_6_io_ins_left[34] ,
    \ces_4_6_io_ins_left[33] ,
    \ces_4_6_io_ins_left[32] ,
    \ces_4_6_io_ins_left[31] ,
    \ces_4_6_io_ins_left[30] ,
    \ces_4_6_io_ins_left[29] ,
    \ces_4_6_io_ins_left[28] ,
    \ces_4_6_io_ins_left[27] ,
    \ces_4_6_io_ins_left[26] ,
    \ces_4_6_io_ins_left[25] ,
    \ces_4_6_io_ins_left[24] ,
    \ces_4_6_io_ins_left[23] ,
    \ces_4_6_io_ins_left[22] ,
    \ces_4_6_io_ins_left[21] ,
    \ces_4_6_io_ins_left[20] ,
    \ces_4_6_io_ins_left[19] ,
    \ces_4_6_io_ins_left[18] ,
    \ces_4_6_io_ins_left[17] ,
    \ces_4_6_io_ins_left[16] ,
    \ces_4_6_io_ins_left[15] ,
    \ces_4_6_io_ins_left[14] ,
    \ces_4_6_io_ins_left[13] ,
    \ces_4_6_io_ins_left[12] ,
    \ces_4_6_io_ins_left[11] ,
    \ces_4_6_io_ins_left[10] ,
    \ces_4_6_io_ins_left[9] ,
    \ces_4_6_io_ins_left[8] ,
    \ces_4_6_io_ins_left[7] ,
    \ces_4_6_io_ins_left[6] ,
    \ces_4_6_io_ins_left[5] ,
    \ces_4_6_io_ins_left[4] ,
    \ces_4_6_io_ins_left[3] ,
    \ces_4_6_io_ins_left[2] ,
    \ces_4_6_io_ins_left[1] ,
    \ces_4_6_io_ins_left[0] }),
    .io_outs_right({net3452,
    net3451,
    net3450,
    net3449,
    net3447,
    net3446,
    net3445,
    net3444,
    net3443,
    net3442,
    net3441,
    net3440,
    net3439,
    net3438,
    net3436,
    net3435,
    net3434,
    net3433,
    net3432,
    net3431,
    net3430,
    net3429,
    net3428,
    net3427,
    net3425,
    net3424,
    net3423,
    net3422,
    net3421,
    net3420,
    net3419,
    net3418,
    net3417,
    net3416,
    net3414,
    net3413,
    net3412,
    net3411,
    net3410,
    net3409,
    net3408,
    net3407,
    net3406,
    net3405,
    net3403,
    net3402,
    net3401,
    net3400,
    net3399,
    net3398,
    net3397,
    net3396,
    net3395,
    net3394,
    net3456,
    net3455,
    net3454,
    net3453,
    net3448,
    net3437,
    net3426,
    net3415,
    net3404,
    net3393}),
    .io_outs_up({\ces_4_7_io_outs_up[63] ,
    \ces_4_7_io_outs_up[62] ,
    \ces_4_7_io_outs_up[61] ,
    \ces_4_7_io_outs_up[60] ,
    \ces_4_7_io_outs_up[59] ,
    \ces_4_7_io_outs_up[58] ,
    \ces_4_7_io_outs_up[57] ,
    \ces_4_7_io_outs_up[56] ,
    \ces_4_7_io_outs_up[55] ,
    \ces_4_7_io_outs_up[54] ,
    \ces_4_7_io_outs_up[53] ,
    \ces_4_7_io_outs_up[52] ,
    \ces_4_7_io_outs_up[51] ,
    \ces_4_7_io_outs_up[50] ,
    \ces_4_7_io_outs_up[49] ,
    \ces_4_7_io_outs_up[48] ,
    \ces_4_7_io_outs_up[47] ,
    \ces_4_7_io_outs_up[46] ,
    \ces_4_7_io_outs_up[45] ,
    \ces_4_7_io_outs_up[44] ,
    \ces_4_7_io_outs_up[43] ,
    \ces_4_7_io_outs_up[42] ,
    \ces_4_7_io_outs_up[41] ,
    \ces_4_7_io_outs_up[40] ,
    \ces_4_7_io_outs_up[39] ,
    \ces_4_7_io_outs_up[38] ,
    \ces_4_7_io_outs_up[37] ,
    \ces_4_7_io_outs_up[36] ,
    \ces_4_7_io_outs_up[35] ,
    \ces_4_7_io_outs_up[34] ,
    \ces_4_7_io_outs_up[33] ,
    \ces_4_7_io_outs_up[32] ,
    \ces_4_7_io_outs_up[31] ,
    \ces_4_7_io_outs_up[30] ,
    \ces_4_7_io_outs_up[29] ,
    \ces_4_7_io_outs_up[28] ,
    \ces_4_7_io_outs_up[27] ,
    \ces_4_7_io_outs_up[26] ,
    \ces_4_7_io_outs_up[25] ,
    \ces_4_7_io_outs_up[24] ,
    \ces_4_7_io_outs_up[23] ,
    \ces_4_7_io_outs_up[22] ,
    \ces_4_7_io_outs_up[21] ,
    \ces_4_7_io_outs_up[20] ,
    \ces_4_7_io_outs_up[19] ,
    \ces_4_7_io_outs_up[18] ,
    \ces_4_7_io_outs_up[17] ,
    \ces_4_7_io_outs_up[16] ,
    \ces_4_7_io_outs_up[15] ,
    \ces_4_7_io_outs_up[14] ,
    \ces_4_7_io_outs_up[13] ,
    \ces_4_7_io_outs_up[12] ,
    \ces_4_7_io_outs_up[11] ,
    \ces_4_7_io_outs_up[10] ,
    \ces_4_7_io_outs_up[9] ,
    \ces_4_7_io_outs_up[8] ,
    \ces_4_7_io_outs_up[7] ,
    \ces_4_7_io_outs_up[6] ,
    \ces_4_7_io_outs_up[5] ,
    \ces_4_7_io_outs_up[4] ,
    \ces_4_7_io_outs_up[3] ,
    \ces_4_7_io_outs_up[2] ,
    \ces_4_7_io_outs_up[1] ,
    \ces_4_7_io_outs_up[0] }));
 Element ces_5_0 (.clock(clknet_3_4_0_clock),
    .io_lsbIns_1(net4196),
    .io_lsbIns_2(net4197),
    .io_lsbIns_3(net4198),
    .io_lsbIns_4(net4199),
    .io_lsbIns_5(net4200),
    .io_lsbIns_6(net4201),
    .io_lsbIns_7(net4202),
    .io_lsbOuts_0(ces_5_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_0_io_lsbOuts_7),
    .io_ins_down({\ces_5_0_io_ins_down[63] ,
    \ces_5_0_io_ins_down[62] ,
    \ces_5_0_io_ins_down[61] ,
    \ces_5_0_io_ins_down[60] ,
    \ces_5_0_io_ins_down[59] ,
    \ces_5_0_io_ins_down[58] ,
    \ces_5_0_io_ins_down[57] ,
    \ces_5_0_io_ins_down[56] ,
    \ces_5_0_io_ins_down[55] ,
    \ces_5_0_io_ins_down[54] ,
    \ces_5_0_io_ins_down[53] ,
    \ces_5_0_io_ins_down[52] ,
    \ces_5_0_io_ins_down[51] ,
    \ces_5_0_io_ins_down[50] ,
    \ces_5_0_io_ins_down[49] ,
    \ces_5_0_io_ins_down[48] ,
    \ces_5_0_io_ins_down[47] ,
    \ces_5_0_io_ins_down[46] ,
    \ces_5_0_io_ins_down[45] ,
    \ces_5_0_io_ins_down[44] ,
    \ces_5_0_io_ins_down[43] ,
    \ces_5_0_io_ins_down[42] ,
    \ces_5_0_io_ins_down[41] ,
    \ces_5_0_io_ins_down[40] ,
    \ces_5_0_io_ins_down[39] ,
    \ces_5_0_io_ins_down[38] ,
    \ces_5_0_io_ins_down[37] ,
    \ces_5_0_io_ins_down[36] ,
    \ces_5_0_io_ins_down[35] ,
    \ces_5_0_io_ins_down[34] ,
    \ces_5_0_io_ins_down[33] ,
    \ces_5_0_io_ins_down[32] ,
    \ces_5_0_io_ins_down[31] ,
    \ces_5_0_io_ins_down[30] ,
    \ces_5_0_io_ins_down[29] ,
    \ces_5_0_io_ins_down[28] ,
    \ces_5_0_io_ins_down[27] ,
    \ces_5_0_io_ins_down[26] ,
    \ces_5_0_io_ins_down[25] ,
    \ces_5_0_io_ins_down[24] ,
    \ces_5_0_io_ins_down[23] ,
    \ces_5_0_io_ins_down[22] ,
    \ces_5_0_io_ins_down[21] ,
    \ces_5_0_io_ins_down[20] ,
    \ces_5_0_io_ins_down[19] ,
    \ces_5_0_io_ins_down[18] ,
    \ces_5_0_io_ins_down[17] ,
    \ces_5_0_io_ins_down[16] ,
    \ces_5_0_io_ins_down[15] ,
    \ces_5_0_io_ins_down[14] ,
    \ces_5_0_io_ins_down[13] ,
    \ces_5_0_io_ins_down[12] ,
    \ces_5_0_io_ins_down[11] ,
    \ces_5_0_io_ins_down[10] ,
    \ces_5_0_io_ins_down[9] ,
    \ces_5_0_io_ins_down[8] ,
    \ces_5_0_io_ins_down[7] ,
    \ces_5_0_io_ins_down[6] ,
    \ces_5_0_io_ins_down[5] ,
    \ces_5_0_io_ins_down[4] ,
    \ces_5_0_io_ins_down[3] ,
    \ces_5_0_io_ins_down[2] ,
    \ces_5_0_io_ins_down[1] ,
    \ces_5_0_io_ins_down[0] }),
    .io_ins_left({\ces_5_0_io_ins_left[63] ,
    \ces_5_0_io_ins_left[62] ,
    \ces_5_0_io_ins_left[61] ,
    \ces_5_0_io_ins_left[60] ,
    \ces_5_0_io_ins_left[59] ,
    \ces_5_0_io_ins_left[58] ,
    \ces_5_0_io_ins_left[57] ,
    \ces_5_0_io_ins_left[56] ,
    \ces_5_0_io_ins_left[55] ,
    \ces_5_0_io_ins_left[54] ,
    \ces_5_0_io_ins_left[53] ,
    \ces_5_0_io_ins_left[52] ,
    \ces_5_0_io_ins_left[51] ,
    \ces_5_0_io_ins_left[50] ,
    \ces_5_0_io_ins_left[49] ,
    \ces_5_0_io_ins_left[48] ,
    \ces_5_0_io_ins_left[47] ,
    \ces_5_0_io_ins_left[46] ,
    \ces_5_0_io_ins_left[45] ,
    \ces_5_0_io_ins_left[44] ,
    \ces_5_0_io_ins_left[43] ,
    \ces_5_0_io_ins_left[42] ,
    \ces_5_0_io_ins_left[41] ,
    \ces_5_0_io_ins_left[40] ,
    \ces_5_0_io_ins_left[39] ,
    \ces_5_0_io_ins_left[38] ,
    \ces_5_0_io_ins_left[37] ,
    \ces_5_0_io_ins_left[36] ,
    \ces_5_0_io_ins_left[35] ,
    \ces_5_0_io_ins_left[34] ,
    \ces_5_0_io_ins_left[33] ,
    \ces_5_0_io_ins_left[32] ,
    \ces_5_0_io_ins_left[31] ,
    \ces_5_0_io_ins_left[30] ,
    \ces_5_0_io_ins_left[29] ,
    \ces_5_0_io_ins_left[28] ,
    \ces_5_0_io_ins_left[27] ,
    \ces_5_0_io_ins_left[26] ,
    \ces_5_0_io_ins_left[25] ,
    \ces_5_0_io_ins_left[24] ,
    \ces_5_0_io_ins_left[23] ,
    \ces_5_0_io_ins_left[22] ,
    \ces_5_0_io_ins_left[21] ,
    \ces_5_0_io_ins_left[20] ,
    \ces_5_0_io_ins_left[19] ,
    \ces_5_0_io_ins_left[18] ,
    \ces_5_0_io_ins_left[17] ,
    \ces_5_0_io_ins_left[16] ,
    \ces_5_0_io_ins_left[15] ,
    \ces_5_0_io_ins_left[14] ,
    \ces_5_0_io_ins_left[13] ,
    \ces_5_0_io_ins_left[12] ,
    \ces_5_0_io_ins_left[11] ,
    \ces_5_0_io_ins_left[10] ,
    \ces_5_0_io_ins_left[9] ,
    \ces_5_0_io_ins_left[8] ,
    \ces_5_0_io_ins_left[7] ,
    \ces_5_0_io_ins_left[6] ,
    \ces_5_0_io_ins_left[5] ,
    \ces_5_0_io_ins_left[4] ,
    \ces_5_0_io_ins_left[3] ,
    \ces_5_0_io_ins_left[2] ,
    \ces_5_0_io_ins_left[1] ,
    \ces_5_0_io_ins_left[0] }),
    .io_ins_right({net1404,
    net1403,
    net1402,
    net1401,
    net1399,
    net1398,
    net1397,
    net1396,
    net1395,
    net1394,
    net1393,
    net1392,
    net1391,
    net1390,
    net1388,
    net1387,
    net1386,
    net1385,
    net1384,
    net1383,
    net1382,
    net1381,
    net1380,
    net1379,
    net1377,
    net1376,
    net1375,
    net1374,
    net1373,
    net1372,
    net1371,
    net1370,
    net1369,
    net1368,
    net1366,
    net1365,
    net1364,
    net1363,
    net1362,
    net1361,
    net1360,
    net1359,
    net1358,
    net1357,
    net1355,
    net1354,
    net1353,
    net1352,
    net1351,
    net1350,
    net1349,
    net1348,
    net1347,
    net1346,
    net1408,
    net1407,
    net1406,
    net1405,
    net1400,
    net1389,
    net1378,
    net1367,
    net1356,
    net1345}),
    .io_ins_up({\ces_4_0_io_outs_up[63] ,
    \ces_4_0_io_outs_up[62] ,
    \ces_4_0_io_outs_up[61] ,
    \ces_4_0_io_outs_up[60] ,
    \ces_4_0_io_outs_up[59] ,
    \ces_4_0_io_outs_up[58] ,
    \ces_4_0_io_outs_up[57] ,
    \ces_4_0_io_outs_up[56] ,
    \ces_4_0_io_outs_up[55] ,
    \ces_4_0_io_outs_up[54] ,
    \ces_4_0_io_outs_up[53] ,
    \ces_4_0_io_outs_up[52] ,
    \ces_4_0_io_outs_up[51] ,
    \ces_4_0_io_outs_up[50] ,
    \ces_4_0_io_outs_up[49] ,
    \ces_4_0_io_outs_up[48] ,
    \ces_4_0_io_outs_up[47] ,
    \ces_4_0_io_outs_up[46] ,
    \ces_4_0_io_outs_up[45] ,
    \ces_4_0_io_outs_up[44] ,
    \ces_4_0_io_outs_up[43] ,
    \ces_4_0_io_outs_up[42] ,
    \ces_4_0_io_outs_up[41] ,
    \ces_4_0_io_outs_up[40] ,
    \ces_4_0_io_outs_up[39] ,
    \ces_4_0_io_outs_up[38] ,
    \ces_4_0_io_outs_up[37] ,
    \ces_4_0_io_outs_up[36] ,
    \ces_4_0_io_outs_up[35] ,
    \ces_4_0_io_outs_up[34] ,
    \ces_4_0_io_outs_up[33] ,
    \ces_4_0_io_outs_up[32] ,
    \ces_4_0_io_outs_up[31] ,
    \ces_4_0_io_outs_up[30] ,
    \ces_4_0_io_outs_up[29] ,
    \ces_4_0_io_outs_up[28] ,
    \ces_4_0_io_outs_up[27] ,
    \ces_4_0_io_outs_up[26] ,
    \ces_4_0_io_outs_up[25] ,
    \ces_4_0_io_outs_up[24] ,
    \ces_4_0_io_outs_up[23] ,
    \ces_4_0_io_outs_up[22] ,
    \ces_4_0_io_outs_up[21] ,
    \ces_4_0_io_outs_up[20] ,
    \ces_4_0_io_outs_up[19] ,
    \ces_4_0_io_outs_up[18] ,
    \ces_4_0_io_outs_up[17] ,
    \ces_4_0_io_outs_up[16] ,
    \ces_4_0_io_outs_up[15] ,
    \ces_4_0_io_outs_up[14] ,
    \ces_4_0_io_outs_up[13] ,
    \ces_4_0_io_outs_up[12] ,
    \ces_4_0_io_outs_up[11] ,
    \ces_4_0_io_outs_up[10] ,
    \ces_4_0_io_outs_up[9] ,
    \ces_4_0_io_outs_up[8] ,
    \ces_4_0_io_outs_up[7] ,
    \ces_4_0_io_outs_up[6] ,
    \ces_4_0_io_outs_up[5] ,
    \ces_4_0_io_outs_up[4] ,
    \ces_4_0_io_outs_up[3] ,
    \ces_4_0_io_outs_up[2] ,
    \ces_4_0_io_outs_up[1] ,
    \ces_4_0_io_outs_up[0] }),
    .io_outs_down({\ces_4_0_io_ins_down[63] ,
    \ces_4_0_io_ins_down[62] ,
    \ces_4_0_io_ins_down[61] ,
    \ces_4_0_io_ins_down[60] ,
    \ces_4_0_io_ins_down[59] ,
    \ces_4_0_io_ins_down[58] ,
    \ces_4_0_io_ins_down[57] ,
    \ces_4_0_io_ins_down[56] ,
    \ces_4_0_io_ins_down[55] ,
    \ces_4_0_io_ins_down[54] ,
    \ces_4_0_io_ins_down[53] ,
    \ces_4_0_io_ins_down[52] ,
    \ces_4_0_io_ins_down[51] ,
    \ces_4_0_io_ins_down[50] ,
    \ces_4_0_io_ins_down[49] ,
    \ces_4_0_io_ins_down[48] ,
    \ces_4_0_io_ins_down[47] ,
    \ces_4_0_io_ins_down[46] ,
    \ces_4_0_io_ins_down[45] ,
    \ces_4_0_io_ins_down[44] ,
    \ces_4_0_io_ins_down[43] ,
    \ces_4_0_io_ins_down[42] ,
    \ces_4_0_io_ins_down[41] ,
    \ces_4_0_io_ins_down[40] ,
    \ces_4_0_io_ins_down[39] ,
    \ces_4_0_io_ins_down[38] ,
    \ces_4_0_io_ins_down[37] ,
    \ces_4_0_io_ins_down[36] ,
    \ces_4_0_io_ins_down[35] ,
    \ces_4_0_io_ins_down[34] ,
    \ces_4_0_io_ins_down[33] ,
    \ces_4_0_io_ins_down[32] ,
    \ces_4_0_io_ins_down[31] ,
    \ces_4_0_io_ins_down[30] ,
    \ces_4_0_io_ins_down[29] ,
    \ces_4_0_io_ins_down[28] ,
    \ces_4_0_io_ins_down[27] ,
    \ces_4_0_io_ins_down[26] ,
    \ces_4_0_io_ins_down[25] ,
    \ces_4_0_io_ins_down[24] ,
    \ces_4_0_io_ins_down[23] ,
    \ces_4_0_io_ins_down[22] ,
    \ces_4_0_io_ins_down[21] ,
    \ces_4_0_io_ins_down[20] ,
    \ces_4_0_io_ins_down[19] ,
    \ces_4_0_io_ins_down[18] ,
    \ces_4_0_io_ins_down[17] ,
    \ces_4_0_io_ins_down[16] ,
    \ces_4_0_io_ins_down[15] ,
    \ces_4_0_io_ins_down[14] ,
    \ces_4_0_io_ins_down[13] ,
    \ces_4_0_io_ins_down[12] ,
    \ces_4_0_io_ins_down[11] ,
    \ces_4_0_io_ins_down[10] ,
    \ces_4_0_io_ins_down[9] ,
    \ces_4_0_io_ins_down[8] ,
    \ces_4_0_io_ins_down[7] ,
    \ces_4_0_io_ins_down[6] ,
    \ces_4_0_io_ins_down[5] ,
    \ces_4_0_io_ins_down[4] ,
    \ces_4_0_io_ins_down[3] ,
    \ces_4_0_io_ins_down[2] ,
    \ces_4_0_io_ins_down[1] ,
    \ces_4_0_io_ins_down[0] }),
    .io_outs_left({net3004,
    net3003,
    net3002,
    net3001,
    net2999,
    net2998,
    net2997,
    net2996,
    net2995,
    net2994,
    net2993,
    net2992,
    net2991,
    net2990,
    net2988,
    net2987,
    net2986,
    net2985,
    net2984,
    net2983,
    net2982,
    net2981,
    net2980,
    net2979,
    net2977,
    net2976,
    net2975,
    net2974,
    net2973,
    net2972,
    net2971,
    net2970,
    net2969,
    net2968,
    net2966,
    net2965,
    net2964,
    net2963,
    net2962,
    net2961,
    net2960,
    net2959,
    net2958,
    net2957,
    net2955,
    net2954,
    net2953,
    net2952,
    net2951,
    net2950,
    net2949,
    net2948,
    net2947,
    net2946,
    net3008,
    net3007,
    net3006,
    net3005,
    net3000,
    net2989,
    net2978,
    net2967,
    net2956,
    net2945}),
    .io_outs_right({\ces_5_0_io_outs_right[63] ,
    \ces_5_0_io_outs_right[62] ,
    \ces_5_0_io_outs_right[61] ,
    \ces_5_0_io_outs_right[60] ,
    \ces_5_0_io_outs_right[59] ,
    \ces_5_0_io_outs_right[58] ,
    \ces_5_0_io_outs_right[57] ,
    \ces_5_0_io_outs_right[56] ,
    \ces_5_0_io_outs_right[55] ,
    \ces_5_0_io_outs_right[54] ,
    \ces_5_0_io_outs_right[53] ,
    \ces_5_0_io_outs_right[52] ,
    \ces_5_0_io_outs_right[51] ,
    \ces_5_0_io_outs_right[50] ,
    \ces_5_0_io_outs_right[49] ,
    \ces_5_0_io_outs_right[48] ,
    \ces_5_0_io_outs_right[47] ,
    \ces_5_0_io_outs_right[46] ,
    \ces_5_0_io_outs_right[45] ,
    \ces_5_0_io_outs_right[44] ,
    \ces_5_0_io_outs_right[43] ,
    \ces_5_0_io_outs_right[42] ,
    \ces_5_0_io_outs_right[41] ,
    \ces_5_0_io_outs_right[40] ,
    \ces_5_0_io_outs_right[39] ,
    \ces_5_0_io_outs_right[38] ,
    \ces_5_0_io_outs_right[37] ,
    \ces_5_0_io_outs_right[36] ,
    \ces_5_0_io_outs_right[35] ,
    \ces_5_0_io_outs_right[34] ,
    \ces_5_0_io_outs_right[33] ,
    \ces_5_0_io_outs_right[32] ,
    \ces_5_0_io_outs_right[31] ,
    \ces_5_0_io_outs_right[30] ,
    \ces_5_0_io_outs_right[29] ,
    \ces_5_0_io_outs_right[28] ,
    \ces_5_0_io_outs_right[27] ,
    \ces_5_0_io_outs_right[26] ,
    \ces_5_0_io_outs_right[25] ,
    \ces_5_0_io_outs_right[24] ,
    \ces_5_0_io_outs_right[23] ,
    \ces_5_0_io_outs_right[22] ,
    \ces_5_0_io_outs_right[21] ,
    \ces_5_0_io_outs_right[20] ,
    \ces_5_0_io_outs_right[19] ,
    \ces_5_0_io_outs_right[18] ,
    \ces_5_0_io_outs_right[17] ,
    \ces_5_0_io_outs_right[16] ,
    \ces_5_0_io_outs_right[15] ,
    \ces_5_0_io_outs_right[14] ,
    \ces_5_0_io_outs_right[13] ,
    \ces_5_0_io_outs_right[12] ,
    \ces_5_0_io_outs_right[11] ,
    \ces_5_0_io_outs_right[10] ,
    \ces_5_0_io_outs_right[9] ,
    \ces_5_0_io_outs_right[8] ,
    \ces_5_0_io_outs_right[7] ,
    \ces_5_0_io_outs_right[6] ,
    \ces_5_0_io_outs_right[5] ,
    \ces_5_0_io_outs_right[4] ,
    \ces_5_0_io_outs_right[3] ,
    \ces_5_0_io_outs_right[2] ,
    \ces_5_0_io_outs_right[1] ,
    \ces_5_0_io_outs_right[0] }),
    .io_outs_up({\ces_5_0_io_outs_up[63] ,
    \ces_5_0_io_outs_up[62] ,
    \ces_5_0_io_outs_up[61] ,
    \ces_5_0_io_outs_up[60] ,
    \ces_5_0_io_outs_up[59] ,
    \ces_5_0_io_outs_up[58] ,
    \ces_5_0_io_outs_up[57] ,
    \ces_5_0_io_outs_up[56] ,
    \ces_5_0_io_outs_up[55] ,
    \ces_5_0_io_outs_up[54] ,
    \ces_5_0_io_outs_up[53] ,
    \ces_5_0_io_outs_up[52] ,
    \ces_5_0_io_outs_up[51] ,
    \ces_5_0_io_outs_up[50] ,
    \ces_5_0_io_outs_up[49] ,
    \ces_5_0_io_outs_up[48] ,
    \ces_5_0_io_outs_up[47] ,
    \ces_5_0_io_outs_up[46] ,
    \ces_5_0_io_outs_up[45] ,
    \ces_5_0_io_outs_up[44] ,
    \ces_5_0_io_outs_up[43] ,
    \ces_5_0_io_outs_up[42] ,
    \ces_5_0_io_outs_up[41] ,
    \ces_5_0_io_outs_up[40] ,
    \ces_5_0_io_outs_up[39] ,
    \ces_5_0_io_outs_up[38] ,
    \ces_5_0_io_outs_up[37] ,
    \ces_5_0_io_outs_up[36] ,
    \ces_5_0_io_outs_up[35] ,
    \ces_5_0_io_outs_up[34] ,
    \ces_5_0_io_outs_up[33] ,
    \ces_5_0_io_outs_up[32] ,
    \ces_5_0_io_outs_up[31] ,
    \ces_5_0_io_outs_up[30] ,
    \ces_5_0_io_outs_up[29] ,
    \ces_5_0_io_outs_up[28] ,
    \ces_5_0_io_outs_up[27] ,
    \ces_5_0_io_outs_up[26] ,
    \ces_5_0_io_outs_up[25] ,
    \ces_5_0_io_outs_up[24] ,
    \ces_5_0_io_outs_up[23] ,
    \ces_5_0_io_outs_up[22] ,
    \ces_5_0_io_outs_up[21] ,
    \ces_5_0_io_outs_up[20] ,
    \ces_5_0_io_outs_up[19] ,
    \ces_5_0_io_outs_up[18] ,
    \ces_5_0_io_outs_up[17] ,
    \ces_5_0_io_outs_up[16] ,
    \ces_5_0_io_outs_up[15] ,
    \ces_5_0_io_outs_up[14] ,
    \ces_5_0_io_outs_up[13] ,
    \ces_5_0_io_outs_up[12] ,
    \ces_5_0_io_outs_up[11] ,
    \ces_5_0_io_outs_up[10] ,
    \ces_5_0_io_outs_up[9] ,
    \ces_5_0_io_outs_up[8] ,
    \ces_5_0_io_outs_up[7] ,
    \ces_5_0_io_outs_up[6] ,
    \ces_5_0_io_outs_up[5] ,
    \ces_5_0_io_outs_up[4] ,
    \ces_5_0_io_outs_up[3] ,
    \ces_5_0_io_outs_up[2] ,
    \ces_5_0_io_outs_up[1] ,
    \ces_5_0_io_outs_up[0] }));
 Element ces_5_1 (.clock(clknet_3_4_0_clock),
    .io_lsbIns_1(ces_5_0_io_lsbOuts_1),
    .io_lsbIns_2(ces_5_0_io_lsbOuts_2),
    .io_lsbIns_3(ces_5_0_io_lsbOuts_3),
    .io_lsbIns_4(ces_5_0_io_lsbOuts_4),
    .io_lsbIns_5(ces_5_0_io_lsbOuts_5),
    .io_lsbIns_6(ces_5_0_io_lsbOuts_6),
    .io_lsbIns_7(ces_5_0_io_lsbOuts_7),
    .io_lsbOuts_0(ces_5_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_1_io_lsbOuts_7),
    .io_ins_down({\ces_5_1_io_ins_down[63] ,
    \ces_5_1_io_ins_down[62] ,
    \ces_5_1_io_ins_down[61] ,
    \ces_5_1_io_ins_down[60] ,
    \ces_5_1_io_ins_down[59] ,
    \ces_5_1_io_ins_down[58] ,
    \ces_5_1_io_ins_down[57] ,
    \ces_5_1_io_ins_down[56] ,
    \ces_5_1_io_ins_down[55] ,
    \ces_5_1_io_ins_down[54] ,
    \ces_5_1_io_ins_down[53] ,
    \ces_5_1_io_ins_down[52] ,
    \ces_5_1_io_ins_down[51] ,
    \ces_5_1_io_ins_down[50] ,
    \ces_5_1_io_ins_down[49] ,
    \ces_5_1_io_ins_down[48] ,
    \ces_5_1_io_ins_down[47] ,
    \ces_5_1_io_ins_down[46] ,
    \ces_5_1_io_ins_down[45] ,
    \ces_5_1_io_ins_down[44] ,
    \ces_5_1_io_ins_down[43] ,
    \ces_5_1_io_ins_down[42] ,
    \ces_5_1_io_ins_down[41] ,
    \ces_5_1_io_ins_down[40] ,
    \ces_5_1_io_ins_down[39] ,
    \ces_5_1_io_ins_down[38] ,
    \ces_5_1_io_ins_down[37] ,
    \ces_5_1_io_ins_down[36] ,
    \ces_5_1_io_ins_down[35] ,
    \ces_5_1_io_ins_down[34] ,
    \ces_5_1_io_ins_down[33] ,
    \ces_5_1_io_ins_down[32] ,
    \ces_5_1_io_ins_down[31] ,
    \ces_5_1_io_ins_down[30] ,
    \ces_5_1_io_ins_down[29] ,
    \ces_5_1_io_ins_down[28] ,
    \ces_5_1_io_ins_down[27] ,
    \ces_5_1_io_ins_down[26] ,
    \ces_5_1_io_ins_down[25] ,
    \ces_5_1_io_ins_down[24] ,
    \ces_5_1_io_ins_down[23] ,
    \ces_5_1_io_ins_down[22] ,
    \ces_5_1_io_ins_down[21] ,
    \ces_5_1_io_ins_down[20] ,
    \ces_5_1_io_ins_down[19] ,
    \ces_5_1_io_ins_down[18] ,
    \ces_5_1_io_ins_down[17] ,
    \ces_5_1_io_ins_down[16] ,
    \ces_5_1_io_ins_down[15] ,
    \ces_5_1_io_ins_down[14] ,
    \ces_5_1_io_ins_down[13] ,
    \ces_5_1_io_ins_down[12] ,
    \ces_5_1_io_ins_down[11] ,
    \ces_5_1_io_ins_down[10] ,
    \ces_5_1_io_ins_down[9] ,
    \ces_5_1_io_ins_down[8] ,
    \ces_5_1_io_ins_down[7] ,
    \ces_5_1_io_ins_down[6] ,
    \ces_5_1_io_ins_down[5] ,
    \ces_5_1_io_ins_down[4] ,
    \ces_5_1_io_ins_down[3] ,
    \ces_5_1_io_ins_down[2] ,
    \ces_5_1_io_ins_down[1] ,
    \ces_5_1_io_ins_down[0] }),
    .io_ins_left({\ces_5_1_io_ins_left[63] ,
    \ces_5_1_io_ins_left[62] ,
    \ces_5_1_io_ins_left[61] ,
    \ces_5_1_io_ins_left[60] ,
    \ces_5_1_io_ins_left[59] ,
    \ces_5_1_io_ins_left[58] ,
    \ces_5_1_io_ins_left[57] ,
    \ces_5_1_io_ins_left[56] ,
    \ces_5_1_io_ins_left[55] ,
    \ces_5_1_io_ins_left[54] ,
    \ces_5_1_io_ins_left[53] ,
    \ces_5_1_io_ins_left[52] ,
    \ces_5_1_io_ins_left[51] ,
    \ces_5_1_io_ins_left[50] ,
    \ces_5_1_io_ins_left[49] ,
    \ces_5_1_io_ins_left[48] ,
    \ces_5_1_io_ins_left[47] ,
    \ces_5_1_io_ins_left[46] ,
    \ces_5_1_io_ins_left[45] ,
    \ces_5_1_io_ins_left[44] ,
    \ces_5_1_io_ins_left[43] ,
    \ces_5_1_io_ins_left[42] ,
    \ces_5_1_io_ins_left[41] ,
    \ces_5_1_io_ins_left[40] ,
    \ces_5_1_io_ins_left[39] ,
    \ces_5_1_io_ins_left[38] ,
    \ces_5_1_io_ins_left[37] ,
    \ces_5_1_io_ins_left[36] ,
    \ces_5_1_io_ins_left[35] ,
    \ces_5_1_io_ins_left[34] ,
    \ces_5_1_io_ins_left[33] ,
    \ces_5_1_io_ins_left[32] ,
    \ces_5_1_io_ins_left[31] ,
    \ces_5_1_io_ins_left[30] ,
    \ces_5_1_io_ins_left[29] ,
    \ces_5_1_io_ins_left[28] ,
    \ces_5_1_io_ins_left[27] ,
    \ces_5_1_io_ins_left[26] ,
    \ces_5_1_io_ins_left[25] ,
    \ces_5_1_io_ins_left[24] ,
    \ces_5_1_io_ins_left[23] ,
    \ces_5_1_io_ins_left[22] ,
    \ces_5_1_io_ins_left[21] ,
    \ces_5_1_io_ins_left[20] ,
    \ces_5_1_io_ins_left[19] ,
    \ces_5_1_io_ins_left[18] ,
    \ces_5_1_io_ins_left[17] ,
    \ces_5_1_io_ins_left[16] ,
    \ces_5_1_io_ins_left[15] ,
    \ces_5_1_io_ins_left[14] ,
    \ces_5_1_io_ins_left[13] ,
    \ces_5_1_io_ins_left[12] ,
    \ces_5_1_io_ins_left[11] ,
    \ces_5_1_io_ins_left[10] ,
    \ces_5_1_io_ins_left[9] ,
    \ces_5_1_io_ins_left[8] ,
    \ces_5_1_io_ins_left[7] ,
    \ces_5_1_io_ins_left[6] ,
    \ces_5_1_io_ins_left[5] ,
    \ces_5_1_io_ins_left[4] ,
    \ces_5_1_io_ins_left[3] ,
    \ces_5_1_io_ins_left[2] ,
    \ces_5_1_io_ins_left[1] ,
    \ces_5_1_io_ins_left[0] }),
    .io_ins_right({\ces_5_0_io_outs_right[63] ,
    \ces_5_0_io_outs_right[62] ,
    \ces_5_0_io_outs_right[61] ,
    \ces_5_0_io_outs_right[60] ,
    \ces_5_0_io_outs_right[59] ,
    \ces_5_0_io_outs_right[58] ,
    \ces_5_0_io_outs_right[57] ,
    \ces_5_0_io_outs_right[56] ,
    \ces_5_0_io_outs_right[55] ,
    \ces_5_0_io_outs_right[54] ,
    \ces_5_0_io_outs_right[53] ,
    \ces_5_0_io_outs_right[52] ,
    \ces_5_0_io_outs_right[51] ,
    \ces_5_0_io_outs_right[50] ,
    \ces_5_0_io_outs_right[49] ,
    \ces_5_0_io_outs_right[48] ,
    \ces_5_0_io_outs_right[47] ,
    \ces_5_0_io_outs_right[46] ,
    \ces_5_0_io_outs_right[45] ,
    \ces_5_0_io_outs_right[44] ,
    \ces_5_0_io_outs_right[43] ,
    \ces_5_0_io_outs_right[42] ,
    \ces_5_0_io_outs_right[41] ,
    \ces_5_0_io_outs_right[40] ,
    \ces_5_0_io_outs_right[39] ,
    \ces_5_0_io_outs_right[38] ,
    \ces_5_0_io_outs_right[37] ,
    \ces_5_0_io_outs_right[36] ,
    \ces_5_0_io_outs_right[35] ,
    \ces_5_0_io_outs_right[34] ,
    \ces_5_0_io_outs_right[33] ,
    \ces_5_0_io_outs_right[32] ,
    \ces_5_0_io_outs_right[31] ,
    \ces_5_0_io_outs_right[30] ,
    \ces_5_0_io_outs_right[29] ,
    \ces_5_0_io_outs_right[28] ,
    \ces_5_0_io_outs_right[27] ,
    \ces_5_0_io_outs_right[26] ,
    \ces_5_0_io_outs_right[25] ,
    \ces_5_0_io_outs_right[24] ,
    \ces_5_0_io_outs_right[23] ,
    \ces_5_0_io_outs_right[22] ,
    \ces_5_0_io_outs_right[21] ,
    \ces_5_0_io_outs_right[20] ,
    \ces_5_0_io_outs_right[19] ,
    \ces_5_0_io_outs_right[18] ,
    \ces_5_0_io_outs_right[17] ,
    \ces_5_0_io_outs_right[16] ,
    \ces_5_0_io_outs_right[15] ,
    \ces_5_0_io_outs_right[14] ,
    \ces_5_0_io_outs_right[13] ,
    \ces_5_0_io_outs_right[12] ,
    \ces_5_0_io_outs_right[11] ,
    \ces_5_0_io_outs_right[10] ,
    \ces_5_0_io_outs_right[9] ,
    \ces_5_0_io_outs_right[8] ,
    \ces_5_0_io_outs_right[7] ,
    \ces_5_0_io_outs_right[6] ,
    \ces_5_0_io_outs_right[5] ,
    \ces_5_0_io_outs_right[4] ,
    \ces_5_0_io_outs_right[3] ,
    \ces_5_0_io_outs_right[2] ,
    \ces_5_0_io_outs_right[1] ,
    \ces_5_0_io_outs_right[0] }),
    .io_ins_up({\ces_4_1_io_outs_up[63] ,
    \ces_4_1_io_outs_up[62] ,
    \ces_4_1_io_outs_up[61] ,
    \ces_4_1_io_outs_up[60] ,
    \ces_4_1_io_outs_up[59] ,
    \ces_4_1_io_outs_up[58] ,
    \ces_4_1_io_outs_up[57] ,
    \ces_4_1_io_outs_up[56] ,
    \ces_4_1_io_outs_up[55] ,
    \ces_4_1_io_outs_up[54] ,
    \ces_4_1_io_outs_up[53] ,
    \ces_4_1_io_outs_up[52] ,
    \ces_4_1_io_outs_up[51] ,
    \ces_4_1_io_outs_up[50] ,
    \ces_4_1_io_outs_up[49] ,
    \ces_4_1_io_outs_up[48] ,
    \ces_4_1_io_outs_up[47] ,
    \ces_4_1_io_outs_up[46] ,
    \ces_4_1_io_outs_up[45] ,
    \ces_4_1_io_outs_up[44] ,
    \ces_4_1_io_outs_up[43] ,
    \ces_4_1_io_outs_up[42] ,
    \ces_4_1_io_outs_up[41] ,
    \ces_4_1_io_outs_up[40] ,
    \ces_4_1_io_outs_up[39] ,
    \ces_4_1_io_outs_up[38] ,
    \ces_4_1_io_outs_up[37] ,
    \ces_4_1_io_outs_up[36] ,
    \ces_4_1_io_outs_up[35] ,
    \ces_4_1_io_outs_up[34] ,
    \ces_4_1_io_outs_up[33] ,
    \ces_4_1_io_outs_up[32] ,
    \ces_4_1_io_outs_up[31] ,
    \ces_4_1_io_outs_up[30] ,
    \ces_4_1_io_outs_up[29] ,
    \ces_4_1_io_outs_up[28] ,
    \ces_4_1_io_outs_up[27] ,
    \ces_4_1_io_outs_up[26] ,
    \ces_4_1_io_outs_up[25] ,
    \ces_4_1_io_outs_up[24] ,
    \ces_4_1_io_outs_up[23] ,
    \ces_4_1_io_outs_up[22] ,
    \ces_4_1_io_outs_up[21] ,
    \ces_4_1_io_outs_up[20] ,
    \ces_4_1_io_outs_up[19] ,
    \ces_4_1_io_outs_up[18] ,
    \ces_4_1_io_outs_up[17] ,
    \ces_4_1_io_outs_up[16] ,
    \ces_4_1_io_outs_up[15] ,
    \ces_4_1_io_outs_up[14] ,
    \ces_4_1_io_outs_up[13] ,
    \ces_4_1_io_outs_up[12] ,
    \ces_4_1_io_outs_up[11] ,
    \ces_4_1_io_outs_up[10] ,
    \ces_4_1_io_outs_up[9] ,
    \ces_4_1_io_outs_up[8] ,
    \ces_4_1_io_outs_up[7] ,
    \ces_4_1_io_outs_up[6] ,
    \ces_4_1_io_outs_up[5] ,
    \ces_4_1_io_outs_up[4] ,
    \ces_4_1_io_outs_up[3] ,
    \ces_4_1_io_outs_up[2] ,
    \ces_4_1_io_outs_up[1] ,
    \ces_4_1_io_outs_up[0] }),
    .io_outs_down({\ces_4_1_io_ins_down[63] ,
    \ces_4_1_io_ins_down[62] ,
    \ces_4_1_io_ins_down[61] ,
    \ces_4_1_io_ins_down[60] ,
    \ces_4_1_io_ins_down[59] ,
    \ces_4_1_io_ins_down[58] ,
    \ces_4_1_io_ins_down[57] ,
    \ces_4_1_io_ins_down[56] ,
    \ces_4_1_io_ins_down[55] ,
    \ces_4_1_io_ins_down[54] ,
    \ces_4_1_io_ins_down[53] ,
    \ces_4_1_io_ins_down[52] ,
    \ces_4_1_io_ins_down[51] ,
    \ces_4_1_io_ins_down[50] ,
    \ces_4_1_io_ins_down[49] ,
    \ces_4_1_io_ins_down[48] ,
    \ces_4_1_io_ins_down[47] ,
    \ces_4_1_io_ins_down[46] ,
    \ces_4_1_io_ins_down[45] ,
    \ces_4_1_io_ins_down[44] ,
    \ces_4_1_io_ins_down[43] ,
    \ces_4_1_io_ins_down[42] ,
    \ces_4_1_io_ins_down[41] ,
    \ces_4_1_io_ins_down[40] ,
    \ces_4_1_io_ins_down[39] ,
    \ces_4_1_io_ins_down[38] ,
    \ces_4_1_io_ins_down[37] ,
    \ces_4_1_io_ins_down[36] ,
    \ces_4_1_io_ins_down[35] ,
    \ces_4_1_io_ins_down[34] ,
    \ces_4_1_io_ins_down[33] ,
    \ces_4_1_io_ins_down[32] ,
    \ces_4_1_io_ins_down[31] ,
    \ces_4_1_io_ins_down[30] ,
    \ces_4_1_io_ins_down[29] ,
    \ces_4_1_io_ins_down[28] ,
    \ces_4_1_io_ins_down[27] ,
    \ces_4_1_io_ins_down[26] ,
    \ces_4_1_io_ins_down[25] ,
    \ces_4_1_io_ins_down[24] ,
    \ces_4_1_io_ins_down[23] ,
    \ces_4_1_io_ins_down[22] ,
    \ces_4_1_io_ins_down[21] ,
    \ces_4_1_io_ins_down[20] ,
    \ces_4_1_io_ins_down[19] ,
    \ces_4_1_io_ins_down[18] ,
    \ces_4_1_io_ins_down[17] ,
    \ces_4_1_io_ins_down[16] ,
    \ces_4_1_io_ins_down[15] ,
    \ces_4_1_io_ins_down[14] ,
    \ces_4_1_io_ins_down[13] ,
    \ces_4_1_io_ins_down[12] ,
    \ces_4_1_io_ins_down[11] ,
    \ces_4_1_io_ins_down[10] ,
    \ces_4_1_io_ins_down[9] ,
    \ces_4_1_io_ins_down[8] ,
    \ces_4_1_io_ins_down[7] ,
    \ces_4_1_io_ins_down[6] ,
    \ces_4_1_io_ins_down[5] ,
    \ces_4_1_io_ins_down[4] ,
    \ces_4_1_io_ins_down[3] ,
    \ces_4_1_io_ins_down[2] ,
    \ces_4_1_io_ins_down[1] ,
    \ces_4_1_io_ins_down[0] }),
    .io_outs_left({\ces_5_0_io_ins_left[63] ,
    \ces_5_0_io_ins_left[62] ,
    \ces_5_0_io_ins_left[61] ,
    \ces_5_0_io_ins_left[60] ,
    \ces_5_0_io_ins_left[59] ,
    \ces_5_0_io_ins_left[58] ,
    \ces_5_0_io_ins_left[57] ,
    \ces_5_0_io_ins_left[56] ,
    \ces_5_0_io_ins_left[55] ,
    \ces_5_0_io_ins_left[54] ,
    \ces_5_0_io_ins_left[53] ,
    \ces_5_0_io_ins_left[52] ,
    \ces_5_0_io_ins_left[51] ,
    \ces_5_0_io_ins_left[50] ,
    \ces_5_0_io_ins_left[49] ,
    \ces_5_0_io_ins_left[48] ,
    \ces_5_0_io_ins_left[47] ,
    \ces_5_0_io_ins_left[46] ,
    \ces_5_0_io_ins_left[45] ,
    \ces_5_0_io_ins_left[44] ,
    \ces_5_0_io_ins_left[43] ,
    \ces_5_0_io_ins_left[42] ,
    \ces_5_0_io_ins_left[41] ,
    \ces_5_0_io_ins_left[40] ,
    \ces_5_0_io_ins_left[39] ,
    \ces_5_0_io_ins_left[38] ,
    \ces_5_0_io_ins_left[37] ,
    \ces_5_0_io_ins_left[36] ,
    \ces_5_0_io_ins_left[35] ,
    \ces_5_0_io_ins_left[34] ,
    \ces_5_0_io_ins_left[33] ,
    \ces_5_0_io_ins_left[32] ,
    \ces_5_0_io_ins_left[31] ,
    \ces_5_0_io_ins_left[30] ,
    \ces_5_0_io_ins_left[29] ,
    \ces_5_0_io_ins_left[28] ,
    \ces_5_0_io_ins_left[27] ,
    \ces_5_0_io_ins_left[26] ,
    \ces_5_0_io_ins_left[25] ,
    \ces_5_0_io_ins_left[24] ,
    \ces_5_0_io_ins_left[23] ,
    \ces_5_0_io_ins_left[22] ,
    \ces_5_0_io_ins_left[21] ,
    \ces_5_0_io_ins_left[20] ,
    \ces_5_0_io_ins_left[19] ,
    \ces_5_0_io_ins_left[18] ,
    \ces_5_0_io_ins_left[17] ,
    \ces_5_0_io_ins_left[16] ,
    \ces_5_0_io_ins_left[15] ,
    \ces_5_0_io_ins_left[14] ,
    \ces_5_0_io_ins_left[13] ,
    \ces_5_0_io_ins_left[12] ,
    \ces_5_0_io_ins_left[11] ,
    \ces_5_0_io_ins_left[10] ,
    \ces_5_0_io_ins_left[9] ,
    \ces_5_0_io_ins_left[8] ,
    \ces_5_0_io_ins_left[7] ,
    \ces_5_0_io_ins_left[6] ,
    \ces_5_0_io_ins_left[5] ,
    \ces_5_0_io_ins_left[4] ,
    \ces_5_0_io_ins_left[3] ,
    \ces_5_0_io_ins_left[2] ,
    \ces_5_0_io_ins_left[1] ,
    \ces_5_0_io_ins_left[0] }),
    .io_outs_right({\ces_5_1_io_outs_right[63] ,
    \ces_5_1_io_outs_right[62] ,
    \ces_5_1_io_outs_right[61] ,
    \ces_5_1_io_outs_right[60] ,
    \ces_5_1_io_outs_right[59] ,
    \ces_5_1_io_outs_right[58] ,
    \ces_5_1_io_outs_right[57] ,
    \ces_5_1_io_outs_right[56] ,
    \ces_5_1_io_outs_right[55] ,
    \ces_5_1_io_outs_right[54] ,
    \ces_5_1_io_outs_right[53] ,
    \ces_5_1_io_outs_right[52] ,
    \ces_5_1_io_outs_right[51] ,
    \ces_5_1_io_outs_right[50] ,
    \ces_5_1_io_outs_right[49] ,
    \ces_5_1_io_outs_right[48] ,
    \ces_5_1_io_outs_right[47] ,
    \ces_5_1_io_outs_right[46] ,
    \ces_5_1_io_outs_right[45] ,
    \ces_5_1_io_outs_right[44] ,
    \ces_5_1_io_outs_right[43] ,
    \ces_5_1_io_outs_right[42] ,
    \ces_5_1_io_outs_right[41] ,
    \ces_5_1_io_outs_right[40] ,
    \ces_5_1_io_outs_right[39] ,
    \ces_5_1_io_outs_right[38] ,
    \ces_5_1_io_outs_right[37] ,
    \ces_5_1_io_outs_right[36] ,
    \ces_5_1_io_outs_right[35] ,
    \ces_5_1_io_outs_right[34] ,
    \ces_5_1_io_outs_right[33] ,
    \ces_5_1_io_outs_right[32] ,
    \ces_5_1_io_outs_right[31] ,
    \ces_5_1_io_outs_right[30] ,
    \ces_5_1_io_outs_right[29] ,
    \ces_5_1_io_outs_right[28] ,
    \ces_5_1_io_outs_right[27] ,
    \ces_5_1_io_outs_right[26] ,
    \ces_5_1_io_outs_right[25] ,
    \ces_5_1_io_outs_right[24] ,
    \ces_5_1_io_outs_right[23] ,
    \ces_5_1_io_outs_right[22] ,
    \ces_5_1_io_outs_right[21] ,
    \ces_5_1_io_outs_right[20] ,
    \ces_5_1_io_outs_right[19] ,
    \ces_5_1_io_outs_right[18] ,
    \ces_5_1_io_outs_right[17] ,
    \ces_5_1_io_outs_right[16] ,
    \ces_5_1_io_outs_right[15] ,
    \ces_5_1_io_outs_right[14] ,
    \ces_5_1_io_outs_right[13] ,
    \ces_5_1_io_outs_right[12] ,
    \ces_5_1_io_outs_right[11] ,
    \ces_5_1_io_outs_right[10] ,
    \ces_5_1_io_outs_right[9] ,
    \ces_5_1_io_outs_right[8] ,
    \ces_5_1_io_outs_right[7] ,
    \ces_5_1_io_outs_right[6] ,
    \ces_5_1_io_outs_right[5] ,
    \ces_5_1_io_outs_right[4] ,
    \ces_5_1_io_outs_right[3] ,
    \ces_5_1_io_outs_right[2] ,
    \ces_5_1_io_outs_right[1] ,
    \ces_5_1_io_outs_right[0] }),
    .io_outs_up({\ces_5_1_io_outs_up[63] ,
    \ces_5_1_io_outs_up[62] ,
    \ces_5_1_io_outs_up[61] ,
    \ces_5_1_io_outs_up[60] ,
    \ces_5_1_io_outs_up[59] ,
    \ces_5_1_io_outs_up[58] ,
    \ces_5_1_io_outs_up[57] ,
    \ces_5_1_io_outs_up[56] ,
    \ces_5_1_io_outs_up[55] ,
    \ces_5_1_io_outs_up[54] ,
    \ces_5_1_io_outs_up[53] ,
    \ces_5_1_io_outs_up[52] ,
    \ces_5_1_io_outs_up[51] ,
    \ces_5_1_io_outs_up[50] ,
    \ces_5_1_io_outs_up[49] ,
    \ces_5_1_io_outs_up[48] ,
    \ces_5_1_io_outs_up[47] ,
    \ces_5_1_io_outs_up[46] ,
    \ces_5_1_io_outs_up[45] ,
    \ces_5_1_io_outs_up[44] ,
    \ces_5_1_io_outs_up[43] ,
    \ces_5_1_io_outs_up[42] ,
    \ces_5_1_io_outs_up[41] ,
    \ces_5_1_io_outs_up[40] ,
    \ces_5_1_io_outs_up[39] ,
    \ces_5_1_io_outs_up[38] ,
    \ces_5_1_io_outs_up[37] ,
    \ces_5_1_io_outs_up[36] ,
    \ces_5_1_io_outs_up[35] ,
    \ces_5_1_io_outs_up[34] ,
    \ces_5_1_io_outs_up[33] ,
    \ces_5_1_io_outs_up[32] ,
    \ces_5_1_io_outs_up[31] ,
    \ces_5_1_io_outs_up[30] ,
    \ces_5_1_io_outs_up[29] ,
    \ces_5_1_io_outs_up[28] ,
    \ces_5_1_io_outs_up[27] ,
    \ces_5_1_io_outs_up[26] ,
    \ces_5_1_io_outs_up[25] ,
    \ces_5_1_io_outs_up[24] ,
    \ces_5_1_io_outs_up[23] ,
    \ces_5_1_io_outs_up[22] ,
    \ces_5_1_io_outs_up[21] ,
    \ces_5_1_io_outs_up[20] ,
    \ces_5_1_io_outs_up[19] ,
    \ces_5_1_io_outs_up[18] ,
    \ces_5_1_io_outs_up[17] ,
    \ces_5_1_io_outs_up[16] ,
    \ces_5_1_io_outs_up[15] ,
    \ces_5_1_io_outs_up[14] ,
    \ces_5_1_io_outs_up[13] ,
    \ces_5_1_io_outs_up[12] ,
    \ces_5_1_io_outs_up[11] ,
    \ces_5_1_io_outs_up[10] ,
    \ces_5_1_io_outs_up[9] ,
    \ces_5_1_io_outs_up[8] ,
    \ces_5_1_io_outs_up[7] ,
    \ces_5_1_io_outs_up[6] ,
    \ces_5_1_io_outs_up[5] ,
    \ces_5_1_io_outs_up[4] ,
    \ces_5_1_io_outs_up[3] ,
    \ces_5_1_io_outs_up[2] ,
    \ces_5_1_io_outs_up[1] ,
    \ces_5_1_io_outs_up[0] }));
 Element ces_5_2 (.clock(clknet_3_4_0_clock),
    .io_lsbIns_1(ces_5_1_io_lsbOuts_1),
    .io_lsbIns_2(ces_5_1_io_lsbOuts_2),
    .io_lsbIns_3(ces_5_1_io_lsbOuts_3),
    .io_lsbIns_4(ces_5_1_io_lsbOuts_4),
    .io_lsbIns_5(ces_5_1_io_lsbOuts_5),
    .io_lsbIns_6(ces_5_1_io_lsbOuts_6),
    .io_lsbIns_7(ces_5_1_io_lsbOuts_7),
    .io_lsbOuts_0(ces_5_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_2_io_lsbOuts_7),
    .io_ins_down({\ces_5_2_io_ins_down[63] ,
    \ces_5_2_io_ins_down[62] ,
    \ces_5_2_io_ins_down[61] ,
    \ces_5_2_io_ins_down[60] ,
    \ces_5_2_io_ins_down[59] ,
    \ces_5_2_io_ins_down[58] ,
    \ces_5_2_io_ins_down[57] ,
    \ces_5_2_io_ins_down[56] ,
    \ces_5_2_io_ins_down[55] ,
    \ces_5_2_io_ins_down[54] ,
    \ces_5_2_io_ins_down[53] ,
    \ces_5_2_io_ins_down[52] ,
    \ces_5_2_io_ins_down[51] ,
    \ces_5_2_io_ins_down[50] ,
    \ces_5_2_io_ins_down[49] ,
    \ces_5_2_io_ins_down[48] ,
    \ces_5_2_io_ins_down[47] ,
    \ces_5_2_io_ins_down[46] ,
    \ces_5_2_io_ins_down[45] ,
    \ces_5_2_io_ins_down[44] ,
    \ces_5_2_io_ins_down[43] ,
    \ces_5_2_io_ins_down[42] ,
    \ces_5_2_io_ins_down[41] ,
    \ces_5_2_io_ins_down[40] ,
    \ces_5_2_io_ins_down[39] ,
    \ces_5_2_io_ins_down[38] ,
    \ces_5_2_io_ins_down[37] ,
    \ces_5_2_io_ins_down[36] ,
    \ces_5_2_io_ins_down[35] ,
    \ces_5_2_io_ins_down[34] ,
    \ces_5_2_io_ins_down[33] ,
    \ces_5_2_io_ins_down[32] ,
    \ces_5_2_io_ins_down[31] ,
    \ces_5_2_io_ins_down[30] ,
    \ces_5_2_io_ins_down[29] ,
    \ces_5_2_io_ins_down[28] ,
    \ces_5_2_io_ins_down[27] ,
    \ces_5_2_io_ins_down[26] ,
    \ces_5_2_io_ins_down[25] ,
    \ces_5_2_io_ins_down[24] ,
    \ces_5_2_io_ins_down[23] ,
    \ces_5_2_io_ins_down[22] ,
    \ces_5_2_io_ins_down[21] ,
    \ces_5_2_io_ins_down[20] ,
    \ces_5_2_io_ins_down[19] ,
    \ces_5_2_io_ins_down[18] ,
    \ces_5_2_io_ins_down[17] ,
    \ces_5_2_io_ins_down[16] ,
    \ces_5_2_io_ins_down[15] ,
    \ces_5_2_io_ins_down[14] ,
    \ces_5_2_io_ins_down[13] ,
    \ces_5_2_io_ins_down[12] ,
    \ces_5_2_io_ins_down[11] ,
    \ces_5_2_io_ins_down[10] ,
    \ces_5_2_io_ins_down[9] ,
    \ces_5_2_io_ins_down[8] ,
    \ces_5_2_io_ins_down[7] ,
    \ces_5_2_io_ins_down[6] ,
    \ces_5_2_io_ins_down[5] ,
    \ces_5_2_io_ins_down[4] ,
    \ces_5_2_io_ins_down[3] ,
    \ces_5_2_io_ins_down[2] ,
    \ces_5_2_io_ins_down[1] ,
    \ces_5_2_io_ins_down[0] }),
    .io_ins_left({\ces_5_2_io_ins_left[63] ,
    \ces_5_2_io_ins_left[62] ,
    \ces_5_2_io_ins_left[61] ,
    \ces_5_2_io_ins_left[60] ,
    \ces_5_2_io_ins_left[59] ,
    \ces_5_2_io_ins_left[58] ,
    \ces_5_2_io_ins_left[57] ,
    \ces_5_2_io_ins_left[56] ,
    \ces_5_2_io_ins_left[55] ,
    \ces_5_2_io_ins_left[54] ,
    \ces_5_2_io_ins_left[53] ,
    \ces_5_2_io_ins_left[52] ,
    \ces_5_2_io_ins_left[51] ,
    \ces_5_2_io_ins_left[50] ,
    \ces_5_2_io_ins_left[49] ,
    \ces_5_2_io_ins_left[48] ,
    \ces_5_2_io_ins_left[47] ,
    \ces_5_2_io_ins_left[46] ,
    \ces_5_2_io_ins_left[45] ,
    \ces_5_2_io_ins_left[44] ,
    \ces_5_2_io_ins_left[43] ,
    \ces_5_2_io_ins_left[42] ,
    \ces_5_2_io_ins_left[41] ,
    \ces_5_2_io_ins_left[40] ,
    \ces_5_2_io_ins_left[39] ,
    \ces_5_2_io_ins_left[38] ,
    \ces_5_2_io_ins_left[37] ,
    \ces_5_2_io_ins_left[36] ,
    \ces_5_2_io_ins_left[35] ,
    \ces_5_2_io_ins_left[34] ,
    \ces_5_2_io_ins_left[33] ,
    \ces_5_2_io_ins_left[32] ,
    \ces_5_2_io_ins_left[31] ,
    \ces_5_2_io_ins_left[30] ,
    \ces_5_2_io_ins_left[29] ,
    \ces_5_2_io_ins_left[28] ,
    \ces_5_2_io_ins_left[27] ,
    \ces_5_2_io_ins_left[26] ,
    \ces_5_2_io_ins_left[25] ,
    \ces_5_2_io_ins_left[24] ,
    \ces_5_2_io_ins_left[23] ,
    \ces_5_2_io_ins_left[22] ,
    \ces_5_2_io_ins_left[21] ,
    \ces_5_2_io_ins_left[20] ,
    \ces_5_2_io_ins_left[19] ,
    \ces_5_2_io_ins_left[18] ,
    \ces_5_2_io_ins_left[17] ,
    \ces_5_2_io_ins_left[16] ,
    \ces_5_2_io_ins_left[15] ,
    \ces_5_2_io_ins_left[14] ,
    \ces_5_2_io_ins_left[13] ,
    \ces_5_2_io_ins_left[12] ,
    \ces_5_2_io_ins_left[11] ,
    \ces_5_2_io_ins_left[10] ,
    \ces_5_2_io_ins_left[9] ,
    \ces_5_2_io_ins_left[8] ,
    \ces_5_2_io_ins_left[7] ,
    \ces_5_2_io_ins_left[6] ,
    \ces_5_2_io_ins_left[5] ,
    \ces_5_2_io_ins_left[4] ,
    \ces_5_2_io_ins_left[3] ,
    \ces_5_2_io_ins_left[2] ,
    \ces_5_2_io_ins_left[1] ,
    \ces_5_2_io_ins_left[0] }),
    .io_ins_right({\ces_5_1_io_outs_right[63] ,
    \ces_5_1_io_outs_right[62] ,
    \ces_5_1_io_outs_right[61] ,
    \ces_5_1_io_outs_right[60] ,
    \ces_5_1_io_outs_right[59] ,
    \ces_5_1_io_outs_right[58] ,
    \ces_5_1_io_outs_right[57] ,
    \ces_5_1_io_outs_right[56] ,
    \ces_5_1_io_outs_right[55] ,
    \ces_5_1_io_outs_right[54] ,
    \ces_5_1_io_outs_right[53] ,
    \ces_5_1_io_outs_right[52] ,
    \ces_5_1_io_outs_right[51] ,
    \ces_5_1_io_outs_right[50] ,
    \ces_5_1_io_outs_right[49] ,
    \ces_5_1_io_outs_right[48] ,
    \ces_5_1_io_outs_right[47] ,
    \ces_5_1_io_outs_right[46] ,
    \ces_5_1_io_outs_right[45] ,
    \ces_5_1_io_outs_right[44] ,
    \ces_5_1_io_outs_right[43] ,
    \ces_5_1_io_outs_right[42] ,
    \ces_5_1_io_outs_right[41] ,
    \ces_5_1_io_outs_right[40] ,
    \ces_5_1_io_outs_right[39] ,
    \ces_5_1_io_outs_right[38] ,
    \ces_5_1_io_outs_right[37] ,
    \ces_5_1_io_outs_right[36] ,
    \ces_5_1_io_outs_right[35] ,
    \ces_5_1_io_outs_right[34] ,
    \ces_5_1_io_outs_right[33] ,
    \ces_5_1_io_outs_right[32] ,
    \ces_5_1_io_outs_right[31] ,
    \ces_5_1_io_outs_right[30] ,
    \ces_5_1_io_outs_right[29] ,
    \ces_5_1_io_outs_right[28] ,
    \ces_5_1_io_outs_right[27] ,
    \ces_5_1_io_outs_right[26] ,
    \ces_5_1_io_outs_right[25] ,
    \ces_5_1_io_outs_right[24] ,
    \ces_5_1_io_outs_right[23] ,
    \ces_5_1_io_outs_right[22] ,
    \ces_5_1_io_outs_right[21] ,
    \ces_5_1_io_outs_right[20] ,
    \ces_5_1_io_outs_right[19] ,
    \ces_5_1_io_outs_right[18] ,
    \ces_5_1_io_outs_right[17] ,
    \ces_5_1_io_outs_right[16] ,
    \ces_5_1_io_outs_right[15] ,
    \ces_5_1_io_outs_right[14] ,
    \ces_5_1_io_outs_right[13] ,
    \ces_5_1_io_outs_right[12] ,
    \ces_5_1_io_outs_right[11] ,
    \ces_5_1_io_outs_right[10] ,
    \ces_5_1_io_outs_right[9] ,
    \ces_5_1_io_outs_right[8] ,
    \ces_5_1_io_outs_right[7] ,
    \ces_5_1_io_outs_right[6] ,
    \ces_5_1_io_outs_right[5] ,
    \ces_5_1_io_outs_right[4] ,
    \ces_5_1_io_outs_right[3] ,
    \ces_5_1_io_outs_right[2] ,
    \ces_5_1_io_outs_right[1] ,
    \ces_5_1_io_outs_right[0] }),
    .io_ins_up({\ces_4_2_io_outs_up[63] ,
    \ces_4_2_io_outs_up[62] ,
    \ces_4_2_io_outs_up[61] ,
    \ces_4_2_io_outs_up[60] ,
    \ces_4_2_io_outs_up[59] ,
    \ces_4_2_io_outs_up[58] ,
    \ces_4_2_io_outs_up[57] ,
    \ces_4_2_io_outs_up[56] ,
    \ces_4_2_io_outs_up[55] ,
    \ces_4_2_io_outs_up[54] ,
    \ces_4_2_io_outs_up[53] ,
    \ces_4_2_io_outs_up[52] ,
    \ces_4_2_io_outs_up[51] ,
    \ces_4_2_io_outs_up[50] ,
    \ces_4_2_io_outs_up[49] ,
    \ces_4_2_io_outs_up[48] ,
    \ces_4_2_io_outs_up[47] ,
    \ces_4_2_io_outs_up[46] ,
    \ces_4_2_io_outs_up[45] ,
    \ces_4_2_io_outs_up[44] ,
    \ces_4_2_io_outs_up[43] ,
    \ces_4_2_io_outs_up[42] ,
    \ces_4_2_io_outs_up[41] ,
    \ces_4_2_io_outs_up[40] ,
    \ces_4_2_io_outs_up[39] ,
    \ces_4_2_io_outs_up[38] ,
    \ces_4_2_io_outs_up[37] ,
    \ces_4_2_io_outs_up[36] ,
    \ces_4_2_io_outs_up[35] ,
    \ces_4_2_io_outs_up[34] ,
    \ces_4_2_io_outs_up[33] ,
    \ces_4_2_io_outs_up[32] ,
    \ces_4_2_io_outs_up[31] ,
    \ces_4_2_io_outs_up[30] ,
    \ces_4_2_io_outs_up[29] ,
    \ces_4_2_io_outs_up[28] ,
    \ces_4_2_io_outs_up[27] ,
    \ces_4_2_io_outs_up[26] ,
    \ces_4_2_io_outs_up[25] ,
    \ces_4_2_io_outs_up[24] ,
    \ces_4_2_io_outs_up[23] ,
    \ces_4_2_io_outs_up[22] ,
    \ces_4_2_io_outs_up[21] ,
    \ces_4_2_io_outs_up[20] ,
    \ces_4_2_io_outs_up[19] ,
    \ces_4_2_io_outs_up[18] ,
    \ces_4_2_io_outs_up[17] ,
    \ces_4_2_io_outs_up[16] ,
    \ces_4_2_io_outs_up[15] ,
    \ces_4_2_io_outs_up[14] ,
    \ces_4_2_io_outs_up[13] ,
    \ces_4_2_io_outs_up[12] ,
    \ces_4_2_io_outs_up[11] ,
    \ces_4_2_io_outs_up[10] ,
    \ces_4_2_io_outs_up[9] ,
    \ces_4_2_io_outs_up[8] ,
    \ces_4_2_io_outs_up[7] ,
    \ces_4_2_io_outs_up[6] ,
    \ces_4_2_io_outs_up[5] ,
    \ces_4_2_io_outs_up[4] ,
    \ces_4_2_io_outs_up[3] ,
    \ces_4_2_io_outs_up[2] ,
    \ces_4_2_io_outs_up[1] ,
    \ces_4_2_io_outs_up[0] }),
    .io_outs_down({\ces_4_2_io_ins_down[63] ,
    \ces_4_2_io_ins_down[62] ,
    \ces_4_2_io_ins_down[61] ,
    \ces_4_2_io_ins_down[60] ,
    \ces_4_2_io_ins_down[59] ,
    \ces_4_2_io_ins_down[58] ,
    \ces_4_2_io_ins_down[57] ,
    \ces_4_2_io_ins_down[56] ,
    \ces_4_2_io_ins_down[55] ,
    \ces_4_2_io_ins_down[54] ,
    \ces_4_2_io_ins_down[53] ,
    \ces_4_2_io_ins_down[52] ,
    \ces_4_2_io_ins_down[51] ,
    \ces_4_2_io_ins_down[50] ,
    \ces_4_2_io_ins_down[49] ,
    \ces_4_2_io_ins_down[48] ,
    \ces_4_2_io_ins_down[47] ,
    \ces_4_2_io_ins_down[46] ,
    \ces_4_2_io_ins_down[45] ,
    \ces_4_2_io_ins_down[44] ,
    \ces_4_2_io_ins_down[43] ,
    \ces_4_2_io_ins_down[42] ,
    \ces_4_2_io_ins_down[41] ,
    \ces_4_2_io_ins_down[40] ,
    \ces_4_2_io_ins_down[39] ,
    \ces_4_2_io_ins_down[38] ,
    \ces_4_2_io_ins_down[37] ,
    \ces_4_2_io_ins_down[36] ,
    \ces_4_2_io_ins_down[35] ,
    \ces_4_2_io_ins_down[34] ,
    \ces_4_2_io_ins_down[33] ,
    \ces_4_2_io_ins_down[32] ,
    \ces_4_2_io_ins_down[31] ,
    \ces_4_2_io_ins_down[30] ,
    \ces_4_2_io_ins_down[29] ,
    \ces_4_2_io_ins_down[28] ,
    \ces_4_2_io_ins_down[27] ,
    \ces_4_2_io_ins_down[26] ,
    \ces_4_2_io_ins_down[25] ,
    \ces_4_2_io_ins_down[24] ,
    \ces_4_2_io_ins_down[23] ,
    \ces_4_2_io_ins_down[22] ,
    \ces_4_2_io_ins_down[21] ,
    \ces_4_2_io_ins_down[20] ,
    \ces_4_2_io_ins_down[19] ,
    \ces_4_2_io_ins_down[18] ,
    \ces_4_2_io_ins_down[17] ,
    \ces_4_2_io_ins_down[16] ,
    \ces_4_2_io_ins_down[15] ,
    \ces_4_2_io_ins_down[14] ,
    \ces_4_2_io_ins_down[13] ,
    \ces_4_2_io_ins_down[12] ,
    \ces_4_2_io_ins_down[11] ,
    \ces_4_2_io_ins_down[10] ,
    \ces_4_2_io_ins_down[9] ,
    \ces_4_2_io_ins_down[8] ,
    \ces_4_2_io_ins_down[7] ,
    \ces_4_2_io_ins_down[6] ,
    \ces_4_2_io_ins_down[5] ,
    \ces_4_2_io_ins_down[4] ,
    \ces_4_2_io_ins_down[3] ,
    \ces_4_2_io_ins_down[2] ,
    \ces_4_2_io_ins_down[1] ,
    \ces_4_2_io_ins_down[0] }),
    .io_outs_left({\ces_5_1_io_ins_left[63] ,
    \ces_5_1_io_ins_left[62] ,
    \ces_5_1_io_ins_left[61] ,
    \ces_5_1_io_ins_left[60] ,
    \ces_5_1_io_ins_left[59] ,
    \ces_5_1_io_ins_left[58] ,
    \ces_5_1_io_ins_left[57] ,
    \ces_5_1_io_ins_left[56] ,
    \ces_5_1_io_ins_left[55] ,
    \ces_5_1_io_ins_left[54] ,
    \ces_5_1_io_ins_left[53] ,
    \ces_5_1_io_ins_left[52] ,
    \ces_5_1_io_ins_left[51] ,
    \ces_5_1_io_ins_left[50] ,
    \ces_5_1_io_ins_left[49] ,
    \ces_5_1_io_ins_left[48] ,
    \ces_5_1_io_ins_left[47] ,
    \ces_5_1_io_ins_left[46] ,
    \ces_5_1_io_ins_left[45] ,
    \ces_5_1_io_ins_left[44] ,
    \ces_5_1_io_ins_left[43] ,
    \ces_5_1_io_ins_left[42] ,
    \ces_5_1_io_ins_left[41] ,
    \ces_5_1_io_ins_left[40] ,
    \ces_5_1_io_ins_left[39] ,
    \ces_5_1_io_ins_left[38] ,
    \ces_5_1_io_ins_left[37] ,
    \ces_5_1_io_ins_left[36] ,
    \ces_5_1_io_ins_left[35] ,
    \ces_5_1_io_ins_left[34] ,
    \ces_5_1_io_ins_left[33] ,
    \ces_5_1_io_ins_left[32] ,
    \ces_5_1_io_ins_left[31] ,
    \ces_5_1_io_ins_left[30] ,
    \ces_5_1_io_ins_left[29] ,
    \ces_5_1_io_ins_left[28] ,
    \ces_5_1_io_ins_left[27] ,
    \ces_5_1_io_ins_left[26] ,
    \ces_5_1_io_ins_left[25] ,
    \ces_5_1_io_ins_left[24] ,
    \ces_5_1_io_ins_left[23] ,
    \ces_5_1_io_ins_left[22] ,
    \ces_5_1_io_ins_left[21] ,
    \ces_5_1_io_ins_left[20] ,
    \ces_5_1_io_ins_left[19] ,
    \ces_5_1_io_ins_left[18] ,
    \ces_5_1_io_ins_left[17] ,
    \ces_5_1_io_ins_left[16] ,
    \ces_5_1_io_ins_left[15] ,
    \ces_5_1_io_ins_left[14] ,
    \ces_5_1_io_ins_left[13] ,
    \ces_5_1_io_ins_left[12] ,
    \ces_5_1_io_ins_left[11] ,
    \ces_5_1_io_ins_left[10] ,
    \ces_5_1_io_ins_left[9] ,
    \ces_5_1_io_ins_left[8] ,
    \ces_5_1_io_ins_left[7] ,
    \ces_5_1_io_ins_left[6] ,
    \ces_5_1_io_ins_left[5] ,
    \ces_5_1_io_ins_left[4] ,
    \ces_5_1_io_ins_left[3] ,
    \ces_5_1_io_ins_left[2] ,
    \ces_5_1_io_ins_left[1] ,
    \ces_5_1_io_ins_left[0] }),
    .io_outs_right({\ces_5_2_io_outs_right[63] ,
    \ces_5_2_io_outs_right[62] ,
    \ces_5_2_io_outs_right[61] ,
    \ces_5_2_io_outs_right[60] ,
    \ces_5_2_io_outs_right[59] ,
    \ces_5_2_io_outs_right[58] ,
    \ces_5_2_io_outs_right[57] ,
    \ces_5_2_io_outs_right[56] ,
    \ces_5_2_io_outs_right[55] ,
    \ces_5_2_io_outs_right[54] ,
    \ces_5_2_io_outs_right[53] ,
    \ces_5_2_io_outs_right[52] ,
    \ces_5_2_io_outs_right[51] ,
    \ces_5_2_io_outs_right[50] ,
    \ces_5_2_io_outs_right[49] ,
    \ces_5_2_io_outs_right[48] ,
    \ces_5_2_io_outs_right[47] ,
    \ces_5_2_io_outs_right[46] ,
    \ces_5_2_io_outs_right[45] ,
    \ces_5_2_io_outs_right[44] ,
    \ces_5_2_io_outs_right[43] ,
    \ces_5_2_io_outs_right[42] ,
    \ces_5_2_io_outs_right[41] ,
    \ces_5_2_io_outs_right[40] ,
    \ces_5_2_io_outs_right[39] ,
    \ces_5_2_io_outs_right[38] ,
    \ces_5_2_io_outs_right[37] ,
    \ces_5_2_io_outs_right[36] ,
    \ces_5_2_io_outs_right[35] ,
    \ces_5_2_io_outs_right[34] ,
    \ces_5_2_io_outs_right[33] ,
    \ces_5_2_io_outs_right[32] ,
    \ces_5_2_io_outs_right[31] ,
    \ces_5_2_io_outs_right[30] ,
    \ces_5_2_io_outs_right[29] ,
    \ces_5_2_io_outs_right[28] ,
    \ces_5_2_io_outs_right[27] ,
    \ces_5_2_io_outs_right[26] ,
    \ces_5_2_io_outs_right[25] ,
    \ces_5_2_io_outs_right[24] ,
    \ces_5_2_io_outs_right[23] ,
    \ces_5_2_io_outs_right[22] ,
    \ces_5_2_io_outs_right[21] ,
    \ces_5_2_io_outs_right[20] ,
    \ces_5_2_io_outs_right[19] ,
    \ces_5_2_io_outs_right[18] ,
    \ces_5_2_io_outs_right[17] ,
    \ces_5_2_io_outs_right[16] ,
    \ces_5_2_io_outs_right[15] ,
    \ces_5_2_io_outs_right[14] ,
    \ces_5_2_io_outs_right[13] ,
    \ces_5_2_io_outs_right[12] ,
    \ces_5_2_io_outs_right[11] ,
    \ces_5_2_io_outs_right[10] ,
    \ces_5_2_io_outs_right[9] ,
    \ces_5_2_io_outs_right[8] ,
    \ces_5_2_io_outs_right[7] ,
    \ces_5_2_io_outs_right[6] ,
    \ces_5_2_io_outs_right[5] ,
    \ces_5_2_io_outs_right[4] ,
    \ces_5_2_io_outs_right[3] ,
    \ces_5_2_io_outs_right[2] ,
    \ces_5_2_io_outs_right[1] ,
    \ces_5_2_io_outs_right[0] }),
    .io_outs_up({\ces_5_2_io_outs_up[63] ,
    \ces_5_2_io_outs_up[62] ,
    \ces_5_2_io_outs_up[61] ,
    \ces_5_2_io_outs_up[60] ,
    \ces_5_2_io_outs_up[59] ,
    \ces_5_2_io_outs_up[58] ,
    \ces_5_2_io_outs_up[57] ,
    \ces_5_2_io_outs_up[56] ,
    \ces_5_2_io_outs_up[55] ,
    \ces_5_2_io_outs_up[54] ,
    \ces_5_2_io_outs_up[53] ,
    \ces_5_2_io_outs_up[52] ,
    \ces_5_2_io_outs_up[51] ,
    \ces_5_2_io_outs_up[50] ,
    \ces_5_2_io_outs_up[49] ,
    \ces_5_2_io_outs_up[48] ,
    \ces_5_2_io_outs_up[47] ,
    \ces_5_2_io_outs_up[46] ,
    \ces_5_2_io_outs_up[45] ,
    \ces_5_2_io_outs_up[44] ,
    \ces_5_2_io_outs_up[43] ,
    \ces_5_2_io_outs_up[42] ,
    \ces_5_2_io_outs_up[41] ,
    \ces_5_2_io_outs_up[40] ,
    \ces_5_2_io_outs_up[39] ,
    \ces_5_2_io_outs_up[38] ,
    \ces_5_2_io_outs_up[37] ,
    \ces_5_2_io_outs_up[36] ,
    \ces_5_2_io_outs_up[35] ,
    \ces_5_2_io_outs_up[34] ,
    \ces_5_2_io_outs_up[33] ,
    \ces_5_2_io_outs_up[32] ,
    \ces_5_2_io_outs_up[31] ,
    \ces_5_2_io_outs_up[30] ,
    \ces_5_2_io_outs_up[29] ,
    \ces_5_2_io_outs_up[28] ,
    \ces_5_2_io_outs_up[27] ,
    \ces_5_2_io_outs_up[26] ,
    \ces_5_2_io_outs_up[25] ,
    \ces_5_2_io_outs_up[24] ,
    \ces_5_2_io_outs_up[23] ,
    \ces_5_2_io_outs_up[22] ,
    \ces_5_2_io_outs_up[21] ,
    \ces_5_2_io_outs_up[20] ,
    \ces_5_2_io_outs_up[19] ,
    \ces_5_2_io_outs_up[18] ,
    \ces_5_2_io_outs_up[17] ,
    \ces_5_2_io_outs_up[16] ,
    \ces_5_2_io_outs_up[15] ,
    \ces_5_2_io_outs_up[14] ,
    \ces_5_2_io_outs_up[13] ,
    \ces_5_2_io_outs_up[12] ,
    \ces_5_2_io_outs_up[11] ,
    \ces_5_2_io_outs_up[10] ,
    \ces_5_2_io_outs_up[9] ,
    \ces_5_2_io_outs_up[8] ,
    \ces_5_2_io_outs_up[7] ,
    \ces_5_2_io_outs_up[6] ,
    \ces_5_2_io_outs_up[5] ,
    \ces_5_2_io_outs_up[4] ,
    \ces_5_2_io_outs_up[3] ,
    \ces_5_2_io_outs_up[2] ,
    \ces_5_2_io_outs_up[1] ,
    \ces_5_2_io_outs_up[0] }));
 Element ces_5_3 (.clock(clknet_3_4_0_clock),
    .io_lsbIns_1(ces_5_2_io_lsbOuts_1),
    .io_lsbIns_2(ces_5_2_io_lsbOuts_2),
    .io_lsbIns_3(ces_5_2_io_lsbOuts_3),
    .io_lsbIns_4(ces_5_2_io_lsbOuts_4),
    .io_lsbIns_5(ces_5_2_io_lsbOuts_5),
    .io_lsbIns_6(ces_5_2_io_lsbOuts_6),
    .io_lsbIns_7(ces_5_2_io_lsbOuts_7),
    .io_lsbOuts_0(ces_5_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_3_io_lsbOuts_7),
    .io_ins_down({\ces_5_3_io_ins_down[63] ,
    \ces_5_3_io_ins_down[62] ,
    \ces_5_3_io_ins_down[61] ,
    \ces_5_3_io_ins_down[60] ,
    \ces_5_3_io_ins_down[59] ,
    \ces_5_3_io_ins_down[58] ,
    \ces_5_3_io_ins_down[57] ,
    \ces_5_3_io_ins_down[56] ,
    \ces_5_3_io_ins_down[55] ,
    \ces_5_3_io_ins_down[54] ,
    \ces_5_3_io_ins_down[53] ,
    \ces_5_3_io_ins_down[52] ,
    \ces_5_3_io_ins_down[51] ,
    \ces_5_3_io_ins_down[50] ,
    \ces_5_3_io_ins_down[49] ,
    \ces_5_3_io_ins_down[48] ,
    \ces_5_3_io_ins_down[47] ,
    \ces_5_3_io_ins_down[46] ,
    \ces_5_3_io_ins_down[45] ,
    \ces_5_3_io_ins_down[44] ,
    \ces_5_3_io_ins_down[43] ,
    \ces_5_3_io_ins_down[42] ,
    \ces_5_3_io_ins_down[41] ,
    \ces_5_3_io_ins_down[40] ,
    \ces_5_3_io_ins_down[39] ,
    \ces_5_3_io_ins_down[38] ,
    \ces_5_3_io_ins_down[37] ,
    \ces_5_3_io_ins_down[36] ,
    \ces_5_3_io_ins_down[35] ,
    \ces_5_3_io_ins_down[34] ,
    \ces_5_3_io_ins_down[33] ,
    \ces_5_3_io_ins_down[32] ,
    \ces_5_3_io_ins_down[31] ,
    \ces_5_3_io_ins_down[30] ,
    \ces_5_3_io_ins_down[29] ,
    \ces_5_3_io_ins_down[28] ,
    \ces_5_3_io_ins_down[27] ,
    \ces_5_3_io_ins_down[26] ,
    \ces_5_3_io_ins_down[25] ,
    \ces_5_3_io_ins_down[24] ,
    \ces_5_3_io_ins_down[23] ,
    \ces_5_3_io_ins_down[22] ,
    \ces_5_3_io_ins_down[21] ,
    \ces_5_3_io_ins_down[20] ,
    \ces_5_3_io_ins_down[19] ,
    \ces_5_3_io_ins_down[18] ,
    \ces_5_3_io_ins_down[17] ,
    \ces_5_3_io_ins_down[16] ,
    \ces_5_3_io_ins_down[15] ,
    \ces_5_3_io_ins_down[14] ,
    \ces_5_3_io_ins_down[13] ,
    \ces_5_3_io_ins_down[12] ,
    \ces_5_3_io_ins_down[11] ,
    \ces_5_3_io_ins_down[10] ,
    \ces_5_3_io_ins_down[9] ,
    \ces_5_3_io_ins_down[8] ,
    \ces_5_3_io_ins_down[7] ,
    \ces_5_3_io_ins_down[6] ,
    \ces_5_3_io_ins_down[5] ,
    \ces_5_3_io_ins_down[4] ,
    \ces_5_3_io_ins_down[3] ,
    \ces_5_3_io_ins_down[2] ,
    \ces_5_3_io_ins_down[1] ,
    \ces_5_3_io_ins_down[0] }),
    .io_ins_left({\ces_5_3_io_ins_left[63] ,
    \ces_5_3_io_ins_left[62] ,
    \ces_5_3_io_ins_left[61] ,
    \ces_5_3_io_ins_left[60] ,
    \ces_5_3_io_ins_left[59] ,
    \ces_5_3_io_ins_left[58] ,
    \ces_5_3_io_ins_left[57] ,
    \ces_5_3_io_ins_left[56] ,
    \ces_5_3_io_ins_left[55] ,
    \ces_5_3_io_ins_left[54] ,
    \ces_5_3_io_ins_left[53] ,
    \ces_5_3_io_ins_left[52] ,
    \ces_5_3_io_ins_left[51] ,
    \ces_5_3_io_ins_left[50] ,
    \ces_5_3_io_ins_left[49] ,
    \ces_5_3_io_ins_left[48] ,
    \ces_5_3_io_ins_left[47] ,
    \ces_5_3_io_ins_left[46] ,
    \ces_5_3_io_ins_left[45] ,
    \ces_5_3_io_ins_left[44] ,
    \ces_5_3_io_ins_left[43] ,
    \ces_5_3_io_ins_left[42] ,
    \ces_5_3_io_ins_left[41] ,
    \ces_5_3_io_ins_left[40] ,
    \ces_5_3_io_ins_left[39] ,
    \ces_5_3_io_ins_left[38] ,
    \ces_5_3_io_ins_left[37] ,
    \ces_5_3_io_ins_left[36] ,
    \ces_5_3_io_ins_left[35] ,
    \ces_5_3_io_ins_left[34] ,
    \ces_5_3_io_ins_left[33] ,
    \ces_5_3_io_ins_left[32] ,
    \ces_5_3_io_ins_left[31] ,
    \ces_5_3_io_ins_left[30] ,
    \ces_5_3_io_ins_left[29] ,
    \ces_5_3_io_ins_left[28] ,
    \ces_5_3_io_ins_left[27] ,
    \ces_5_3_io_ins_left[26] ,
    \ces_5_3_io_ins_left[25] ,
    \ces_5_3_io_ins_left[24] ,
    \ces_5_3_io_ins_left[23] ,
    \ces_5_3_io_ins_left[22] ,
    \ces_5_3_io_ins_left[21] ,
    \ces_5_3_io_ins_left[20] ,
    \ces_5_3_io_ins_left[19] ,
    \ces_5_3_io_ins_left[18] ,
    \ces_5_3_io_ins_left[17] ,
    \ces_5_3_io_ins_left[16] ,
    \ces_5_3_io_ins_left[15] ,
    \ces_5_3_io_ins_left[14] ,
    \ces_5_3_io_ins_left[13] ,
    \ces_5_3_io_ins_left[12] ,
    \ces_5_3_io_ins_left[11] ,
    \ces_5_3_io_ins_left[10] ,
    \ces_5_3_io_ins_left[9] ,
    \ces_5_3_io_ins_left[8] ,
    \ces_5_3_io_ins_left[7] ,
    \ces_5_3_io_ins_left[6] ,
    \ces_5_3_io_ins_left[5] ,
    \ces_5_3_io_ins_left[4] ,
    \ces_5_3_io_ins_left[3] ,
    \ces_5_3_io_ins_left[2] ,
    \ces_5_3_io_ins_left[1] ,
    \ces_5_3_io_ins_left[0] }),
    .io_ins_right({\ces_5_2_io_outs_right[63] ,
    \ces_5_2_io_outs_right[62] ,
    \ces_5_2_io_outs_right[61] ,
    \ces_5_2_io_outs_right[60] ,
    \ces_5_2_io_outs_right[59] ,
    \ces_5_2_io_outs_right[58] ,
    \ces_5_2_io_outs_right[57] ,
    \ces_5_2_io_outs_right[56] ,
    \ces_5_2_io_outs_right[55] ,
    \ces_5_2_io_outs_right[54] ,
    \ces_5_2_io_outs_right[53] ,
    \ces_5_2_io_outs_right[52] ,
    \ces_5_2_io_outs_right[51] ,
    \ces_5_2_io_outs_right[50] ,
    \ces_5_2_io_outs_right[49] ,
    \ces_5_2_io_outs_right[48] ,
    \ces_5_2_io_outs_right[47] ,
    \ces_5_2_io_outs_right[46] ,
    \ces_5_2_io_outs_right[45] ,
    \ces_5_2_io_outs_right[44] ,
    \ces_5_2_io_outs_right[43] ,
    \ces_5_2_io_outs_right[42] ,
    \ces_5_2_io_outs_right[41] ,
    \ces_5_2_io_outs_right[40] ,
    \ces_5_2_io_outs_right[39] ,
    \ces_5_2_io_outs_right[38] ,
    \ces_5_2_io_outs_right[37] ,
    \ces_5_2_io_outs_right[36] ,
    \ces_5_2_io_outs_right[35] ,
    \ces_5_2_io_outs_right[34] ,
    \ces_5_2_io_outs_right[33] ,
    \ces_5_2_io_outs_right[32] ,
    \ces_5_2_io_outs_right[31] ,
    \ces_5_2_io_outs_right[30] ,
    \ces_5_2_io_outs_right[29] ,
    \ces_5_2_io_outs_right[28] ,
    \ces_5_2_io_outs_right[27] ,
    \ces_5_2_io_outs_right[26] ,
    \ces_5_2_io_outs_right[25] ,
    \ces_5_2_io_outs_right[24] ,
    \ces_5_2_io_outs_right[23] ,
    \ces_5_2_io_outs_right[22] ,
    \ces_5_2_io_outs_right[21] ,
    \ces_5_2_io_outs_right[20] ,
    \ces_5_2_io_outs_right[19] ,
    \ces_5_2_io_outs_right[18] ,
    \ces_5_2_io_outs_right[17] ,
    \ces_5_2_io_outs_right[16] ,
    \ces_5_2_io_outs_right[15] ,
    \ces_5_2_io_outs_right[14] ,
    \ces_5_2_io_outs_right[13] ,
    \ces_5_2_io_outs_right[12] ,
    \ces_5_2_io_outs_right[11] ,
    \ces_5_2_io_outs_right[10] ,
    \ces_5_2_io_outs_right[9] ,
    \ces_5_2_io_outs_right[8] ,
    \ces_5_2_io_outs_right[7] ,
    \ces_5_2_io_outs_right[6] ,
    \ces_5_2_io_outs_right[5] ,
    \ces_5_2_io_outs_right[4] ,
    \ces_5_2_io_outs_right[3] ,
    \ces_5_2_io_outs_right[2] ,
    \ces_5_2_io_outs_right[1] ,
    \ces_5_2_io_outs_right[0] }),
    .io_ins_up({\ces_4_3_io_outs_up[63] ,
    \ces_4_3_io_outs_up[62] ,
    \ces_4_3_io_outs_up[61] ,
    \ces_4_3_io_outs_up[60] ,
    \ces_4_3_io_outs_up[59] ,
    \ces_4_3_io_outs_up[58] ,
    \ces_4_3_io_outs_up[57] ,
    \ces_4_3_io_outs_up[56] ,
    \ces_4_3_io_outs_up[55] ,
    \ces_4_3_io_outs_up[54] ,
    \ces_4_3_io_outs_up[53] ,
    \ces_4_3_io_outs_up[52] ,
    \ces_4_3_io_outs_up[51] ,
    \ces_4_3_io_outs_up[50] ,
    \ces_4_3_io_outs_up[49] ,
    \ces_4_3_io_outs_up[48] ,
    \ces_4_3_io_outs_up[47] ,
    \ces_4_3_io_outs_up[46] ,
    \ces_4_3_io_outs_up[45] ,
    \ces_4_3_io_outs_up[44] ,
    \ces_4_3_io_outs_up[43] ,
    \ces_4_3_io_outs_up[42] ,
    \ces_4_3_io_outs_up[41] ,
    \ces_4_3_io_outs_up[40] ,
    \ces_4_3_io_outs_up[39] ,
    \ces_4_3_io_outs_up[38] ,
    \ces_4_3_io_outs_up[37] ,
    \ces_4_3_io_outs_up[36] ,
    \ces_4_3_io_outs_up[35] ,
    \ces_4_3_io_outs_up[34] ,
    \ces_4_3_io_outs_up[33] ,
    \ces_4_3_io_outs_up[32] ,
    \ces_4_3_io_outs_up[31] ,
    \ces_4_3_io_outs_up[30] ,
    \ces_4_3_io_outs_up[29] ,
    \ces_4_3_io_outs_up[28] ,
    \ces_4_3_io_outs_up[27] ,
    \ces_4_3_io_outs_up[26] ,
    \ces_4_3_io_outs_up[25] ,
    \ces_4_3_io_outs_up[24] ,
    \ces_4_3_io_outs_up[23] ,
    \ces_4_3_io_outs_up[22] ,
    \ces_4_3_io_outs_up[21] ,
    \ces_4_3_io_outs_up[20] ,
    \ces_4_3_io_outs_up[19] ,
    \ces_4_3_io_outs_up[18] ,
    \ces_4_3_io_outs_up[17] ,
    \ces_4_3_io_outs_up[16] ,
    \ces_4_3_io_outs_up[15] ,
    \ces_4_3_io_outs_up[14] ,
    \ces_4_3_io_outs_up[13] ,
    \ces_4_3_io_outs_up[12] ,
    \ces_4_3_io_outs_up[11] ,
    \ces_4_3_io_outs_up[10] ,
    \ces_4_3_io_outs_up[9] ,
    \ces_4_3_io_outs_up[8] ,
    \ces_4_3_io_outs_up[7] ,
    \ces_4_3_io_outs_up[6] ,
    \ces_4_3_io_outs_up[5] ,
    \ces_4_3_io_outs_up[4] ,
    \ces_4_3_io_outs_up[3] ,
    \ces_4_3_io_outs_up[2] ,
    \ces_4_3_io_outs_up[1] ,
    \ces_4_3_io_outs_up[0] }),
    .io_outs_down({\ces_4_3_io_ins_down[63] ,
    \ces_4_3_io_ins_down[62] ,
    \ces_4_3_io_ins_down[61] ,
    \ces_4_3_io_ins_down[60] ,
    \ces_4_3_io_ins_down[59] ,
    \ces_4_3_io_ins_down[58] ,
    \ces_4_3_io_ins_down[57] ,
    \ces_4_3_io_ins_down[56] ,
    \ces_4_3_io_ins_down[55] ,
    \ces_4_3_io_ins_down[54] ,
    \ces_4_3_io_ins_down[53] ,
    \ces_4_3_io_ins_down[52] ,
    \ces_4_3_io_ins_down[51] ,
    \ces_4_3_io_ins_down[50] ,
    \ces_4_3_io_ins_down[49] ,
    \ces_4_3_io_ins_down[48] ,
    \ces_4_3_io_ins_down[47] ,
    \ces_4_3_io_ins_down[46] ,
    \ces_4_3_io_ins_down[45] ,
    \ces_4_3_io_ins_down[44] ,
    \ces_4_3_io_ins_down[43] ,
    \ces_4_3_io_ins_down[42] ,
    \ces_4_3_io_ins_down[41] ,
    \ces_4_3_io_ins_down[40] ,
    \ces_4_3_io_ins_down[39] ,
    \ces_4_3_io_ins_down[38] ,
    \ces_4_3_io_ins_down[37] ,
    \ces_4_3_io_ins_down[36] ,
    \ces_4_3_io_ins_down[35] ,
    \ces_4_3_io_ins_down[34] ,
    \ces_4_3_io_ins_down[33] ,
    \ces_4_3_io_ins_down[32] ,
    \ces_4_3_io_ins_down[31] ,
    \ces_4_3_io_ins_down[30] ,
    \ces_4_3_io_ins_down[29] ,
    \ces_4_3_io_ins_down[28] ,
    \ces_4_3_io_ins_down[27] ,
    \ces_4_3_io_ins_down[26] ,
    \ces_4_3_io_ins_down[25] ,
    \ces_4_3_io_ins_down[24] ,
    \ces_4_3_io_ins_down[23] ,
    \ces_4_3_io_ins_down[22] ,
    \ces_4_3_io_ins_down[21] ,
    \ces_4_3_io_ins_down[20] ,
    \ces_4_3_io_ins_down[19] ,
    \ces_4_3_io_ins_down[18] ,
    \ces_4_3_io_ins_down[17] ,
    \ces_4_3_io_ins_down[16] ,
    \ces_4_3_io_ins_down[15] ,
    \ces_4_3_io_ins_down[14] ,
    \ces_4_3_io_ins_down[13] ,
    \ces_4_3_io_ins_down[12] ,
    \ces_4_3_io_ins_down[11] ,
    \ces_4_3_io_ins_down[10] ,
    \ces_4_3_io_ins_down[9] ,
    \ces_4_3_io_ins_down[8] ,
    \ces_4_3_io_ins_down[7] ,
    \ces_4_3_io_ins_down[6] ,
    \ces_4_3_io_ins_down[5] ,
    \ces_4_3_io_ins_down[4] ,
    \ces_4_3_io_ins_down[3] ,
    \ces_4_3_io_ins_down[2] ,
    \ces_4_3_io_ins_down[1] ,
    \ces_4_3_io_ins_down[0] }),
    .io_outs_left({\ces_5_2_io_ins_left[63] ,
    \ces_5_2_io_ins_left[62] ,
    \ces_5_2_io_ins_left[61] ,
    \ces_5_2_io_ins_left[60] ,
    \ces_5_2_io_ins_left[59] ,
    \ces_5_2_io_ins_left[58] ,
    \ces_5_2_io_ins_left[57] ,
    \ces_5_2_io_ins_left[56] ,
    \ces_5_2_io_ins_left[55] ,
    \ces_5_2_io_ins_left[54] ,
    \ces_5_2_io_ins_left[53] ,
    \ces_5_2_io_ins_left[52] ,
    \ces_5_2_io_ins_left[51] ,
    \ces_5_2_io_ins_left[50] ,
    \ces_5_2_io_ins_left[49] ,
    \ces_5_2_io_ins_left[48] ,
    \ces_5_2_io_ins_left[47] ,
    \ces_5_2_io_ins_left[46] ,
    \ces_5_2_io_ins_left[45] ,
    \ces_5_2_io_ins_left[44] ,
    \ces_5_2_io_ins_left[43] ,
    \ces_5_2_io_ins_left[42] ,
    \ces_5_2_io_ins_left[41] ,
    \ces_5_2_io_ins_left[40] ,
    \ces_5_2_io_ins_left[39] ,
    \ces_5_2_io_ins_left[38] ,
    \ces_5_2_io_ins_left[37] ,
    \ces_5_2_io_ins_left[36] ,
    \ces_5_2_io_ins_left[35] ,
    \ces_5_2_io_ins_left[34] ,
    \ces_5_2_io_ins_left[33] ,
    \ces_5_2_io_ins_left[32] ,
    \ces_5_2_io_ins_left[31] ,
    \ces_5_2_io_ins_left[30] ,
    \ces_5_2_io_ins_left[29] ,
    \ces_5_2_io_ins_left[28] ,
    \ces_5_2_io_ins_left[27] ,
    \ces_5_2_io_ins_left[26] ,
    \ces_5_2_io_ins_left[25] ,
    \ces_5_2_io_ins_left[24] ,
    \ces_5_2_io_ins_left[23] ,
    \ces_5_2_io_ins_left[22] ,
    \ces_5_2_io_ins_left[21] ,
    \ces_5_2_io_ins_left[20] ,
    \ces_5_2_io_ins_left[19] ,
    \ces_5_2_io_ins_left[18] ,
    \ces_5_2_io_ins_left[17] ,
    \ces_5_2_io_ins_left[16] ,
    \ces_5_2_io_ins_left[15] ,
    \ces_5_2_io_ins_left[14] ,
    \ces_5_2_io_ins_left[13] ,
    \ces_5_2_io_ins_left[12] ,
    \ces_5_2_io_ins_left[11] ,
    \ces_5_2_io_ins_left[10] ,
    \ces_5_2_io_ins_left[9] ,
    \ces_5_2_io_ins_left[8] ,
    \ces_5_2_io_ins_left[7] ,
    \ces_5_2_io_ins_left[6] ,
    \ces_5_2_io_ins_left[5] ,
    \ces_5_2_io_ins_left[4] ,
    \ces_5_2_io_ins_left[3] ,
    \ces_5_2_io_ins_left[2] ,
    \ces_5_2_io_ins_left[1] ,
    \ces_5_2_io_ins_left[0] }),
    .io_outs_right({\ces_5_3_io_outs_right[63] ,
    \ces_5_3_io_outs_right[62] ,
    \ces_5_3_io_outs_right[61] ,
    \ces_5_3_io_outs_right[60] ,
    \ces_5_3_io_outs_right[59] ,
    \ces_5_3_io_outs_right[58] ,
    \ces_5_3_io_outs_right[57] ,
    \ces_5_3_io_outs_right[56] ,
    \ces_5_3_io_outs_right[55] ,
    \ces_5_3_io_outs_right[54] ,
    \ces_5_3_io_outs_right[53] ,
    \ces_5_3_io_outs_right[52] ,
    \ces_5_3_io_outs_right[51] ,
    \ces_5_3_io_outs_right[50] ,
    \ces_5_3_io_outs_right[49] ,
    \ces_5_3_io_outs_right[48] ,
    \ces_5_3_io_outs_right[47] ,
    \ces_5_3_io_outs_right[46] ,
    \ces_5_3_io_outs_right[45] ,
    \ces_5_3_io_outs_right[44] ,
    \ces_5_3_io_outs_right[43] ,
    \ces_5_3_io_outs_right[42] ,
    \ces_5_3_io_outs_right[41] ,
    \ces_5_3_io_outs_right[40] ,
    \ces_5_3_io_outs_right[39] ,
    \ces_5_3_io_outs_right[38] ,
    \ces_5_3_io_outs_right[37] ,
    \ces_5_3_io_outs_right[36] ,
    \ces_5_3_io_outs_right[35] ,
    \ces_5_3_io_outs_right[34] ,
    \ces_5_3_io_outs_right[33] ,
    \ces_5_3_io_outs_right[32] ,
    \ces_5_3_io_outs_right[31] ,
    \ces_5_3_io_outs_right[30] ,
    \ces_5_3_io_outs_right[29] ,
    \ces_5_3_io_outs_right[28] ,
    \ces_5_3_io_outs_right[27] ,
    \ces_5_3_io_outs_right[26] ,
    \ces_5_3_io_outs_right[25] ,
    \ces_5_3_io_outs_right[24] ,
    \ces_5_3_io_outs_right[23] ,
    \ces_5_3_io_outs_right[22] ,
    \ces_5_3_io_outs_right[21] ,
    \ces_5_3_io_outs_right[20] ,
    \ces_5_3_io_outs_right[19] ,
    \ces_5_3_io_outs_right[18] ,
    \ces_5_3_io_outs_right[17] ,
    \ces_5_3_io_outs_right[16] ,
    \ces_5_3_io_outs_right[15] ,
    \ces_5_3_io_outs_right[14] ,
    \ces_5_3_io_outs_right[13] ,
    \ces_5_3_io_outs_right[12] ,
    \ces_5_3_io_outs_right[11] ,
    \ces_5_3_io_outs_right[10] ,
    \ces_5_3_io_outs_right[9] ,
    \ces_5_3_io_outs_right[8] ,
    \ces_5_3_io_outs_right[7] ,
    \ces_5_3_io_outs_right[6] ,
    \ces_5_3_io_outs_right[5] ,
    \ces_5_3_io_outs_right[4] ,
    \ces_5_3_io_outs_right[3] ,
    \ces_5_3_io_outs_right[2] ,
    \ces_5_3_io_outs_right[1] ,
    \ces_5_3_io_outs_right[0] }),
    .io_outs_up({\ces_5_3_io_outs_up[63] ,
    \ces_5_3_io_outs_up[62] ,
    \ces_5_3_io_outs_up[61] ,
    \ces_5_3_io_outs_up[60] ,
    \ces_5_3_io_outs_up[59] ,
    \ces_5_3_io_outs_up[58] ,
    \ces_5_3_io_outs_up[57] ,
    \ces_5_3_io_outs_up[56] ,
    \ces_5_3_io_outs_up[55] ,
    \ces_5_3_io_outs_up[54] ,
    \ces_5_3_io_outs_up[53] ,
    \ces_5_3_io_outs_up[52] ,
    \ces_5_3_io_outs_up[51] ,
    \ces_5_3_io_outs_up[50] ,
    \ces_5_3_io_outs_up[49] ,
    \ces_5_3_io_outs_up[48] ,
    \ces_5_3_io_outs_up[47] ,
    \ces_5_3_io_outs_up[46] ,
    \ces_5_3_io_outs_up[45] ,
    \ces_5_3_io_outs_up[44] ,
    \ces_5_3_io_outs_up[43] ,
    \ces_5_3_io_outs_up[42] ,
    \ces_5_3_io_outs_up[41] ,
    \ces_5_3_io_outs_up[40] ,
    \ces_5_3_io_outs_up[39] ,
    \ces_5_3_io_outs_up[38] ,
    \ces_5_3_io_outs_up[37] ,
    \ces_5_3_io_outs_up[36] ,
    \ces_5_3_io_outs_up[35] ,
    \ces_5_3_io_outs_up[34] ,
    \ces_5_3_io_outs_up[33] ,
    \ces_5_3_io_outs_up[32] ,
    \ces_5_3_io_outs_up[31] ,
    \ces_5_3_io_outs_up[30] ,
    \ces_5_3_io_outs_up[29] ,
    \ces_5_3_io_outs_up[28] ,
    \ces_5_3_io_outs_up[27] ,
    \ces_5_3_io_outs_up[26] ,
    \ces_5_3_io_outs_up[25] ,
    \ces_5_3_io_outs_up[24] ,
    \ces_5_3_io_outs_up[23] ,
    \ces_5_3_io_outs_up[22] ,
    \ces_5_3_io_outs_up[21] ,
    \ces_5_3_io_outs_up[20] ,
    \ces_5_3_io_outs_up[19] ,
    \ces_5_3_io_outs_up[18] ,
    \ces_5_3_io_outs_up[17] ,
    \ces_5_3_io_outs_up[16] ,
    \ces_5_3_io_outs_up[15] ,
    \ces_5_3_io_outs_up[14] ,
    \ces_5_3_io_outs_up[13] ,
    \ces_5_3_io_outs_up[12] ,
    \ces_5_3_io_outs_up[11] ,
    \ces_5_3_io_outs_up[10] ,
    \ces_5_3_io_outs_up[9] ,
    \ces_5_3_io_outs_up[8] ,
    \ces_5_3_io_outs_up[7] ,
    \ces_5_3_io_outs_up[6] ,
    \ces_5_3_io_outs_up[5] ,
    \ces_5_3_io_outs_up[4] ,
    \ces_5_3_io_outs_up[3] ,
    \ces_5_3_io_outs_up[2] ,
    \ces_5_3_io_outs_up[1] ,
    \ces_5_3_io_outs_up[0] }));
 Element ces_5_4 (.clock(clknet_3_6_0_clock),
    .io_lsbIns_1(ces_5_3_io_lsbOuts_1),
    .io_lsbIns_2(ces_5_3_io_lsbOuts_2),
    .io_lsbIns_3(ces_5_3_io_lsbOuts_3),
    .io_lsbIns_4(ces_5_3_io_lsbOuts_4),
    .io_lsbIns_5(ces_5_3_io_lsbOuts_5),
    .io_lsbIns_6(ces_5_3_io_lsbOuts_6),
    .io_lsbIns_7(ces_5_3_io_lsbOuts_7),
    .io_lsbOuts_0(ces_5_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_4_io_lsbOuts_7),
    .io_ins_down({\ces_5_4_io_ins_down[63] ,
    \ces_5_4_io_ins_down[62] ,
    \ces_5_4_io_ins_down[61] ,
    \ces_5_4_io_ins_down[60] ,
    \ces_5_4_io_ins_down[59] ,
    \ces_5_4_io_ins_down[58] ,
    \ces_5_4_io_ins_down[57] ,
    \ces_5_4_io_ins_down[56] ,
    \ces_5_4_io_ins_down[55] ,
    \ces_5_4_io_ins_down[54] ,
    \ces_5_4_io_ins_down[53] ,
    \ces_5_4_io_ins_down[52] ,
    \ces_5_4_io_ins_down[51] ,
    \ces_5_4_io_ins_down[50] ,
    \ces_5_4_io_ins_down[49] ,
    \ces_5_4_io_ins_down[48] ,
    \ces_5_4_io_ins_down[47] ,
    \ces_5_4_io_ins_down[46] ,
    \ces_5_4_io_ins_down[45] ,
    \ces_5_4_io_ins_down[44] ,
    \ces_5_4_io_ins_down[43] ,
    \ces_5_4_io_ins_down[42] ,
    \ces_5_4_io_ins_down[41] ,
    \ces_5_4_io_ins_down[40] ,
    \ces_5_4_io_ins_down[39] ,
    \ces_5_4_io_ins_down[38] ,
    \ces_5_4_io_ins_down[37] ,
    \ces_5_4_io_ins_down[36] ,
    \ces_5_4_io_ins_down[35] ,
    \ces_5_4_io_ins_down[34] ,
    \ces_5_4_io_ins_down[33] ,
    \ces_5_4_io_ins_down[32] ,
    \ces_5_4_io_ins_down[31] ,
    \ces_5_4_io_ins_down[30] ,
    \ces_5_4_io_ins_down[29] ,
    \ces_5_4_io_ins_down[28] ,
    \ces_5_4_io_ins_down[27] ,
    \ces_5_4_io_ins_down[26] ,
    \ces_5_4_io_ins_down[25] ,
    \ces_5_4_io_ins_down[24] ,
    \ces_5_4_io_ins_down[23] ,
    \ces_5_4_io_ins_down[22] ,
    \ces_5_4_io_ins_down[21] ,
    \ces_5_4_io_ins_down[20] ,
    \ces_5_4_io_ins_down[19] ,
    \ces_5_4_io_ins_down[18] ,
    \ces_5_4_io_ins_down[17] ,
    \ces_5_4_io_ins_down[16] ,
    \ces_5_4_io_ins_down[15] ,
    \ces_5_4_io_ins_down[14] ,
    \ces_5_4_io_ins_down[13] ,
    \ces_5_4_io_ins_down[12] ,
    \ces_5_4_io_ins_down[11] ,
    \ces_5_4_io_ins_down[10] ,
    \ces_5_4_io_ins_down[9] ,
    \ces_5_4_io_ins_down[8] ,
    \ces_5_4_io_ins_down[7] ,
    \ces_5_4_io_ins_down[6] ,
    \ces_5_4_io_ins_down[5] ,
    \ces_5_4_io_ins_down[4] ,
    \ces_5_4_io_ins_down[3] ,
    \ces_5_4_io_ins_down[2] ,
    \ces_5_4_io_ins_down[1] ,
    \ces_5_4_io_ins_down[0] }),
    .io_ins_left({\ces_5_4_io_ins_left[63] ,
    \ces_5_4_io_ins_left[62] ,
    \ces_5_4_io_ins_left[61] ,
    \ces_5_4_io_ins_left[60] ,
    \ces_5_4_io_ins_left[59] ,
    \ces_5_4_io_ins_left[58] ,
    \ces_5_4_io_ins_left[57] ,
    \ces_5_4_io_ins_left[56] ,
    \ces_5_4_io_ins_left[55] ,
    \ces_5_4_io_ins_left[54] ,
    \ces_5_4_io_ins_left[53] ,
    \ces_5_4_io_ins_left[52] ,
    \ces_5_4_io_ins_left[51] ,
    \ces_5_4_io_ins_left[50] ,
    \ces_5_4_io_ins_left[49] ,
    \ces_5_4_io_ins_left[48] ,
    \ces_5_4_io_ins_left[47] ,
    \ces_5_4_io_ins_left[46] ,
    \ces_5_4_io_ins_left[45] ,
    \ces_5_4_io_ins_left[44] ,
    \ces_5_4_io_ins_left[43] ,
    \ces_5_4_io_ins_left[42] ,
    \ces_5_4_io_ins_left[41] ,
    \ces_5_4_io_ins_left[40] ,
    \ces_5_4_io_ins_left[39] ,
    \ces_5_4_io_ins_left[38] ,
    \ces_5_4_io_ins_left[37] ,
    \ces_5_4_io_ins_left[36] ,
    \ces_5_4_io_ins_left[35] ,
    \ces_5_4_io_ins_left[34] ,
    \ces_5_4_io_ins_left[33] ,
    \ces_5_4_io_ins_left[32] ,
    \ces_5_4_io_ins_left[31] ,
    \ces_5_4_io_ins_left[30] ,
    \ces_5_4_io_ins_left[29] ,
    \ces_5_4_io_ins_left[28] ,
    \ces_5_4_io_ins_left[27] ,
    \ces_5_4_io_ins_left[26] ,
    \ces_5_4_io_ins_left[25] ,
    \ces_5_4_io_ins_left[24] ,
    \ces_5_4_io_ins_left[23] ,
    \ces_5_4_io_ins_left[22] ,
    \ces_5_4_io_ins_left[21] ,
    \ces_5_4_io_ins_left[20] ,
    \ces_5_4_io_ins_left[19] ,
    \ces_5_4_io_ins_left[18] ,
    \ces_5_4_io_ins_left[17] ,
    \ces_5_4_io_ins_left[16] ,
    \ces_5_4_io_ins_left[15] ,
    \ces_5_4_io_ins_left[14] ,
    \ces_5_4_io_ins_left[13] ,
    \ces_5_4_io_ins_left[12] ,
    \ces_5_4_io_ins_left[11] ,
    \ces_5_4_io_ins_left[10] ,
    \ces_5_4_io_ins_left[9] ,
    \ces_5_4_io_ins_left[8] ,
    \ces_5_4_io_ins_left[7] ,
    \ces_5_4_io_ins_left[6] ,
    \ces_5_4_io_ins_left[5] ,
    \ces_5_4_io_ins_left[4] ,
    \ces_5_4_io_ins_left[3] ,
    \ces_5_4_io_ins_left[2] ,
    \ces_5_4_io_ins_left[1] ,
    \ces_5_4_io_ins_left[0] }),
    .io_ins_right({\ces_5_3_io_outs_right[63] ,
    \ces_5_3_io_outs_right[62] ,
    \ces_5_3_io_outs_right[61] ,
    \ces_5_3_io_outs_right[60] ,
    \ces_5_3_io_outs_right[59] ,
    \ces_5_3_io_outs_right[58] ,
    \ces_5_3_io_outs_right[57] ,
    \ces_5_3_io_outs_right[56] ,
    \ces_5_3_io_outs_right[55] ,
    \ces_5_3_io_outs_right[54] ,
    \ces_5_3_io_outs_right[53] ,
    \ces_5_3_io_outs_right[52] ,
    \ces_5_3_io_outs_right[51] ,
    \ces_5_3_io_outs_right[50] ,
    \ces_5_3_io_outs_right[49] ,
    \ces_5_3_io_outs_right[48] ,
    \ces_5_3_io_outs_right[47] ,
    \ces_5_3_io_outs_right[46] ,
    \ces_5_3_io_outs_right[45] ,
    \ces_5_3_io_outs_right[44] ,
    \ces_5_3_io_outs_right[43] ,
    \ces_5_3_io_outs_right[42] ,
    \ces_5_3_io_outs_right[41] ,
    \ces_5_3_io_outs_right[40] ,
    \ces_5_3_io_outs_right[39] ,
    \ces_5_3_io_outs_right[38] ,
    \ces_5_3_io_outs_right[37] ,
    \ces_5_3_io_outs_right[36] ,
    \ces_5_3_io_outs_right[35] ,
    \ces_5_3_io_outs_right[34] ,
    \ces_5_3_io_outs_right[33] ,
    \ces_5_3_io_outs_right[32] ,
    \ces_5_3_io_outs_right[31] ,
    \ces_5_3_io_outs_right[30] ,
    \ces_5_3_io_outs_right[29] ,
    \ces_5_3_io_outs_right[28] ,
    \ces_5_3_io_outs_right[27] ,
    \ces_5_3_io_outs_right[26] ,
    \ces_5_3_io_outs_right[25] ,
    \ces_5_3_io_outs_right[24] ,
    \ces_5_3_io_outs_right[23] ,
    \ces_5_3_io_outs_right[22] ,
    \ces_5_3_io_outs_right[21] ,
    \ces_5_3_io_outs_right[20] ,
    \ces_5_3_io_outs_right[19] ,
    \ces_5_3_io_outs_right[18] ,
    \ces_5_3_io_outs_right[17] ,
    \ces_5_3_io_outs_right[16] ,
    \ces_5_3_io_outs_right[15] ,
    \ces_5_3_io_outs_right[14] ,
    \ces_5_3_io_outs_right[13] ,
    \ces_5_3_io_outs_right[12] ,
    \ces_5_3_io_outs_right[11] ,
    \ces_5_3_io_outs_right[10] ,
    \ces_5_3_io_outs_right[9] ,
    \ces_5_3_io_outs_right[8] ,
    \ces_5_3_io_outs_right[7] ,
    \ces_5_3_io_outs_right[6] ,
    \ces_5_3_io_outs_right[5] ,
    \ces_5_3_io_outs_right[4] ,
    \ces_5_3_io_outs_right[3] ,
    \ces_5_3_io_outs_right[2] ,
    \ces_5_3_io_outs_right[1] ,
    \ces_5_3_io_outs_right[0] }),
    .io_ins_up({\ces_4_4_io_outs_up[63] ,
    \ces_4_4_io_outs_up[62] ,
    \ces_4_4_io_outs_up[61] ,
    \ces_4_4_io_outs_up[60] ,
    \ces_4_4_io_outs_up[59] ,
    \ces_4_4_io_outs_up[58] ,
    \ces_4_4_io_outs_up[57] ,
    \ces_4_4_io_outs_up[56] ,
    \ces_4_4_io_outs_up[55] ,
    \ces_4_4_io_outs_up[54] ,
    \ces_4_4_io_outs_up[53] ,
    \ces_4_4_io_outs_up[52] ,
    \ces_4_4_io_outs_up[51] ,
    \ces_4_4_io_outs_up[50] ,
    \ces_4_4_io_outs_up[49] ,
    \ces_4_4_io_outs_up[48] ,
    \ces_4_4_io_outs_up[47] ,
    \ces_4_4_io_outs_up[46] ,
    \ces_4_4_io_outs_up[45] ,
    \ces_4_4_io_outs_up[44] ,
    \ces_4_4_io_outs_up[43] ,
    \ces_4_4_io_outs_up[42] ,
    \ces_4_4_io_outs_up[41] ,
    \ces_4_4_io_outs_up[40] ,
    \ces_4_4_io_outs_up[39] ,
    \ces_4_4_io_outs_up[38] ,
    \ces_4_4_io_outs_up[37] ,
    \ces_4_4_io_outs_up[36] ,
    \ces_4_4_io_outs_up[35] ,
    \ces_4_4_io_outs_up[34] ,
    \ces_4_4_io_outs_up[33] ,
    \ces_4_4_io_outs_up[32] ,
    \ces_4_4_io_outs_up[31] ,
    \ces_4_4_io_outs_up[30] ,
    \ces_4_4_io_outs_up[29] ,
    \ces_4_4_io_outs_up[28] ,
    \ces_4_4_io_outs_up[27] ,
    \ces_4_4_io_outs_up[26] ,
    \ces_4_4_io_outs_up[25] ,
    \ces_4_4_io_outs_up[24] ,
    \ces_4_4_io_outs_up[23] ,
    \ces_4_4_io_outs_up[22] ,
    \ces_4_4_io_outs_up[21] ,
    \ces_4_4_io_outs_up[20] ,
    \ces_4_4_io_outs_up[19] ,
    \ces_4_4_io_outs_up[18] ,
    \ces_4_4_io_outs_up[17] ,
    \ces_4_4_io_outs_up[16] ,
    \ces_4_4_io_outs_up[15] ,
    \ces_4_4_io_outs_up[14] ,
    \ces_4_4_io_outs_up[13] ,
    \ces_4_4_io_outs_up[12] ,
    \ces_4_4_io_outs_up[11] ,
    \ces_4_4_io_outs_up[10] ,
    \ces_4_4_io_outs_up[9] ,
    \ces_4_4_io_outs_up[8] ,
    \ces_4_4_io_outs_up[7] ,
    \ces_4_4_io_outs_up[6] ,
    \ces_4_4_io_outs_up[5] ,
    \ces_4_4_io_outs_up[4] ,
    \ces_4_4_io_outs_up[3] ,
    \ces_4_4_io_outs_up[2] ,
    \ces_4_4_io_outs_up[1] ,
    \ces_4_4_io_outs_up[0] }),
    .io_outs_down({\ces_4_4_io_ins_down[63] ,
    \ces_4_4_io_ins_down[62] ,
    \ces_4_4_io_ins_down[61] ,
    \ces_4_4_io_ins_down[60] ,
    \ces_4_4_io_ins_down[59] ,
    \ces_4_4_io_ins_down[58] ,
    \ces_4_4_io_ins_down[57] ,
    \ces_4_4_io_ins_down[56] ,
    \ces_4_4_io_ins_down[55] ,
    \ces_4_4_io_ins_down[54] ,
    \ces_4_4_io_ins_down[53] ,
    \ces_4_4_io_ins_down[52] ,
    \ces_4_4_io_ins_down[51] ,
    \ces_4_4_io_ins_down[50] ,
    \ces_4_4_io_ins_down[49] ,
    \ces_4_4_io_ins_down[48] ,
    \ces_4_4_io_ins_down[47] ,
    \ces_4_4_io_ins_down[46] ,
    \ces_4_4_io_ins_down[45] ,
    \ces_4_4_io_ins_down[44] ,
    \ces_4_4_io_ins_down[43] ,
    \ces_4_4_io_ins_down[42] ,
    \ces_4_4_io_ins_down[41] ,
    \ces_4_4_io_ins_down[40] ,
    \ces_4_4_io_ins_down[39] ,
    \ces_4_4_io_ins_down[38] ,
    \ces_4_4_io_ins_down[37] ,
    \ces_4_4_io_ins_down[36] ,
    \ces_4_4_io_ins_down[35] ,
    \ces_4_4_io_ins_down[34] ,
    \ces_4_4_io_ins_down[33] ,
    \ces_4_4_io_ins_down[32] ,
    \ces_4_4_io_ins_down[31] ,
    \ces_4_4_io_ins_down[30] ,
    \ces_4_4_io_ins_down[29] ,
    \ces_4_4_io_ins_down[28] ,
    \ces_4_4_io_ins_down[27] ,
    \ces_4_4_io_ins_down[26] ,
    \ces_4_4_io_ins_down[25] ,
    \ces_4_4_io_ins_down[24] ,
    \ces_4_4_io_ins_down[23] ,
    \ces_4_4_io_ins_down[22] ,
    \ces_4_4_io_ins_down[21] ,
    \ces_4_4_io_ins_down[20] ,
    \ces_4_4_io_ins_down[19] ,
    \ces_4_4_io_ins_down[18] ,
    \ces_4_4_io_ins_down[17] ,
    \ces_4_4_io_ins_down[16] ,
    \ces_4_4_io_ins_down[15] ,
    \ces_4_4_io_ins_down[14] ,
    \ces_4_4_io_ins_down[13] ,
    \ces_4_4_io_ins_down[12] ,
    \ces_4_4_io_ins_down[11] ,
    \ces_4_4_io_ins_down[10] ,
    \ces_4_4_io_ins_down[9] ,
    \ces_4_4_io_ins_down[8] ,
    \ces_4_4_io_ins_down[7] ,
    \ces_4_4_io_ins_down[6] ,
    \ces_4_4_io_ins_down[5] ,
    \ces_4_4_io_ins_down[4] ,
    \ces_4_4_io_ins_down[3] ,
    \ces_4_4_io_ins_down[2] ,
    \ces_4_4_io_ins_down[1] ,
    \ces_4_4_io_ins_down[0] }),
    .io_outs_left({\ces_5_3_io_ins_left[63] ,
    \ces_5_3_io_ins_left[62] ,
    \ces_5_3_io_ins_left[61] ,
    \ces_5_3_io_ins_left[60] ,
    \ces_5_3_io_ins_left[59] ,
    \ces_5_3_io_ins_left[58] ,
    \ces_5_3_io_ins_left[57] ,
    \ces_5_3_io_ins_left[56] ,
    \ces_5_3_io_ins_left[55] ,
    \ces_5_3_io_ins_left[54] ,
    \ces_5_3_io_ins_left[53] ,
    \ces_5_3_io_ins_left[52] ,
    \ces_5_3_io_ins_left[51] ,
    \ces_5_3_io_ins_left[50] ,
    \ces_5_3_io_ins_left[49] ,
    \ces_5_3_io_ins_left[48] ,
    \ces_5_3_io_ins_left[47] ,
    \ces_5_3_io_ins_left[46] ,
    \ces_5_3_io_ins_left[45] ,
    \ces_5_3_io_ins_left[44] ,
    \ces_5_3_io_ins_left[43] ,
    \ces_5_3_io_ins_left[42] ,
    \ces_5_3_io_ins_left[41] ,
    \ces_5_3_io_ins_left[40] ,
    \ces_5_3_io_ins_left[39] ,
    \ces_5_3_io_ins_left[38] ,
    \ces_5_3_io_ins_left[37] ,
    \ces_5_3_io_ins_left[36] ,
    \ces_5_3_io_ins_left[35] ,
    \ces_5_3_io_ins_left[34] ,
    \ces_5_3_io_ins_left[33] ,
    \ces_5_3_io_ins_left[32] ,
    \ces_5_3_io_ins_left[31] ,
    \ces_5_3_io_ins_left[30] ,
    \ces_5_3_io_ins_left[29] ,
    \ces_5_3_io_ins_left[28] ,
    \ces_5_3_io_ins_left[27] ,
    \ces_5_3_io_ins_left[26] ,
    \ces_5_3_io_ins_left[25] ,
    \ces_5_3_io_ins_left[24] ,
    \ces_5_3_io_ins_left[23] ,
    \ces_5_3_io_ins_left[22] ,
    \ces_5_3_io_ins_left[21] ,
    \ces_5_3_io_ins_left[20] ,
    \ces_5_3_io_ins_left[19] ,
    \ces_5_3_io_ins_left[18] ,
    \ces_5_3_io_ins_left[17] ,
    \ces_5_3_io_ins_left[16] ,
    \ces_5_3_io_ins_left[15] ,
    \ces_5_3_io_ins_left[14] ,
    \ces_5_3_io_ins_left[13] ,
    \ces_5_3_io_ins_left[12] ,
    \ces_5_3_io_ins_left[11] ,
    \ces_5_3_io_ins_left[10] ,
    \ces_5_3_io_ins_left[9] ,
    \ces_5_3_io_ins_left[8] ,
    \ces_5_3_io_ins_left[7] ,
    \ces_5_3_io_ins_left[6] ,
    \ces_5_3_io_ins_left[5] ,
    \ces_5_3_io_ins_left[4] ,
    \ces_5_3_io_ins_left[3] ,
    \ces_5_3_io_ins_left[2] ,
    \ces_5_3_io_ins_left[1] ,
    \ces_5_3_io_ins_left[0] }),
    .io_outs_right({\ces_5_4_io_outs_right[63] ,
    \ces_5_4_io_outs_right[62] ,
    \ces_5_4_io_outs_right[61] ,
    \ces_5_4_io_outs_right[60] ,
    \ces_5_4_io_outs_right[59] ,
    \ces_5_4_io_outs_right[58] ,
    \ces_5_4_io_outs_right[57] ,
    \ces_5_4_io_outs_right[56] ,
    \ces_5_4_io_outs_right[55] ,
    \ces_5_4_io_outs_right[54] ,
    \ces_5_4_io_outs_right[53] ,
    \ces_5_4_io_outs_right[52] ,
    \ces_5_4_io_outs_right[51] ,
    \ces_5_4_io_outs_right[50] ,
    \ces_5_4_io_outs_right[49] ,
    \ces_5_4_io_outs_right[48] ,
    \ces_5_4_io_outs_right[47] ,
    \ces_5_4_io_outs_right[46] ,
    \ces_5_4_io_outs_right[45] ,
    \ces_5_4_io_outs_right[44] ,
    \ces_5_4_io_outs_right[43] ,
    \ces_5_4_io_outs_right[42] ,
    \ces_5_4_io_outs_right[41] ,
    \ces_5_4_io_outs_right[40] ,
    \ces_5_4_io_outs_right[39] ,
    \ces_5_4_io_outs_right[38] ,
    \ces_5_4_io_outs_right[37] ,
    \ces_5_4_io_outs_right[36] ,
    \ces_5_4_io_outs_right[35] ,
    \ces_5_4_io_outs_right[34] ,
    \ces_5_4_io_outs_right[33] ,
    \ces_5_4_io_outs_right[32] ,
    \ces_5_4_io_outs_right[31] ,
    \ces_5_4_io_outs_right[30] ,
    \ces_5_4_io_outs_right[29] ,
    \ces_5_4_io_outs_right[28] ,
    \ces_5_4_io_outs_right[27] ,
    \ces_5_4_io_outs_right[26] ,
    \ces_5_4_io_outs_right[25] ,
    \ces_5_4_io_outs_right[24] ,
    \ces_5_4_io_outs_right[23] ,
    \ces_5_4_io_outs_right[22] ,
    \ces_5_4_io_outs_right[21] ,
    \ces_5_4_io_outs_right[20] ,
    \ces_5_4_io_outs_right[19] ,
    \ces_5_4_io_outs_right[18] ,
    \ces_5_4_io_outs_right[17] ,
    \ces_5_4_io_outs_right[16] ,
    \ces_5_4_io_outs_right[15] ,
    \ces_5_4_io_outs_right[14] ,
    \ces_5_4_io_outs_right[13] ,
    \ces_5_4_io_outs_right[12] ,
    \ces_5_4_io_outs_right[11] ,
    \ces_5_4_io_outs_right[10] ,
    \ces_5_4_io_outs_right[9] ,
    \ces_5_4_io_outs_right[8] ,
    \ces_5_4_io_outs_right[7] ,
    \ces_5_4_io_outs_right[6] ,
    \ces_5_4_io_outs_right[5] ,
    \ces_5_4_io_outs_right[4] ,
    \ces_5_4_io_outs_right[3] ,
    \ces_5_4_io_outs_right[2] ,
    \ces_5_4_io_outs_right[1] ,
    \ces_5_4_io_outs_right[0] }),
    .io_outs_up({\ces_5_4_io_outs_up[63] ,
    \ces_5_4_io_outs_up[62] ,
    \ces_5_4_io_outs_up[61] ,
    \ces_5_4_io_outs_up[60] ,
    \ces_5_4_io_outs_up[59] ,
    \ces_5_4_io_outs_up[58] ,
    \ces_5_4_io_outs_up[57] ,
    \ces_5_4_io_outs_up[56] ,
    \ces_5_4_io_outs_up[55] ,
    \ces_5_4_io_outs_up[54] ,
    \ces_5_4_io_outs_up[53] ,
    \ces_5_4_io_outs_up[52] ,
    \ces_5_4_io_outs_up[51] ,
    \ces_5_4_io_outs_up[50] ,
    \ces_5_4_io_outs_up[49] ,
    \ces_5_4_io_outs_up[48] ,
    \ces_5_4_io_outs_up[47] ,
    \ces_5_4_io_outs_up[46] ,
    \ces_5_4_io_outs_up[45] ,
    \ces_5_4_io_outs_up[44] ,
    \ces_5_4_io_outs_up[43] ,
    \ces_5_4_io_outs_up[42] ,
    \ces_5_4_io_outs_up[41] ,
    \ces_5_4_io_outs_up[40] ,
    \ces_5_4_io_outs_up[39] ,
    \ces_5_4_io_outs_up[38] ,
    \ces_5_4_io_outs_up[37] ,
    \ces_5_4_io_outs_up[36] ,
    \ces_5_4_io_outs_up[35] ,
    \ces_5_4_io_outs_up[34] ,
    \ces_5_4_io_outs_up[33] ,
    \ces_5_4_io_outs_up[32] ,
    \ces_5_4_io_outs_up[31] ,
    \ces_5_4_io_outs_up[30] ,
    \ces_5_4_io_outs_up[29] ,
    \ces_5_4_io_outs_up[28] ,
    \ces_5_4_io_outs_up[27] ,
    \ces_5_4_io_outs_up[26] ,
    \ces_5_4_io_outs_up[25] ,
    \ces_5_4_io_outs_up[24] ,
    \ces_5_4_io_outs_up[23] ,
    \ces_5_4_io_outs_up[22] ,
    \ces_5_4_io_outs_up[21] ,
    \ces_5_4_io_outs_up[20] ,
    \ces_5_4_io_outs_up[19] ,
    \ces_5_4_io_outs_up[18] ,
    \ces_5_4_io_outs_up[17] ,
    \ces_5_4_io_outs_up[16] ,
    \ces_5_4_io_outs_up[15] ,
    \ces_5_4_io_outs_up[14] ,
    \ces_5_4_io_outs_up[13] ,
    \ces_5_4_io_outs_up[12] ,
    \ces_5_4_io_outs_up[11] ,
    \ces_5_4_io_outs_up[10] ,
    \ces_5_4_io_outs_up[9] ,
    \ces_5_4_io_outs_up[8] ,
    \ces_5_4_io_outs_up[7] ,
    \ces_5_4_io_outs_up[6] ,
    \ces_5_4_io_outs_up[5] ,
    \ces_5_4_io_outs_up[4] ,
    \ces_5_4_io_outs_up[3] ,
    \ces_5_4_io_outs_up[2] ,
    \ces_5_4_io_outs_up[1] ,
    \ces_5_4_io_outs_up[0] }));
 Element ces_5_5 (.clock(clknet_3_6_0_clock),
    .io_lsbIns_1(ces_5_4_io_lsbOuts_1),
    .io_lsbIns_2(ces_5_4_io_lsbOuts_2),
    .io_lsbIns_3(ces_5_4_io_lsbOuts_3),
    .io_lsbIns_4(ces_5_4_io_lsbOuts_4),
    .io_lsbIns_5(ces_5_4_io_lsbOuts_5),
    .io_lsbIns_6(ces_5_4_io_lsbOuts_6),
    .io_lsbIns_7(ces_5_4_io_lsbOuts_7),
    .io_lsbOuts_0(ces_5_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_5_io_lsbOuts_7),
    .io_ins_down({\ces_5_5_io_ins_down[63] ,
    \ces_5_5_io_ins_down[62] ,
    \ces_5_5_io_ins_down[61] ,
    \ces_5_5_io_ins_down[60] ,
    \ces_5_5_io_ins_down[59] ,
    \ces_5_5_io_ins_down[58] ,
    \ces_5_5_io_ins_down[57] ,
    \ces_5_5_io_ins_down[56] ,
    \ces_5_5_io_ins_down[55] ,
    \ces_5_5_io_ins_down[54] ,
    \ces_5_5_io_ins_down[53] ,
    \ces_5_5_io_ins_down[52] ,
    \ces_5_5_io_ins_down[51] ,
    \ces_5_5_io_ins_down[50] ,
    \ces_5_5_io_ins_down[49] ,
    \ces_5_5_io_ins_down[48] ,
    \ces_5_5_io_ins_down[47] ,
    \ces_5_5_io_ins_down[46] ,
    \ces_5_5_io_ins_down[45] ,
    \ces_5_5_io_ins_down[44] ,
    \ces_5_5_io_ins_down[43] ,
    \ces_5_5_io_ins_down[42] ,
    \ces_5_5_io_ins_down[41] ,
    \ces_5_5_io_ins_down[40] ,
    \ces_5_5_io_ins_down[39] ,
    \ces_5_5_io_ins_down[38] ,
    \ces_5_5_io_ins_down[37] ,
    \ces_5_5_io_ins_down[36] ,
    \ces_5_5_io_ins_down[35] ,
    \ces_5_5_io_ins_down[34] ,
    \ces_5_5_io_ins_down[33] ,
    \ces_5_5_io_ins_down[32] ,
    \ces_5_5_io_ins_down[31] ,
    \ces_5_5_io_ins_down[30] ,
    \ces_5_5_io_ins_down[29] ,
    \ces_5_5_io_ins_down[28] ,
    \ces_5_5_io_ins_down[27] ,
    \ces_5_5_io_ins_down[26] ,
    \ces_5_5_io_ins_down[25] ,
    \ces_5_5_io_ins_down[24] ,
    \ces_5_5_io_ins_down[23] ,
    \ces_5_5_io_ins_down[22] ,
    \ces_5_5_io_ins_down[21] ,
    \ces_5_5_io_ins_down[20] ,
    \ces_5_5_io_ins_down[19] ,
    \ces_5_5_io_ins_down[18] ,
    \ces_5_5_io_ins_down[17] ,
    \ces_5_5_io_ins_down[16] ,
    \ces_5_5_io_ins_down[15] ,
    \ces_5_5_io_ins_down[14] ,
    \ces_5_5_io_ins_down[13] ,
    \ces_5_5_io_ins_down[12] ,
    \ces_5_5_io_ins_down[11] ,
    \ces_5_5_io_ins_down[10] ,
    \ces_5_5_io_ins_down[9] ,
    \ces_5_5_io_ins_down[8] ,
    \ces_5_5_io_ins_down[7] ,
    \ces_5_5_io_ins_down[6] ,
    \ces_5_5_io_ins_down[5] ,
    \ces_5_5_io_ins_down[4] ,
    \ces_5_5_io_ins_down[3] ,
    \ces_5_5_io_ins_down[2] ,
    \ces_5_5_io_ins_down[1] ,
    \ces_5_5_io_ins_down[0] }),
    .io_ins_left({\ces_5_5_io_ins_left[63] ,
    \ces_5_5_io_ins_left[62] ,
    \ces_5_5_io_ins_left[61] ,
    \ces_5_5_io_ins_left[60] ,
    \ces_5_5_io_ins_left[59] ,
    \ces_5_5_io_ins_left[58] ,
    \ces_5_5_io_ins_left[57] ,
    \ces_5_5_io_ins_left[56] ,
    \ces_5_5_io_ins_left[55] ,
    \ces_5_5_io_ins_left[54] ,
    \ces_5_5_io_ins_left[53] ,
    \ces_5_5_io_ins_left[52] ,
    \ces_5_5_io_ins_left[51] ,
    \ces_5_5_io_ins_left[50] ,
    \ces_5_5_io_ins_left[49] ,
    \ces_5_5_io_ins_left[48] ,
    \ces_5_5_io_ins_left[47] ,
    \ces_5_5_io_ins_left[46] ,
    \ces_5_5_io_ins_left[45] ,
    \ces_5_5_io_ins_left[44] ,
    \ces_5_5_io_ins_left[43] ,
    \ces_5_5_io_ins_left[42] ,
    \ces_5_5_io_ins_left[41] ,
    \ces_5_5_io_ins_left[40] ,
    \ces_5_5_io_ins_left[39] ,
    \ces_5_5_io_ins_left[38] ,
    \ces_5_5_io_ins_left[37] ,
    \ces_5_5_io_ins_left[36] ,
    \ces_5_5_io_ins_left[35] ,
    \ces_5_5_io_ins_left[34] ,
    \ces_5_5_io_ins_left[33] ,
    \ces_5_5_io_ins_left[32] ,
    \ces_5_5_io_ins_left[31] ,
    \ces_5_5_io_ins_left[30] ,
    \ces_5_5_io_ins_left[29] ,
    \ces_5_5_io_ins_left[28] ,
    \ces_5_5_io_ins_left[27] ,
    \ces_5_5_io_ins_left[26] ,
    \ces_5_5_io_ins_left[25] ,
    \ces_5_5_io_ins_left[24] ,
    \ces_5_5_io_ins_left[23] ,
    \ces_5_5_io_ins_left[22] ,
    \ces_5_5_io_ins_left[21] ,
    \ces_5_5_io_ins_left[20] ,
    \ces_5_5_io_ins_left[19] ,
    \ces_5_5_io_ins_left[18] ,
    \ces_5_5_io_ins_left[17] ,
    \ces_5_5_io_ins_left[16] ,
    \ces_5_5_io_ins_left[15] ,
    \ces_5_5_io_ins_left[14] ,
    \ces_5_5_io_ins_left[13] ,
    \ces_5_5_io_ins_left[12] ,
    \ces_5_5_io_ins_left[11] ,
    \ces_5_5_io_ins_left[10] ,
    \ces_5_5_io_ins_left[9] ,
    \ces_5_5_io_ins_left[8] ,
    \ces_5_5_io_ins_left[7] ,
    \ces_5_5_io_ins_left[6] ,
    \ces_5_5_io_ins_left[5] ,
    \ces_5_5_io_ins_left[4] ,
    \ces_5_5_io_ins_left[3] ,
    \ces_5_5_io_ins_left[2] ,
    \ces_5_5_io_ins_left[1] ,
    \ces_5_5_io_ins_left[0] }),
    .io_ins_right({\ces_5_4_io_outs_right[63] ,
    \ces_5_4_io_outs_right[62] ,
    \ces_5_4_io_outs_right[61] ,
    \ces_5_4_io_outs_right[60] ,
    \ces_5_4_io_outs_right[59] ,
    \ces_5_4_io_outs_right[58] ,
    \ces_5_4_io_outs_right[57] ,
    \ces_5_4_io_outs_right[56] ,
    \ces_5_4_io_outs_right[55] ,
    \ces_5_4_io_outs_right[54] ,
    \ces_5_4_io_outs_right[53] ,
    \ces_5_4_io_outs_right[52] ,
    \ces_5_4_io_outs_right[51] ,
    \ces_5_4_io_outs_right[50] ,
    \ces_5_4_io_outs_right[49] ,
    \ces_5_4_io_outs_right[48] ,
    \ces_5_4_io_outs_right[47] ,
    \ces_5_4_io_outs_right[46] ,
    \ces_5_4_io_outs_right[45] ,
    \ces_5_4_io_outs_right[44] ,
    \ces_5_4_io_outs_right[43] ,
    \ces_5_4_io_outs_right[42] ,
    \ces_5_4_io_outs_right[41] ,
    \ces_5_4_io_outs_right[40] ,
    \ces_5_4_io_outs_right[39] ,
    \ces_5_4_io_outs_right[38] ,
    \ces_5_4_io_outs_right[37] ,
    \ces_5_4_io_outs_right[36] ,
    \ces_5_4_io_outs_right[35] ,
    \ces_5_4_io_outs_right[34] ,
    \ces_5_4_io_outs_right[33] ,
    \ces_5_4_io_outs_right[32] ,
    \ces_5_4_io_outs_right[31] ,
    \ces_5_4_io_outs_right[30] ,
    \ces_5_4_io_outs_right[29] ,
    \ces_5_4_io_outs_right[28] ,
    \ces_5_4_io_outs_right[27] ,
    \ces_5_4_io_outs_right[26] ,
    \ces_5_4_io_outs_right[25] ,
    \ces_5_4_io_outs_right[24] ,
    \ces_5_4_io_outs_right[23] ,
    \ces_5_4_io_outs_right[22] ,
    \ces_5_4_io_outs_right[21] ,
    \ces_5_4_io_outs_right[20] ,
    \ces_5_4_io_outs_right[19] ,
    \ces_5_4_io_outs_right[18] ,
    \ces_5_4_io_outs_right[17] ,
    \ces_5_4_io_outs_right[16] ,
    \ces_5_4_io_outs_right[15] ,
    \ces_5_4_io_outs_right[14] ,
    \ces_5_4_io_outs_right[13] ,
    \ces_5_4_io_outs_right[12] ,
    \ces_5_4_io_outs_right[11] ,
    \ces_5_4_io_outs_right[10] ,
    \ces_5_4_io_outs_right[9] ,
    \ces_5_4_io_outs_right[8] ,
    \ces_5_4_io_outs_right[7] ,
    \ces_5_4_io_outs_right[6] ,
    \ces_5_4_io_outs_right[5] ,
    \ces_5_4_io_outs_right[4] ,
    \ces_5_4_io_outs_right[3] ,
    \ces_5_4_io_outs_right[2] ,
    \ces_5_4_io_outs_right[1] ,
    \ces_5_4_io_outs_right[0] }),
    .io_ins_up({\ces_4_5_io_outs_up[63] ,
    \ces_4_5_io_outs_up[62] ,
    \ces_4_5_io_outs_up[61] ,
    \ces_4_5_io_outs_up[60] ,
    \ces_4_5_io_outs_up[59] ,
    \ces_4_5_io_outs_up[58] ,
    \ces_4_5_io_outs_up[57] ,
    \ces_4_5_io_outs_up[56] ,
    \ces_4_5_io_outs_up[55] ,
    \ces_4_5_io_outs_up[54] ,
    \ces_4_5_io_outs_up[53] ,
    \ces_4_5_io_outs_up[52] ,
    \ces_4_5_io_outs_up[51] ,
    \ces_4_5_io_outs_up[50] ,
    \ces_4_5_io_outs_up[49] ,
    \ces_4_5_io_outs_up[48] ,
    \ces_4_5_io_outs_up[47] ,
    \ces_4_5_io_outs_up[46] ,
    \ces_4_5_io_outs_up[45] ,
    \ces_4_5_io_outs_up[44] ,
    \ces_4_5_io_outs_up[43] ,
    \ces_4_5_io_outs_up[42] ,
    \ces_4_5_io_outs_up[41] ,
    \ces_4_5_io_outs_up[40] ,
    \ces_4_5_io_outs_up[39] ,
    \ces_4_5_io_outs_up[38] ,
    \ces_4_5_io_outs_up[37] ,
    \ces_4_5_io_outs_up[36] ,
    \ces_4_5_io_outs_up[35] ,
    \ces_4_5_io_outs_up[34] ,
    \ces_4_5_io_outs_up[33] ,
    \ces_4_5_io_outs_up[32] ,
    \ces_4_5_io_outs_up[31] ,
    \ces_4_5_io_outs_up[30] ,
    \ces_4_5_io_outs_up[29] ,
    \ces_4_5_io_outs_up[28] ,
    \ces_4_5_io_outs_up[27] ,
    \ces_4_5_io_outs_up[26] ,
    \ces_4_5_io_outs_up[25] ,
    \ces_4_5_io_outs_up[24] ,
    \ces_4_5_io_outs_up[23] ,
    \ces_4_5_io_outs_up[22] ,
    \ces_4_5_io_outs_up[21] ,
    \ces_4_5_io_outs_up[20] ,
    \ces_4_5_io_outs_up[19] ,
    \ces_4_5_io_outs_up[18] ,
    \ces_4_5_io_outs_up[17] ,
    \ces_4_5_io_outs_up[16] ,
    \ces_4_5_io_outs_up[15] ,
    \ces_4_5_io_outs_up[14] ,
    \ces_4_5_io_outs_up[13] ,
    \ces_4_5_io_outs_up[12] ,
    \ces_4_5_io_outs_up[11] ,
    \ces_4_5_io_outs_up[10] ,
    \ces_4_5_io_outs_up[9] ,
    \ces_4_5_io_outs_up[8] ,
    \ces_4_5_io_outs_up[7] ,
    \ces_4_5_io_outs_up[6] ,
    \ces_4_5_io_outs_up[5] ,
    \ces_4_5_io_outs_up[4] ,
    \ces_4_5_io_outs_up[3] ,
    \ces_4_5_io_outs_up[2] ,
    \ces_4_5_io_outs_up[1] ,
    \ces_4_5_io_outs_up[0] }),
    .io_outs_down({\ces_4_5_io_ins_down[63] ,
    \ces_4_5_io_ins_down[62] ,
    \ces_4_5_io_ins_down[61] ,
    \ces_4_5_io_ins_down[60] ,
    \ces_4_5_io_ins_down[59] ,
    \ces_4_5_io_ins_down[58] ,
    \ces_4_5_io_ins_down[57] ,
    \ces_4_5_io_ins_down[56] ,
    \ces_4_5_io_ins_down[55] ,
    \ces_4_5_io_ins_down[54] ,
    \ces_4_5_io_ins_down[53] ,
    \ces_4_5_io_ins_down[52] ,
    \ces_4_5_io_ins_down[51] ,
    \ces_4_5_io_ins_down[50] ,
    \ces_4_5_io_ins_down[49] ,
    \ces_4_5_io_ins_down[48] ,
    \ces_4_5_io_ins_down[47] ,
    \ces_4_5_io_ins_down[46] ,
    \ces_4_5_io_ins_down[45] ,
    \ces_4_5_io_ins_down[44] ,
    \ces_4_5_io_ins_down[43] ,
    \ces_4_5_io_ins_down[42] ,
    \ces_4_5_io_ins_down[41] ,
    \ces_4_5_io_ins_down[40] ,
    \ces_4_5_io_ins_down[39] ,
    \ces_4_5_io_ins_down[38] ,
    \ces_4_5_io_ins_down[37] ,
    \ces_4_5_io_ins_down[36] ,
    \ces_4_5_io_ins_down[35] ,
    \ces_4_5_io_ins_down[34] ,
    \ces_4_5_io_ins_down[33] ,
    \ces_4_5_io_ins_down[32] ,
    \ces_4_5_io_ins_down[31] ,
    \ces_4_5_io_ins_down[30] ,
    \ces_4_5_io_ins_down[29] ,
    \ces_4_5_io_ins_down[28] ,
    \ces_4_5_io_ins_down[27] ,
    \ces_4_5_io_ins_down[26] ,
    \ces_4_5_io_ins_down[25] ,
    \ces_4_5_io_ins_down[24] ,
    \ces_4_5_io_ins_down[23] ,
    \ces_4_5_io_ins_down[22] ,
    \ces_4_5_io_ins_down[21] ,
    \ces_4_5_io_ins_down[20] ,
    \ces_4_5_io_ins_down[19] ,
    \ces_4_5_io_ins_down[18] ,
    \ces_4_5_io_ins_down[17] ,
    \ces_4_5_io_ins_down[16] ,
    \ces_4_5_io_ins_down[15] ,
    \ces_4_5_io_ins_down[14] ,
    \ces_4_5_io_ins_down[13] ,
    \ces_4_5_io_ins_down[12] ,
    \ces_4_5_io_ins_down[11] ,
    \ces_4_5_io_ins_down[10] ,
    \ces_4_5_io_ins_down[9] ,
    \ces_4_5_io_ins_down[8] ,
    \ces_4_5_io_ins_down[7] ,
    \ces_4_5_io_ins_down[6] ,
    \ces_4_5_io_ins_down[5] ,
    \ces_4_5_io_ins_down[4] ,
    \ces_4_5_io_ins_down[3] ,
    \ces_4_5_io_ins_down[2] ,
    \ces_4_5_io_ins_down[1] ,
    \ces_4_5_io_ins_down[0] }),
    .io_outs_left({\ces_5_4_io_ins_left[63] ,
    \ces_5_4_io_ins_left[62] ,
    \ces_5_4_io_ins_left[61] ,
    \ces_5_4_io_ins_left[60] ,
    \ces_5_4_io_ins_left[59] ,
    \ces_5_4_io_ins_left[58] ,
    \ces_5_4_io_ins_left[57] ,
    \ces_5_4_io_ins_left[56] ,
    \ces_5_4_io_ins_left[55] ,
    \ces_5_4_io_ins_left[54] ,
    \ces_5_4_io_ins_left[53] ,
    \ces_5_4_io_ins_left[52] ,
    \ces_5_4_io_ins_left[51] ,
    \ces_5_4_io_ins_left[50] ,
    \ces_5_4_io_ins_left[49] ,
    \ces_5_4_io_ins_left[48] ,
    \ces_5_4_io_ins_left[47] ,
    \ces_5_4_io_ins_left[46] ,
    \ces_5_4_io_ins_left[45] ,
    \ces_5_4_io_ins_left[44] ,
    \ces_5_4_io_ins_left[43] ,
    \ces_5_4_io_ins_left[42] ,
    \ces_5_4_io_ins_left[41] ,
    \ces_5_4_io_ins_left[40] ,
    \ces_5_4_io_ins_left[39] ,
    \ces_5_4_io_ins_left[38] ,
    \ces_5_4_io_ins_left[37] ,
    \ces_5_4_io_ins_left[36] ,
    \ces_5_4_io_ins_left[35] ,
    \ces_5_4_io_ins_left[34] ,
    \ces_5_4_io_ins_left[33] ,
    \ces_5_4_io_ins_left[32] ,
    \ces_5_4_io_ins_left[31] ,
    \ces_5_4_io_ins_left[30] ,
    \ces_5_4_io_ins_left[29] ,
    \ces_5_4_io_ins_left[28] ,
    \ces_5_4_io_ins_left[27] ,
    \ces_5_4_io_ins_left[26] ,
    \ces_5_4_io_ins_left[25] ,
    \ces_5_4_io_ins_left[24] ,
    \ces_5_4_io_ins_left[23] ,
    \ces_5_4_io_ins_left[22] ,
    \ces_5_4_io_ins_left[21] ,
    \ces_5_4_io_ins_left[20] ,
    \ces_5_4_io_ins_left[19] ,
    \ces_5_4_io_ins_left[18] ,
    \ces_5_4_io_ins_left[17] ,
    \ces_5_4_io_ins_left[16] ,
    \ces_5_4_io_ins_left[15] ,
    \ces_5_4_io_ins_left[14] ,
    \ces_5_4_io_ins_left[13] ,
    \ces_5_4_io_ins_left[12] ,
    \ces_5_4_io_ins_left[11] ,
    \ces_5_4_io_ins_left[10] ,
    \ces_5_4_io_ins_left[9] ,
    \ces_5_4_io_ins_left[8] ,
    \ces_5_4_io_ins_left[7] ,
    \ces_5_4_io_ins_left[6] ,
    \ces_5_4_io_ins_left[5] ,
    \ces_5_4_io_ins_left[4] ,
    \ces_5_4_io_ins_left[3] ,
    \ces_5_4_io_ins_left[2] ,
    \ces_5_4_io_ins_left[1] ,
    \ces_5_4_io_ins_left[0] }),
    .io_outs_right({\ces_5_5_io_outs_right[63] ,
    \ces_5_5_io_outs_right[62] ,
    \ces_5_5_io_outs_right[61] ,
    \ces_5_5_io_outs_right[60] ,
    \ces_5_5_io_outs_right[59] ,
    \ces_5_5_io_outs_right[58] ,
    \ces_5_5_io_outs_right[57] ,
    \ces_5_5_io_outs_right[56] ,
    \ces_5_5_io_outs_right[55] ,
    \ces_5_5_io_outs_right[54] ,
    \ces_5_5_io_outs_right[53] ,
    \ces_5_5_io_outs_right[52] ,
    \ces_5_5_io_outs_right[51] ,
    \ces_5_5_io_outs_right[50] ,
    \ces_5_5_io_outs_right[49] ,
    \ces_5_5_io_outs_right[48] ,
    \ces_5_5_io_outs_right[47] ,
    \ces_5_5_io_outs_right[46] ,
    \ces_5_5_io_outs_right[45] ,
    \ces_5_5_io_outs_right[44] ,
    \ces_5_5_io_outs_right[43] ,
    \ces_5_5_io_outs_right[42] ,
    \ces_5_5_io_outs_right[41] ,
    \ces_5_5_io_outs_right[40] ,
    \ces_5_5_io_outs_right[39] ,
    \ces_5_5_io_outs_right[38] ,
    \ces_5_5_io_outs_right[37] ,
    \ces_5_5_io_outs_right[36] ,
    \ces_5_5_io_outs_right[35] ,
    \ces_5_5_io_outs_right[34] ,
    \ces_5_5_io_outs_right[33] ,
    \ces_5_5_io_outs_right[32] ,
    \ces_5_5_io_outs_right[31] ,
    \ces_5_5_io_outs_right[30] ,
    \ces_5_5_io_outs_right[29] ,
    \ces_5_5_io_outs_right[28] ,
    \ces_5_5_io_outs_right[27] ,
    \ces_5_5_io_outs_right[26] ,
    \ces_5_5_io_outs_right[25] ,
    \ces_5_5_io_outs_right[24] ,
    \ces_5_5_io_outs_right[23] ,
    \ces_5_5_io_outs_right[22] ,
    \ces_5_5_io_outs_right[21] ,
    \ces_5_5_io_outs_right[20] ,
    \ces_5_5_io_outs_right[19] ,
    \ces_5_5_io_outs_right[18] ,
    \ces_5_5_io_outs_right[17] ,
    \ces_5_5_io_outs_right[16] ,
    \ces_5_5_io_outs_right[15] ,
    \ces_5_5_io_outs_right[14] ,
    \ces_5_5_io_outs_right[13] ,
    \ces_5_5_io_outs_right[12] ,
    \ces_5_5_io_outs_right[11] ,
    \ces_5_5_io_outs_right[10] ,
    \ces_5_5_io_outs_right[9] ,
    \ces_5_5_io_outs_right[8] ,
    \ces_5_5_io_outs_right[7] ,
    \ces_5_5_io_outs_right[6] ,
    \ces_5_5_io_outs_right[5] ,
    \ces_5_5_io_outs_right[4] ,
    \ces_5_5_io_outs_right[3] ,
    \ces_5_5_io_outs_right[2] ,
    \ces_5_5_io_outs_right[1] ,
    \ces_5_5_io_outs_right[0] }),
    .io_outs_up({\ces_5_5_io_outs_up[63] ,
    \ces_5_5_io_outs_up[62] ,
    \ces_5_5_io_outs_up[61] ,
    \ces_5_5_io_outs_up[60] ,
    \ces_5_5_io_outs_up[59] ,
    \ces_5_5_io_outs_up[58] ,
    \ces_5_5_io_outs_up[57] ,
    \ces_5_5_io_outs_up[56] ,
    \ces_5_5_io_outs_up[55] ,
    \ces_5_5_io_outs_up[54] ,
    \ces_5_5_io_outs_up[53] ,
    \ces_5_5_io_outs_up[52] ,
    \ces_5_5_io_outs_up[51] ,
    \ces_5_5_io_outs_up[50] ,
    \ces_5_5_io_outs_up[49] ,
    \ces_5_5_io_outs_up[48] ,
    \ces_5_5_io_outs_up[47] ,
    \ces_5_5_io_outs_up[46] ,
    \ces_5_5_io_outs_up[45] ,
    \ces_5_5_io_outs_up[44] ,
    \ces_5_5_io_outs_up[43] ,
    \ces_5_5_io_outs_up[42] ,
    \ces_5_5_io_outs_up[41] ,
    \ces_5_5_io_outs_up[40] ,
    \ces_5_5_io_outs_up[39] ,
    \ces_5_5_io_outs_up[38] ,
    \ces_5_5_io_outs_up[37] ,
    \ces_5_5_io_outs_up[36] ,
    \ces_5_5_io_outs_up[35] ,
    \ces_5_5_io_outs_up[34] ,
    \ces_5_5_io_outs_up[33] ,
    \ces_5_5_io_outs_up[32] ,
    \ces_5_5_io_outs_up[31] ,
    \ces_5_5_io_outs_up[30] ,
    \ces_5_5_io_outs_up[29] ,
    \ces_5_5_io_outs_up[28] ,
    \ces_5_5_io_outs_up[27] ,
    \ces_5_5_io_outs_up[26] ,
    \ces_5_5_io_outs_up[25] ,
    \ces_5_5_io_outs_up[24] ,
    \ces_5_5_io_outs_up[23] ,
    \ces_5_5_io_outs_up[22] ,
    \ces_5_5_io_outs_up[21] ,
    \ces_5_5_io_outs_up[20] ,
    \ces_5_5_io_outs_up[19] ,
    \ces_5_5_io_outs_up[18] ,
    \ces_5_5_io_outs_up[17] ,
    \ces_5_5_io_outs_up[16] ,
    \ces_5_5_io_outs_up[15] ,
    \ces_5_5_io_outs_up[14] ,
    \ces_5_5_io_outs_up[13] ,
    \ces_5_5_io_outs_up[12] ,
    \ces_5_5_io_outs_up[11] ,
    \ces_5_5_io_outs_up[10] ,
    \ces_5_5_io_outs_up[9] ,
    \ces_5_5_io_outs_up[8] ,
    \ces_5_5_io_outs_up[7] ,
    \ces_5_5_io_outs_up[6] ,
    \ces_5_5_io_outs_up[5] ,
    \ces_5_5_io_outs_up[4] ,
    \ces_5_5_io_outs_up[3] ,
    \ces_5_5_io_outs_up[2] ,
    \ces_5_5_io_outs_up[1] ,
    \ces_5_5_io_outs_up[0] }));
 Element ces_5_6 (.clock(clknet_3_6_0_clock),
    .io_lsbIns_1(ces_5_5_io_lsbOuts_1),
    .io_lsbIns_2(ces_5_5_io_lsbOuts_2),
    .io_lsbIns_3(ces_5_5_io_lsbOuts_3),
    .io_lsbIns_4(ces_5_5_io_lsbOuts_4),
    .io_lsbIns_5(ces_5_5_io_lsbOuts_5),
    .io_lsbIns_6(ces_5_5_io_lsbOuts_6),
    .io_lsbIns_7(ces_5_5_io_lsbOuts_7),
    .io_lsbOuts_0(ces_5_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_6_io_lsbOuts_7),
    .io_ins_down({\ces_5_6_io_ins_down[63] ,
    \ces_5_6_io_ins_down[62] ,
    \ces_5_6_io_ins_down[61] ,
    \ces_5_6_io_ins_down[60] ,
    \ces_5_6_io_ins_down[59] ,
    \ces_5_6_io_ins_down[58] ,
    \ces_5_6_io_ins_down[57] ,
    \ces_5_6_io_ins_down[56] ,
    \ces_5_6_io_ins_down[55] ,
    \ces_5_6_io_ins_down[54] ,
    \ces_5_6_io_ins_down[53] ,
    \ces_5_6_io_ins_down[52] ,
    \ces_5_6_io_ins_down[51] ,
    \ces_5_6_io_ins_down[50] ,
    \ces_5_6_io_ins_down[49] ,
    \ces_5_6_io_ins_down[48] ,
    \ces_5_6_io_ins_down[47] ,
    \ces_5_6_io_ins_down[46] ,
    \ces_5_6_io_ins_down[45] ,
    \ces_5_6_io_ins_down[44] ,
    \ces_5_6_io_ins_down[43] ,
    \ces_5_6_io_ins_down[42] ,
    \ces_5_6_io_ins_down[41] ,
    \ces_5_6_io_ins_down[40] ,
    \ces_5_6_io_ins_down[39] ,
    \ces_5_6_io_ins_down[38] ,
    \ces_5_6_io_ins_down[37] ,
    \ces_5_6_io_ins_down[36] ,
    \ces_5_6_io_ins_down[35] ,
    \ces_5_6_io_ins_down[34] ,
    \ces_5_6_io_ins_down[33] ,
    \ces_5_6_io_ins_down[32] ,
    \ces_5_6_io_ins_down[31] ,
    \ces_5_6_io_ins_down[30] ,
    \ces_5_6_io_ins_down[29] ,
    \ces_5_6_io_ins_down[28] ,
    \ces_5_6_io_ins_down[27] ,
    \ces_5_6_io_ins_down[26] ,
    \ces_5_6_io_ins_down[25] ,
    \ces_5_6_io_ins_down[24] ,
    \ces_5_6_io_ins_down[23] ,
    \ces_5_6_io_ins_down[22] ,
    \ces_5_6_io_ins_down[21] ,
    \ces_5_6_io_ins_down[20] ,
    \ces_5_6_io_ins_down[19] ,
    \ces_5_6_io_ins_down[18] ,
    \ces_5_6_io_ins_down[17] ,
    \ces_5_6_io_ins_down[16] ,
    \ces_5_6_io_ins_down[15] ,
    \ces_5_6_io_ins_down[14] ,
    \ces_5_6_io_ins_down[13] ,
    \ces_5_6_io_ins_down[12] ,
    \ces_5_6_io_ins_down[11] ,
    \ces_5_6_io_ins_down[10] ,
    \ces_5_6_io_ins_down[9] ,
    \ces_5_6_io_ins_down[8] ,
    \ces_5_6_io_ins_down[7] ,
    \ces_5_6_io_ins_down[6] ,
    \ces_5_6_io_ins_down[5] ,
    \ces_5_6_io_ins_down[4] ,
    \ces_5_6_io_ins_down[3] ,
    \ces_5_6_io_ins_down[2] ,
    \ces_5_6_io_ins_down[1] ,
    \ces_5_6_io_ins_down[0] }),
    .io_ins_left({\ces_5_6_io_ins_left[63] ,
    \ces_5_6_io_ins_left[62] ,
    \ces_5_6_io_ins_left[61] ,
    \ces_5_6_io_ins_left[60] ,
    \ces_5_6_io_ins_left[59] ,
    \ces_5_6_io_ins_left[58] ,
    \ces_5_6_io_ins_left[57] ,
    \ces_5_6_io_ins_left[56] ,
    \ces_5_6_io_ins_left[55] ,
    \ces_5_6_io_ins_left[54] ,
    \ces_5_6_io_ins_left[53] ,
    \ces_5_6_io_ins_left[52] ,
    \ces_5_6_io_ins_left[51] ,
    \ces_5_6_io_ins_left[50] ,
    \ces_5_6_io_ins_left[49] ,
    \ces_5_6_io_ins_left[48] ,
    \ces_5_6_io_ins_left[47] ,
    \ces_5_6_io_ins_left[46] ,
    \ces_5_6_io_ins_left[45] ,
    \ces_5_6_io_ins_left[44] ,
    \ces_5_6_io_ins_left[43] ,
    \ces_5_6_io_ins_left[42] ,
    \ces_5_6_io_ins_left[41] ,
    \ces_5_6_io_ins_left[40] ,
    \ces_5_6_io_ins_left[39] ,
    \ces_5_6_io_ins_left[38] ,
    \ces_5_6_io_ins_left[37] ,
    \ces_5_6_io_ins_left[36] ,
    \ces_5_6_io_ins_left[35] ,
    \ces_5_6_io_ins_left[34] ,
    \ces_5_6_io_ins_left[33] ,
    \ces_5_6_io_ins_left[32] ,
    \ces_5_6_io_ins_left[31] ,
    \ces_5_6_io_ins_left[30] ,
    \ces_5_6_io_ins_left[29] ,
    \ces_5_6_io_ins_left[28] ,
    \ces_5_6_io_ins_left[27] ,
    \ces_5_6_io_ins_left[26] ,
    \ces_5_6_io_ins_left[25] ,
    \ces_5_6_io_ins_left[24] ,
    \ces_5_6_io_ins_left[23] ,
    \ces_5_6_io_ins_left[22] ,
    \ces_5_6_io_ins_left[21] ,
    \ces_5_6_io_ins_left[20] ,
    \ces_5_6_io_ins_left[19] ,
    \ces_5_6_io_ins_left[18] ,
    \ces_5_6_io_ins_left[17] ,
    \ces_5_6_io_ins_left[16] ,
    \ces_5_6_io_ins_left[15] ,
    \ces_5_6_io_ins_left[14] ,
    \ces_5_6_io_ins_left[13] ,
    \ces_5_6_io_ins_left[12] ,
    \ces_5_6_io_ins_left[11] ,
    \ces_5_6_io_ins_left[10] ,
    \ces_5_6_io_ins_left[9] ,
    \ces_5_6_io_ins_left[8] ,
    \ces_5_6_io_ins_left[7] ,
    \ces_5_6_io_ins_left[6] ,
    \ces_5_6_io_ins_left[5] ,
    \ces_5_6_io_ins_left[4] ,
    \ces_5_6_io_ins_left[3] ,
    \ces_5_6_io_ins_left[2] ,
    \ces_5_6_io_ins_left[1] ,
    \ces_5_6_io_ins_left[0] }),
    .io_ins_right({\ces_5_5_io_outs_right[63] ,
    \ces_5_5_io_outs_right[62] ,
    \ces_5_5_io_outs_right[61] ,
    \ces_5_5_io_outs_right[60] ,
    \ces_5_5_io_outs_right[59] ,
    \ces_5_5_io_outs_right[58] ,
    \ces_5_5_io_outs_right[57] ,
    \ces_5_5_io_outs_right[56] ,
    \ces_5_5_io_outs_right[55] ,
    \ces_5_5_io_outs_right[54] ,
    \ces_5_5_io_outs_right[53] ,
    \ces_5_5_io_outs_right[52] ,
    \ces_5_5_io_outs_right[51] ,
    \ces_5_5_io_outs_right[50] ,
    \ces_5_5_io_outs_right[49] ,
    \ces_5_5_io_outs_right[48] ,
    \ces_5_5_io_outs_right[47] ,
    \ces_5_5_io_outs_right[46] ,
    \ces_5_5_io_outs_right[45] ,
    \ces_5_5_io_outs_right[44] ,
    \ces_5_5_io_outs_right[43] ,
    \ces_5_5_io_outs_right[42] ,
    \ces_5_5_io_outs_right[41] ,
    \ces_5_5_io_outs_right[40] ,
    \ces_5_5_io_outs_right[39] ,
    \ces_5_5_io_outs_right[38] ,
    \ces_5_5_io_outs_right[37] ,
    \ces_5_5_io_outs_right[36] ,
    \ces_5_5_io_outs_right[35] ,
    \ces_5_5_io_outs_right[34] ,
    \ces_5_5_io_outs_right[33] ,
    \ces_5_5_io_outs_right[32] ,
    \ces_5_5_io_outs_right[31] ,
    \ces_5_5_io_outs_right[30] ,
    \ces_5_5_io_outs_right[29] ,
    \ces_5_5_io_outs_right[28] ,
    \ces_5_5_io_outs_right[27] ,
    \ces_5_5_io_outs_right[26] ,
    \ces_5_5_io_outs_right[25] ,
    \ces_5_5_io_outs_right[24] ,
    \ces_5_5_io_outs_right[23] ,
    \ces_5_5_io_outs_right[22] ,
    \ces_5_5_io_outs_right[21] ,
    \ces_5_5_io_outs_right[20] ,
    \ces_5_5_io_outs_right[19] ,
    \ces_5_5_io_outs_right[18] ,
    \ces_5_5_io_outs_right[17] ,
    \ces_5_5_io_outs_right[16] ,
    \ces_5_5_io_outs_right[15] ,
    \ces_5_5_io_outs_right[14] ,
    \ces_5_5_io_outs_right[13] ,
    \ces_5_5_io_outs_right[12] ,
    \ces_5_5_io_outs_right[11] ,
    \ces_5_5_io_outs_right[10] ,
    \ces_5_5_io_outs_right[9] ,
    \ces_5_5_io_outs_right[8] ,
    \ces_5_5_io_outs_right[7] ,
    \ces_5_5_io_outs_right[6] ,
    \ces_5_5_io_outs_right[5] ,
    \ces_5_5_io_outs_right[4] ,
    \ces_5_5_io_outs_right[3] ,
    \ces_5_5_io_outs_right[2] ,
    \ces_5_5_io_outs_right[1] ,
    \ces_5_5_io_outs_right[0] }),
    .io_ins_up({\ces_4_6_io_outs_up[63] ,
    \ces_4_6_io_outs_up[62] ,
    \ces_4_6_io_outs_up[61] ,
    \ces_4_6_io_outs_up[60] ,
    \ces_4_6_io_outs_up[59] ,
    \ces_4_6_io_outs_up[58] ,
    \ces_4_6_io_outs_up[57] ,
    \ces_4_6_io_outs_up[56] ,
    \ces_4_6_io_outs_up[55] ,
    \ces_4_6_io_outs_up[54] ,
    \ces_4_6_io_outs_up[53] ,
    \ces_4_6_io_outs_up[52] ,
    \ces_4_6_io_outs_up[51] ,
    \ces_4_6_io_outs_up[50] ,
    \ces_4_6_io_outs_up[49] ,
    \ces_4_6_io_outs_up[48] ,
    \ces_4_6_io_outs_up[47] ,
    \ces_4_6_io_outs_up[46] ,
    \ces_4_6_io_outs_up[45] ,
    \ces_4_6_io_outs_up[44] ,
    \ces_4_6_io_outs_up[43] ,
    \ces_4_6_io_outs_up[42] ,
    \ces_4_6_io_outs_up[41] ,
    \ces_4_6_io_outs_up[40] ,
    \ces_4_6_io_outs_up[39] ,
    \ces_4_6_io_outs_up[38] ,
    \ces_4_6_io_outs_up[37] ,
    \ces_4_6_io_outs_up[36] ,
    \ces_4_6_io_outs_up[35] ,
    \ces_4_6_io_outs_up[34] ,
    \ces_4_6_io_outs_up[33] ,
    \ces_4_6_io_outs_up[32] ,
    \ces_4_6_io_outs_up[31] ,
    \ces_4_6_io_outs_up[30] ,
    \ces_4_6_io_outs_up[29] ,
    \ces_4_6_io_outs_up[28] ,
    \ces_4_6_io_outs_up[27] ,
    \ces_4_6_io_outs_up[26] ,
    \ces_4_6_io_outs_up[25] ,
    \ces_4_6_io_outs_up[24] ,
    \ces_4_6_io_outs_up[23] ,
    \ces_4_6_io_outs_up[22] ,
    \ces_4_6_io_outs_up[21] ,
    \ces_4_6_io_outs_up[20] ,
    \ces_4_6_io_outs_up[19] ,
    \ces_4_6_io_outs_up[18] ,
    \ces_4_6_io_outs_up[17] ,
    \ces_4_6_io_outs_up[16] ,
    \ces_4_6_io_outs_up[15] ,
    \ces_4_6_io_outs_up[14] ,
    \ces_4_6_io_outs_up[13] ,
    \ces_4_6_io_outs_up[12] ,
    \ces_4_6_io_outs_up[11] ,
    \ces_4_6_io_outs_up[10] ,
    \ces_4_6_io_outs_up[9] ,
    \ces_4_6_io_outs_up[8] ,
    \ces_4_6_io_outs_up[7] ,
    \ces_4_6_io_outs_up[6] ,
    \ces_4_6_io_outs_up[5] ,
    \ces_4_6_io_outs_up[4] ,
    \ces_4_6_io_outs_up[3] ,
    \ces_4_6_io_outs_up[2] ,
    \ces_4_6_io_outs_up[1] ,
    \ces_4_6_io_outs_up[0] }),
    .io_outs_down({\ces_4_6_io_ins_down[63] ,
    \ces_4_6_io_ins_down[62] ,
    \ces_4_6_io_ins_down[61] ,
    \ces_4_6_io_ins_down[60] ,
    \ces_4_6_io_ins_down[59] ,
    \ces_4_6_io_ins_down[58] ,
    \ces_4_6_io_ins_down[57] ,
    \ces_4_6_io_ins_down[56] ,
    \ces_4_6_io_ins_down[55] ,
    \ces_4_6_io_ins_down[54] ,
    \ces_4_6_io_ins_down[53] ,
    \ces_4_6_io_ins_down[52] ,
    \ces_4_6_io_ins_down[51] ,
    \ces_4_6_io_ins_down[50] ,
    \ces_4_6_io_ins_down[49] ,
    \ces_4_6_io_ins_down[48] ,
    \ces_4_6_io_ins_down[47] ,
    \ces_4_6_io_ins_down[46] ,
    \ces_4_6_io_ins_down[45] ,
    \ces_4_6_io_ins_down[44] ,
    \ces_4_6_io_ins_down[43] ,
    \ces_4_6_io_ins_down[42] ,
    \ces_4_6_io_ins_down[41] ,
    \ces_4_6_io_ins_down[40] ,
    \ces_4_6_io_ins_down[39] ,
    \ces_4_6_io_ins_down[38] ,
    \ces_4_6_io_ins_down[37] ,
    \ces_4_6_io_ins_down[36] ,
    \ces_4_6_io_ins_down[35] ,
    \ces_4_6_io_ins_down[34] ,
    \ces_4_6_io_ins_down[33] ,
    \ces_4_6_io_ins_down[32] ,
    \ces_4_6_io_ins_down[31] ,
    \ces_4_6_io_ins_down[30] ,
    \ces_4_6_io_ins_down[29] ,
    \ces_4_6_io_ins_down[28] ,
    \ces_4_6_io_ins_down[27] ,
    \ces_4_6_io_ins_down[26] ,
    \ces_4_6_io_ins_down[25] ,
    \ces_4_6_io_ins_down[24] ,
    \ces_4_6_io_ins_down[23] ,
    \ces_4_6_io_ins_down[22] ,
    \ces_4_6_io_ins_down[21] ,
    \ces_4_6_io_ins_down[20] ,
    \ces_4_6_io_ins_down[19] ,
    \ces_4_6_io_ins_down[18] ,
    \ces_4_6_io_ins_down[17] ,
    \ces_4_6_io_ins_down[16] ,
    \ces_4_6_io_ins_down[15] ,
    \ces_4_6_io_ins_down[14] ,
    \ces_4_6_io_ins_down[13] ,
    \ces_4_6_io_ins_down[12] ,
    \ces_4_6_io_ins_down[11] ,
    \ces_4_6_io_ins_down[10] ,
    \ces_4_6_io_ins_down[9] ,
    \ces_4_6_io_ins_down[8] ,
    \ces_4_6_io_ins_down[7] ,
    \ces_4_6_io_ins_down[6] ,
    \ces_4_6_io_ins_down[5] ,
    \ces_4_6_io_ins_down[4] ,
    \ces_4_6_io_ins_down[3] ,
    \ces_4_6_io_ins_down[2] ,
    \ces_4_6_io_ins_down[1] ,
    \ces_4_6_io_ins_down[0] }),
    .io_outs_left({\ces_5_5_io_ins_left[63] ,
    \ces_5_5_io_ins_left[62] ,
    \ces_5_5_io_ins_left[61] ,
    \ces_5_5_io_ins_left[60] ,
    \ces_5_5_io_ins_left[59] ,
    \ces_5_5_io_ins_left[58] ,
    \ces_5_5_io_ins_left[57] ,
    \ces_5_5_io_ins_left[56] ,
    \ces_5_5_io_ins_left[55] ,
    \ces_5_5_io_ins_left[54] ,
    \ces_5_5_io_ins_left[53] ,
    \ces_5_5_io_ins_left[52] ,
    \ces_5_5_io_ins_left[51] ,
    \ces_5_5_io_ins_left[50] ,
    \ces_5_5_io_ins_left[49] ,
    \ces_5_5_io_ins_left[48] ,
    \ces_5_5_io_ins_left[47] ,
    \ces_5_5_io_ins_left[46] ,
    \ces_5_5_io_ins_left[45] ,
    \ces_5_5_io_ins_left[44] ,
    \ces_5_5_io_ins_left[43] ,
    \ces_5_5_io_ins_left[42] ,
    \ces_5_5_io_ins_left[41] ,
    \ces_5_5_io_ins_left[40] ,
    \ces_5_5_io_ins_left[39] ,
    \ces_5_5_io_ins_left[38] ,
    \ces_5_5_io_ins_left[37] ,
    \ces_5_5_io_ins_left[36] ,
    \ces_5_5_io_ins_left[35] ,
    \ces_5_5_io_ins_left[34] ,
    \ces_5_5_io_ins_left[33] ,
    \ces_5_5_io_ins_left[32] ,
    \ces_5_5_io_ins_left[31] ,
    \ces_5_5_io_ins_left[30] ,
    \ces_5_5_io_ins_left[29] ,
    \ces_5_5_io_ins_left[28] ,
    \ces_5_5_io_ins_left[27] ,
    \ces_5_5_io_ins_left[26] ,
    \ces_5_5_io_ins_left[25] ,
    \ces_5_5_io_ins_left[24] ,
    \ces_5_5_io_ins_left[23] ,
    \ces_5_5_io_ins_left[22] ,
    \ces_5_5_io_ins_left[21] ,
    \ces_5_5_io_ins_left[20] ,
    \ces_5_5_io_ins_left[19] ,
    \ces_5_5_io_ins_left[18] ,
    \ces_5_5_io_ins_left[17] ,
    \ces_5_5_io_ins_left[16] ,
    \ces_5_5_io_ins_left[15] ,
    \ces_5_5_io_ins_left[14] ,
    \ces_5_5_io_ins_left[13] ,
    \ces_5_5_io_ins_left[12] ,
    \ces_5_5_io_ins_left[11] ,
    \ces_5_5_io_ins_left[10] ,
    \ces_5_5_io_ins_left[9] ,
    \ces_5_5_io_ins_left[8] ,
    \ces_5_5_io_ins_left[7] ,
    \ces_5_5_io_ins_left[6] ,
    \ces_5_5_io_ins_left[5] ,
    \ces_5_5_io_ins_left[4] ,
    \ces_5_5_io_ins_left[3] ,
    \ces_5_5_io_ins_left[2] ,
    \ces_5_5_io_ins_left[1] ,
    \ces_5_5_io_ins_left[0] }),
    .io_outs_right({\ces_5_6_io_outs_right[63] ,
    \ces_5_6_io_outs_right[62] ,
    \ces_5_6_io_outs_right[61] ,
    \ces_5_6_io_outs_right[60] ,
    \ces_5_6_io_outs_right[59] ,
    \ces_5_6_io_outs_right[58] ,
    \ces_5_6_io_outs_right[57] ,
    \ces_5_6_io_outs_right[56] ,
    \ces_5_6_io_outs_right[55] ,
    \ces_5_6_io_outs_right[54] ,
    \ces_5_6_io_outs_right[53] ,
    \ces_5_6_io_outs_right[52] ,
    \ces_5_6_io_outs_right[51] ,
    \ces_5_6_io_outs_right[50] ,
    \ces_5_6_io_outs_right[49] ,
    \ces_5_6_io_outs_right[48] ,
    \ces_5_6_io_outs_right[47] ,
    \ces_5_6_io_outs_right[46] ,
    \ces_5_6_io_outs_right[45] ,
    \ces_5_6_io_outs_right[44] ,
    \ces_5_6_io_outs_right[43] ,
    \ces_5_6_io_outs_right[42] ,
    \ces_5_6_io_outs_right[41] ,
    \ces_5_6_io_outs_right[40] ,
    \ces_5_6_io_outs_right[39] ,
    \ces_5_6_io_outs_right[38] ,
    \ces_5_6_io_outs_right[37] ,
    \ces_5_6_io_outs_right[36] ,
    \ces_5_6_io_outs_right[35] ,
    \ces_5_6_io_outs_right[34] ,
    \ces_5_6_io_outs_right[33] ,
    \ces_5_6_io_outs_right[32] ,
    \ces_5_6_io_outs_right[31] ,
    \ces_5_6_io_outs_right[30] ,
    \ces_5_6_io_outs_right[29] ,
    \ces_5_6_io_outs_right[28] ,
    \ces_5_6_io_outs_right[27] ,
    \ces_5_6_io_outs_right[26] ,
    \ces_5_6_io_outs_right[25] ,
    \ces_5_6_io_outs_right[24] ,
    \ces_5_6_io_outs_right[23] ,
    \ces_5_6_io_outs_right[22] ,
    \ces_5_6_io_outs_right[21] ,
    \ces_5_6_io_outs_right[20] ,
    \ces_5_6_io_outs_right[19] ,
    \ces_5_6_io_outs_right[18] ,
    \ces_5_6_io_outs_right[17] ,
    \ces_5_6_io_outs_right[16] ,
    \ces_5_6_io_outs_right[15] ,
    \ces_5_6_io_outs_right[14] ,
    \ces_5_6_io_outs_right[13] ,
    \ces_5_6_io_outs_right[12] ,
    \ces_5_6_io_outs_right[11] ,
    \ces_5_6_io_outs_right[10] ,
    \ces_5_6_io_outs_right[9] ,
    \ces_5_6_io_outs_right[8] ,
    \ces_5_6_io_outs_right[7] ,
    \ces_5_6_io_outs_right[6] ,
    \ces_5_6_io_outs_right[5] ,
    \ces_5_6_io_outs_right[4] ,
    \ces_5_6_io_outs_right[3] ,
    \ces_5_6_io_outs_right[2] ,
    \ces_5_6_io_outs_right[1] ,
    \ces_5_6_io_outs_right[0] }),
    .io_outs_up({\ces_5_6_io_outs_up[63] ,
    \ces_5_6_io_outs_up[62] ,
    \ces_5_6_io_outs_up[61] ,
    \ces_5_6_io_outs_up[60] ,
    \ces_5_6_io_outs_up[59] ,
    \ces_5_6_io_outs_up[58] ,
    \ces_5_6_io_outs_up[57] ,
    \ces_5_6_io_outs_up[56] ,
    \ces_5_6_io_outs_up[55] ,
    \ces_5_6_io_outs_up[54] ,
    \ces_5_6_io_outs_up[53] ,
    \ces_5_6_io_outs_up[52] ,
    \ces_5_6_io_outs_up[51] ,
    \ces_5_6_io_outs_up[50] ,
    \ces_5_6_io_outs_up[49] ,
    \ces_5_6_io_outs_up[48] ,
    \ces_5_6_io_outs_up[47] ,
    \ces_5_6_io_outs_up[46] ,
    \ces_5_6_io_outs_up[45] ,
    \ces_5_6_io_outs_up[44] ,
    \ces_5_6_io_outs_up[43] ,
    \ces_5_6_io_outs_up[42] ,
    \ces_5_6_io_outs_up[41] ,
    \ces_5_6_io_outs_up[40] ,
    \ces_5_6_io_outs_up[39] ,
    \ces_5_6_io_outs_up[38] ,
    \ces_5_6_io_outs_up[37] ,
    \ces_5_6_io_outs_up[36] ,
    \ces_5_6_io_outs_up[35] ,
    \ces_5_6_io_outs_up[34] ,
    \ces_5_6_io_outs_up[33] ,
    \ces_5_6_io_outs_up[32] ,
    \ces_5_6_io_outs_up[31] ,
    \ces_5_6_io_outs_up[30] ,
    \ces_5_6_io_outs_up[29] ,
    \ces_5_6_io_outs_up[28] ,
    \ces_5_6_io_outs_up[27] ,
    \ces_5_6_io_outs_up[26] ,
    \ces_5_6_io_outs_up[25] ,
    \ces_5_6_io_outs_up[24] ,
    \ces_5_6_io_outs_up[23] ,
    \ces_5_6_io_outs_up[22] ,
    \ces_5_6_io_outs_up[21] ,
    \ces_5_6_io_outs_up[20] ,
    \ces_5_6_io_outs_up[19] ,
    \ces_5_6_io_outs_up[18] ,
    \ces_5_6_io_outs_up[17] ,
    \ces_5_6_io_outs_up[16] ,
    \ces_5_6_io_outs_up[15] ,
    \ces_5_6_io_outs_up[14] ,
    \ces_5_6_io_outs_up[13] ,
    \ces_5_6_io_outs_up[12] ,
    \ces_5_6_io_outs_up[11] ,
    \ces_5_6_io_outs_up[10] ,
    \ces_5_6_io_outs_up[9] ,
    \ces_5_6_io_outs_up[8] ,
    \ces_5_6_io_outs_up[7] ,
    \ces_5_6_io_outs_up[6] ,
    \ces_5_6_io_outs_up[5] ,
    \ces_5_6_io_outs_up[4] ,
    \ces_5_6_io_outs_up[3] ,
    \ces_5_6_io_outs_up[2] ,
    \ces_5_6_io_outs_up[1] ,
    \ces_5_6_io_outs_up[0] }));
 Element ces_5_7 (.clock(clknet_3_6_0_clock),
    .io_lsbIns_1(ces_5_6_io_lsbOuts_1),
    .io_lsbIns_2(ces_5_6_io_lsbOuts_2),
    .io_lsbIns_3(ces_5_6_io_lsbOuts_3),
    .io_lsbIns_4(ces_5_6_io_lsbOuts_4),
    .io_lsbIns_5(ces_5_6_io_lsbOuts_5),
    .io_lsbIns_6(ces_5_6_io_lsbOuts_6),
    .io_lsbIns_7(ces_5_6_io_lsbOuts_7),
    .io_lsbOuts_0(ces_5_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_5_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_5_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_5_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_5_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_5_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_5_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_5_7_io_lsbOuts_7),
    .io_ins_down({\ces_5_7_io_ins_down[63] ,
    \ces_5_7_io_ins_down[62] ,
    \ces_5_7_io_ins_down[61] ,
    \ces_5_7_io_ins_down[60] ,
    \ces_5_7_io_ins_down[59] ,
    \ces_5_7_io_ins_down[58] ,
    \ces_5_7_io_ins_down[57] ,
    \ces_5_7_io_ins_down[56] ,
    \ces_5_7_io_ins_down[55] ,
    \ces_5_7_io_ins_down[54] ,
    \ces_5_7_io_ins_down[53] ,
    \ces_5_7_io_ins_down[52] ,
    \ces_5_7_io_ins_down[51] ,
    \ces_5_7_io_ins_down[50] ,
    \ces_5_7_io_ins_down[49] ,
    \ces_5_7_io_ins_down[48] ,
    \ces_5_7_io_ins_down[47] ,
    \ces_5_7_io_ins_down[46] ,
    \ces_5_7_io_ins_down[45] ,
    \ces_5_7_io_ins_down[44] ,
    \ces_5_7_io_ins_down[43] ,
    \ces_5_7_io_ins_down[42] ,
    \ces_5_7_io_ins_down[41] ,
    \ces_5_7_io_ins_down[40] ,
    \ces_5_7_io_ins_down[39] ,
    \ces_5_7_io_ins_down[38] ,
    \ces_5_7_io_ins_down[37] ,
    \ces_5_7_io_ins_down[36] ,
    \ces_5_7_io_ins_down[35] ,
    \ces_5_7_io_ins_down[34] ,
    \ces_5_7_io_ins_down[33] ,
    \ces_5_7_io_ins_down[32] ,
    \ces_5_7_io_ins_down[31] ,
    \ces_5_7_io_ins_down[30] ,
    \ces_5_7_io_ins_down[29] ,
    \ces_5_7_io_ins_down[28] ,
    \ces_5_7_io_ins_down[27] ,
    \ces_5_7_io_ins_down[26] ,
    \ces_5_7_io_ins_down[25] ,
    \ces_5_7_io_ins_down[24] ,
    \ces_5_7_io_ins_down[23] ,
    \ces_5_7_io_ins_down[22] ,
    \ces_5_7_io_ins_down[21] ,
    \ces_5_7_io_ins_down[20] ,
    \ces_5_7_io_ins_down[19] ,
    \ces_5_7_io_ins_down[18] ,
    \ces_5_7_io_ins_down[17] ,
    \ces_5_7_io_ins_down[16] ,
    \ces_5_7_io_ins_down[15] ,
    \ces_5_7_io_ins_down[14] ,
    \ces_5_7_io_ins_down[13] ,
    \ces_5_7_io_ins_down[12] ,
    \ces_5_7_io_ins_down[11] ,
    \ces_5_7_io_ins_down[10] ,
    \ces_5_7_io_ins_down[9] ,
    \ces_5_7_io_ins_down[8] ,
    \ces_5_7_io_ins_down[7] ,
    \ces_5_7_io_ins_down[6] ,
    \ces_5_7_io_ins_down[5] ,
    \ces_5_7_io_ins_down[4] ,
    \ces_5_7_io_ins_down[3] ,
    \ces_5_7_io_ins_down[2] ,
    \ces_5_7_io_ins_down[1] ,
    \ces_5_7_io_ins_down[0] }),
    .io_ins_left({net892,
    net891,
    net890,
    net889,
    net887,
    net886,
    net885,
    net884,
    net883,
    net882,
    net881,
    net880,
    net879,
    net878,
    net876,
    net875,
    net874,
    net873,
    net872,
    net871,
    net870,
    net869,
    net868,
    net867,
    net865,
    net864,
    net863,
    net862,
    net861,
    net860,
    net859,
    net858,
    net857,
    net856,
    net854,
    net853,
    net852,
    net851,
    net850,
    net849,
    net848,
    net847,
    net846,
    net845,
    net843,
    net842,
    net841,
    net840,
    net839,
    net838,
    net837,
    net836,
    net835,
    net834,
    net896,
    net895,
    net894,
    net893,
    net888,
    net877,
    net866,
    net855,
    net844,
    net833}),
    .io_ins_right({\ces_5_6_io_outs_right[63] ,
    \ces_5_6_io_outs_right[62] ,
    \ces_5_6_io_outs_right[61] ,
    \ces_5_6_io_outs_right[60] ,
    \ces_5_6_io_outs_right[59] ,
    \ces_5_6_io_outs_right[58] ,
    \ces_5_6_io_outs_right[57] ,
    \ces_5_6_io_outs_right[56] ,
    \ces_5_6_io_outs_right[55] ,
    \ces_5_6_io_outs_right[54] ,
    \ces_5_6_io_outs_right[53] ,
    \ces_5_6_io_outs_right[52] ,
    \ces_5_6_io_outs_right[51] ,
    \ces_5_6_io_outs_right[50] ,
    \ces_5_6_io_outs_right[49] ,
    \ces_5_6_io_outs_right[48] ,
    \ces_5_6_io_outs_right[47] ,
    \ces_5_6_io_outs_right[46] ,
    \ces_5_6_io_outs_right[45] ,
    \ces_5_6_io_outs_right[44] ,
    \ces_5_6_io_outs_right[43] ,
    \ces_5_6_io_outs_right[42] ,
    \ces_5_6_io_outs_right[41] ,
    \ces_5_6_io_outs_right[40] ,
    \ces_5_6_io_outs_right[39] ,
    \ces_5_6_io_outs_right[38] ,
    \ces_5_6_io_outs_right[37] ,
    \ces_5_6_io_outs_right[36] ,
    \ces_5_6_io_outs_right[35] ,
    \ces_5_6_io_outs_right[34] ,
    \ces_5_6_io_outs_right[33] ,
    \ces_5_6_io_outs_right[32] ,
    \ces_5_6_io_outs_right[31] ,
    \ces_5_6_io_outs_right[30] ,
    \ces_5_6_io_outs_right[29] ,
    \ces_5_6_io_outs_right[28] ,
    \ces_5_6_io_outs_right[27] ,
    \ces_5_6_io_outs_right[26] ,
    \ces_5_6_io_outs_right[25] ,
    \ces_5_6_io_outs_right[24] ,
    \ces_5_6_io_outs_right[23] ,
    \ces_5_6_io_outs_right[22] ,
    \ces_5_6_io_outs_right[21] ,
    \ces_5_6_io_outs_right[20] ,
    \ces_5_6_io_outs_right[19] ,
    \ces_5_6_io_outs_right[18] ,
    \ces_5_6_io_outs_right[17] ,
    \ces_5_6_io_outs_right[16] ,
    \ces_5_6_io_outs_right[15] ,
    \ces_5_6_io_outs_right[14] ,
    \ces_5_6_io_outs_right[13] ,
    \ces_5_6_io_outs_right[12] ,
    \ces_5_6_io_outs_right[11] ,
    \ces_5_6_io_outs_right[10] ,
    \ces_5_6_io_outs_right[9] ,
    \ces_5_6_io_outs_right[8] ,
    \ces_5_6_io_outs_right[7] ,
    \ces_5_6_io_outs_right[6] ,
    \ces_5_6_io_outs_right[5] ,
    \ces_5_6_io_outs_right[4] ,
    \ces_5_6_io_outs_right[3] ,
    \ces_5_6_io_outs_right[2] ,
    \ces_5_6_io_outs_right[1] ,
    \ces_5_6_io_outs_right[0] }),
    .io_ins_up({\ces_4_7_io_outs_up[63] ,
    \ces_4_7_io_outs_up[62] ,
    \ces_4_7_io_outs_up[61] ,
    \ces_4_7_io_outs_up[60] ,
    \ces_4_7_io_outs_up[59] ,
    \ces_4_7_io_outs_up[58] ,
    \ces_4_7_io_outs_up[57] ,
    \ces_4_7_io_outs_up[56] ,
    \ces_4_7_io_outs_up[55] ,
    \ces_4_7_io_outs_up[54] ,
    \ces_4_7_io_outs_up[53] ,
    \ces_4_7_io_outs_up[52] ,
    \ces_4_7_io_outs_up[51] ,
    \ces_4_7_io_outs_up[50] ,
    \ces_4_7_io_outs_up[49] ,
    \ces_4_7_io_outs_up[48] ,
    \ces_4_7_io_outs_up[47] ,
    \ces_4_7_io_outs_up[46] ,
    \ces_4_7_io_outs_up[45] ,
    \ces_4_7_io_outs_up[44] ,
    \ces_4_7_io_outs_up[43] ,
    \ces_4_7_io_outs_up[42] ,
    \ces_4_7_io_outs_up[41] ,
    \ces_4_7_io_outs_up[40] ,
    \ces_4_7_io_outs_up[39] ,
    \ces_4_7_io_outs_up[38] ,
    \ces_4_7_io_outs_up[37] ,
    \ces_4_7_io_outs_up[36] ,
    \ces_4_7_io_outs_up[35] ,
    \ces_4_7_io_outs_up[34] ,
    \ces_4_7_io_outs_up[33] ,
    \ces_4_7_io_outs_up[32] ,
    \ces_4_7_io_outs_up[31] ,
    \ces_4_7_io_outs_up[30] ,
    \ces_4_7_io_outs_up[29] ,
    \ces_4_7_io_outs_up[28] ,
    \ces_4_7_io_outs_up[27] ,
    \ces_4_7_io_outs_up[26] ,
    \ces_4_7_io_outs_up[25] ,
    \ces_4_7_io_outs_up[24] ,
    \ces_4_7_io_outs_up[23] ,
    \ces_4_7_io_outs_up[22] ,
    \ces_4_7_io_outs_up[21] ,
    \ces_4_7_io_outs_up[20] ,
    \ces_4_7_io_outs_up[19] ,
    \ces_4_7_io_outs_up[18] ,
    \ces_4_7_io_outs_up[17] ,
    \ces_4_7_io_outs_up[16] ,
    \ces_4_7_io_outs_up[15] ,
    \ces_4_7_io_outs_up[14] ,
    \ces_4_7_io_outs_up[13] ,
    \ces_4_7_io_outs_up[12] ,
    \ces_4_7_io_outs_up[11] ,
    \ces_4_7_io_outs_up[10] ,
    \ces_4_7_io_outs_up[9] ,
    \ces_4_7_io_outs_up[8] ,
    \ces_4_7_io_outs_up[7] ,
    \ces_4_7_io_outs_up[6] ,
    \ces_4_7_io_outs_up[5] ,
    \ces_4_7_io_outs_up[4] ,
    \ces_4_7_io_outs_up[3] ,
    \ces_4_7_io_outs_up[2] ,
    \ces_4_7_io_outs_up[1] ,
    \ces_4_7_io_outs_up[0] }),
    .io_outs_down({\ces_4_7_io_ins_down[63] ,
    \ces_4_7_io_ins_down[62] ,
    \ces_4_7_io_ins_down[61] ,
    \ces_4_7_io_ins_down[60] ,
    \ces_4_7_io_ins_down[59] ,
    \ces_4_7_io_ins_down[58] ,
    \ces_4_7_io_ins_down[57] ,
    \ces_4_7_io_ins_down[56] ,
    \ces_4_7_io_ins_down[55] ,
    \ces_4_7_io_ins_down[54] ,
    \ces_4_7_io_ins_down[53] ,
    \ces_4_7_io_ins_down[52] ,
    \ces_4_7_io_ins_down[51] ,
    \ces_4_7_io_ins_down[50] ,
    \ces_4_7_io_ins_down[49] ,
    \ces_4_7_io_ins_down[48] ,
    \ces_4_7_io_ins_down[47] ,
    \ces_4_7_io_ins_down[46] ,
    \ces_4_7_io_ins_down[45] ,
    \ces_4_7_io_ins_down[44] ,
    \ces_4_7_io_ins_down[43] ,
    \ces_4_7_io_ins_down[42] ,
    \ces_4_7_io_ins_down[41] ,
    \ces_4_7_io_ins_down[40] ,
    \ces_4_7_io_ins_down[39] ,
    \ces_4_7_io_ins_down[38] ,
    \ces_4_7_io_ins_down[37] ,
    \ces_4_7_io_ins_down[36] ,
    \ces_4_7_io_ins_down[35] ,
    \ces_4_7_io_ins_down[34] ,
    \ces_4_7_io_ins_down[33] ,
    \ces_4_7_io_ins_down[32] ,
    \ces_4_7_io_ins_down[31] ,
    \ces_4_7_io_ins_down[30] ,
    \ces_4_7_io_ins_down[29] ,
    \ces_4_7_io_ins_down[28] ,
    \ces_4_7_io_ins_down[27] ,
    \ces_4_7_io_ins_down[26] ,
    \ces_4_7_io_ins_down[25] ,
    \ces_4_7_io_ins_down[24] ,
    \ces_4_7_io_ins_down[23] ,
    \ces_4_7_io_ins_down[22] ,
    \ces_4_7_io_ins_down[21] ,
    \ces_4_7_io_ins_down[20] ,
    \ces_4_7_io_ins_down[19] ,
    \ces_4_7_io_ins_down[18] ,
    \ces_4_7_io_ins_down[17] ,
    \ces_4_7_io_ins_down[16] ,
    \ces_4_7_io_ins_down[15] ,
    \ces_4_7_io_ins_down[14] ,
    \ces_4_7_io_ins_down[13] ,
    \ces_4_7_io_ins_down[12] ,
    \ces_4_7_io_ins_down[11] ,
    \ces_4_7_io_ins_down[10] ,
    \ces_4_7_io_ins_down[9] ,
    \ces_4_7_io_ins_down[8] ,
    \ces_4_7_io_ins_down[7] ,
    \ces_4_7_io_ins_down[6] ,
    \ces_4_7_io_ins_down[5] ,
    \ces_4_7_io_ins_down[4] ,
    \ces_4_7_io_ins_down[3] ,
    \ces_4_7_io_ins_down[2] ,
    \ces_4_7_io_ins_down[1] ,
    \ces_4_7_io_ins_down[0] }),
    .io_outs_left({\ces_5_6_io_ins_left[63] ,
    \ces_5_6_io_ins_left[62] ,
    \ces_5_6_io_ins_left[61] ,
    \ces_5_6_io_ins_left[60] ,
    \ces_5_6_io_ins_left[59] ,
    \ces_5_6_io_ins_left[58] ,
    \ces_5_6_io_ins_left[57] ,
    \ces_5_6_io_ins_left[56] ,
    \ces_5_6_io_ins_left[55] ,
    \ces_5_6_io_ins_left[54] ,
    \ces_5_6_io_ins_left[53] ,
    \ces_5_6_io_ins_left[52] ,
    \ces_5_6_io_ins_left[51] ,
    \ces_5_6_io_ins_left[50] ,
    \ces_5_6_io_ins_left[49] ,
    \ces_5_6_io_ins_left[48] ,
    \ces_5_6_io_ins_left[47] ,
    \ces_5_6_io_ins_left[46] ,
    \ces_5_6_io_ins_left[45] ,
    \ces_5_6_io_ins_left[44] ,
    \ces_5_6_io_ins_left[43] ,
    \ces_5_6_io_ins_left[42] ,
    \ces_5_6_io_ins_left[41] ,
    \ces_5_6_io_ins_left[40] ,
    \ces_5_6_io_ins_left[39] ,
    \ces_5_6_io_ins_left[38] ,
    \ces_5_6_io_ins_left[37] ,
    \ces_5_6_io_ins_left[36] ,
    \ces_5_6_io_ins_left[35] ,
    \ces_5_6_io_ins_left[34] ,
    \ces_5_6_io_ins_left[33] ,
    \ces_5_6_io_ins_left[32] ,
    \ces_5_6_io_ins_left[31] ,
    \ces_5_6_io_ins_left[30] ,
    \ces_5_6_io_ins_left[29] ,
    \ces_5_6_io_ins_left[28] ,
    \ces_5_6_io_ins_left[27] ,
    \ces_5_6_io_ins_left[26] ,
    \ces_5_6_io_ins_left[25] ,
    \ces_5_6_io_ins_left[24] ,
    \ces_5_6_io_ins_left[23] ,
    \ces_5_6_io_ins_left[22] ,
    \ces_5_6_io_ins_left[21] ,
    \ces_5_6_io_ins_left[20] ,
    \ces_5_6_io_ins_left[19] ,
    \ces_5_6_io_ins_left[18] ,
    \ces_5_6_io_ins_left[17] ,
    \ces_5_6_io_ins_left[16] ,
    \ces_5_6_io_ins_left[15] ,
    \ces_5_6_io_ins_left[14] ,
    \ces_5_6_io_ins_left[13] ,
    \ces_5_6_io_ins_left[12] ,
    \ces_5_6_io_ins_left[11] ,
    \ces_5_6_io_ins_left[10] ,
    \ces_5_6_io_ins_left[9] ,
    \ces_5_6_io_ins_left[8] ,
    \ces_5_6_io_ins_left[7] ,
    \ces_5_6_io_ins_left[6] ,
    \ces_5_6_io_ins_left[5] ,
    \ces_5_6_io_ins_left[4] ,
    \ces_5_6_io_ins_left[3] ,
    \ces_5_6_io_ins_left[2] ,
    \ces_5_6_io_ins_left[1] ,
    \ces_5_6_io_ins_left[0] }),
    .io_outs_right({net3516,
    net3515,
    net3514,
    net3513,
    net3511,
    net3510,
    net3509,
    net3508,
    net3507,
    net3506,
    net3505,
    net3504,
    net3503,
    net3502,
    net3500,
    net3499,
    net3498,
    net3497,
    net3496,
    net3495,
    net3494,
    net3493,
    net3492,
    net3491,
    net3489,
    net3488,
    net3487,
    net3486,
    net3485,
    net3484,
    net3483,
    net3482,
    net3481,
    net3480,
    net3478,
    net3477,
    net3476,
    net3475,
    net3474,
    net3473,
    net3472,
    net3471,
    net3470,
    net3469,
    net3467,
    net3466,
    net3465,
    net3464,
    net3463,
    net3462,
    net3461,
    net3460,
    net3459,
    net3458,
    net3520,
    net3519,
    net3518,
    net3517,
    net3512,
    net3501,
    net3490,
    net3479,
    net3468,
    net3457}),
    .io_outs_up({\ces_5_7_io_outs_up[63] ,
    \ces_5_7_io_outs_up[62] ,
    \ces_5_7_io_outs_up[61] ,
    \ces_5_7_io_outs_up[60] ,
    \ces_5_7_io_outs_up[59] ,
    \ces_5_7_io_outs_up[58] ,
    \ces_5_7_io_outs_up[57] ,
    \ces_5_7_io_outs_up[56] ,
    \ces_5_7_io_outs_up[55] ,
    \ces_5_7_io_outs_up[54] ,
    \ces_5_7_io_outs_up[53] ,
    \ces_5_7_io_outs_up[52] ,
    \ces_5_7_io_outs_up[51] ,
    \ces_5_7_io_outs_up[50] ,
    \ces_5_7_io_outs_up[49] ,
    \ces_5_7_io_outs_up[48] ,
    \ces_5_7_io_outs_up[47] ,
    \ces_5_7_io_outs_up[46] ,
    \ces_5_7_io_outs_up[45] ,
    \ces_5_7_io_outs_up[44] ,
    \ces_5_7_io_outs_up[43] ,
    \ces_5_7_io_outs_up[42] ,
    \ces_5_7_io_outs_up[41] ,
    \ces_5_7_io_outs_up[40] ,
    \ces_5_7_io_outs_up[39] ,
    \ces_5_7_io_outs_up[38] ,
    \ces_5_7_io_outs_up[37] ,
    \ces_5_7_io_outs_up[36] ,
    \ces_5_7_io_outs_up[35] ,
    \ces_5_7_io_outs_up[34] ,
    \ces_5_7_io_outs_up[33] ,
    \ces_5_7_io_outs_up[32] ,
    \ces_5_7_io_outs_up[31] ,
    \ces_5_7_io_outs_up[30] ,
    \ces_5_7_io_outs_up[29] ,
    \ces_5_7_io_outs_up[28] ,
    \ces_5_7_io_outs_up[27] ,
    \ces_5_7_io_outs_up[26] ,
    \ces_5_7_io_outs_up[25] ,
    \ces_5_7_io_outs_up[24] ,
    \ces_5_7_io_outs_up[23] ,
    \ces_5_7_io_outs_up[22] ,
    \ces_5_7_io_outs_up[21] ,
    \ces_5_7_io_outs_up[20] ,
    \ces_5_7_io_outs_up[19] ,
    \ces_5_7_io_outs_up[18] ,
    \ces_5_7_io_outs_up[17] ,
    \ces_5_7_io_outs_up[16] ,
    \ces_5_7_io_outs_up[15] ,
    \ces_5_7_io_outs_up[14] ,
    \ces_5_7_io_outs_up[13] ,
    \ces_5_7_io_outs_up[12] ,
    \ces_5_7_io_outs_up[11] ,
    \ces_5_7_io_outs_up[10] ,
    \ces_5_7_io_outs_up[9] ,
    \ces_5_7_io_outs_up[8] ,
    \ces_5_7_io_outs_up[7] ,
    \ces_5_7_io_outs_up[6] ,
    \ces_5_7_io_outs_up[5] ,
    \ces_5_7_io_outs_up[4] ,
    \ces_5_7_io_outs_up[3] ,
    \ces_5_7_io_outs_up[2] ,
    \ces_5_7_io_outs_up[1] ,
    \ces_5_7_io_outs_up[0] }));
 Element ces_6_0 (.clock(clknet_3_5_0_clock),
    .io_lsbIns_1(net4203),
    .io_lsbIns_2(net4204),
    .io_lsbIns_3(net4205),
    .io_lsbIns_4(net4206),
    .io_lsbIns_5(net4207),
    .io_lsbIns_6(net4208),
    .io_lsbIns_7(net4209),
    .io_lsbOuts_0(ces_6_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_0_io_lsbOuts_7),
    .io_ins_down({\ces_6_0_io_ins_down[63] ,
    \ces_6_0_io_ins_down[62] ,
    \ces_6_0_io_ins_down[61] ,
    \ces_6_0_io_ins_down[60] ,
    \ces_6_0_io_ins_down[59] ,
    \ces_6_0_io_ins_down[58] ,
    \ces_6_0_io_ins_down[57] ,
    \ces_6_0_io_ins_down[56] ,
    \ces_6_0_io_ins_down[55] ,
    \ces_6_0_io_ins_down[54] ,
    \ces_6_0_io_ins_down[53] ,
    \ces_6_0_io_ins_down[52] ,
    \ces_6_0_io_ins_down[51] ,
    \ces_6_0_io_ins_down[50] ,
    \ces_6_0_io_ins_down[49] ,
    \ces_6_0_io_ins_down[48] ,
    \ces_6_0_io_ins_down[47] ,
    \ces_6_0_io_ins_down[46] ,
    \ces_6_0_io_ins_down[45] ,
    \ces_6_0_io_ins_down[44] ,
    \ces_6_0_io_ins_down[43] ,
    \ces_6_0_io_ins_down[42] ,
    \ces_6_0_io_ins_down[41] ,
    \ces_6_0_io_ins_down[40] ,
    \ces_6_0_io_ins_down[39] ,
    \ces_6_0_io_ins_down[38] ,
    \ces_6_0_io_ins_down[37] ,
    \ces_6_0_io_ins_down[36] ,
    \ces_6_0_io_ins_down[35] ,
    \ces_6_0_io_ins_down[34] ,
    \ces_6_0_io_ins_down[33] ,
    \ces_6_0_io_ins_down[32] ,
    \ces_6_0_io_ins_down[31] ,
    \ces_6_0_io_ins_down[30] ,
    \ces_6_0_io_ins_down[29] ,
    \ces_6_0_io_ins_down[28] ,
    \ces_6_0_io_ins_down[27] ,
    \ces_6_0_io_ins_down[26] ,
    \ces_6_0_io_ins_down[25] ,
    \ces_6_0_io_ins_down[24] ,
    \ces_6_0_io_ins_down[23] ,
    \ces_6_0_io_ins_down[22] ,
    \ces_6_0_io_ins_down[21] ,
    \ces_6_0_io_ins_down[20] ,
    \ces_6_0_io_ins_down[19] ,
    \ces_6_0_io_ins_down[18] ,
    \ces_6_0_io_ins_down[17] ,
    \ces_6_0_io_ins_down[16] ,
    \ces_6_0_io_ins_down[15] ,
    \ces_6_0_io_ins_down[14] ,
    \ces_6_0_io_ins_down[13] ,
    \ces_6_0_io_ins_down[12] ,
    \ces_6_0_io_ins_down[11] ,
    \ces_6_0_io_ins_down[10] ,
    \ces_6_0_io_ins_down[9] ,
    \ces_6_0_io_ins_down[8] ,
    \ces_6_0_io_ins_down[7] ,
    \ces_6_0_io_ins_down[6] ,
    \ces_6_0_io_ins_down[5] ,
    \ces_6_0_io_ins_down[4] ,
    \ces_6_0_io_ins_down[3] ,
    \ces_6_0_io_ins_down[2] ,
    \ces_6_0_io_ins_down[1] ,
    \ces_6_0_io_ins_down[0] }),
    .io_ins_left({\ces_6_0_io_ins_left[63] ,
    \ces_6_0_io_ins_left[62] ,
    \ces_6_0_io_ins_left[61] ,
    \ces_6_0_io_ins_left[60] ,
    \ces_6_0_io_ins_left[59] ,
    \ces_6_0_io_ins_left[58] ,
    \ces_6_0_io_ins_left[57] ,
    \ces_6_0_io_ins_left[56] ,
    \ces_6_0_io_ins_left[55] ,
    \ces_6_0_io_ins_left[54] ,
    \ces_6_0_io_ins_left[53] ,
    \ces_6_0_io_ins_left[52] ,
    \ces_6_0_io_ins_left[51] ,
    \ces_6_0_io_ins_left[50] ,
    \ces_6_0_io_ins_left[49] ,
    \ces_6_0_io_ins_left[48] ,
    \ces_6_0_io_ins_left[47] ,
    \ces_6_0_io_ins_left[46] ,
    \ces_6_0_io_ins_left[45] ,
    \ces_6_0_io_ins_left[44] ,
    \ces_6_0_io_ins_left[43] ,
    \ces_6_0_io_ins_left[42] ,
    \ces_6_0_io_ins_left[41] ,
    \ces_6_0_io_ins_left[40] ,
    \ces_6_0_io_ins_left[39] ,
    \ces_6_0_io_ins_left[38] ,
    \ces_6_0_io_ins_left[37] ,
    \ces_6_0_io_ins_left[36] ,
    \ces_6_0_io_ins_left[35] ,
    \ces_6_0_io_ins_left[34] ,
    \ces_6_0_io_ins_left[33] ,
    \ces_6_0_io_ins_left[32] ,
    \ces_6_0_io_ins_left[31] ,
    \ces_6_0_io_ins_left[30] ,
    \ces_6_0_io_ins_left[29] ,
    \ces_6_0_io_ins_left[28] ,
    \ces_6_0_io_ins_left[27] ,
    \ces_6_0_io_ins_left[26] ,
    \ces_6_0_io_ins_left[25] ,
    \ces_6_0_io_ins_left[24] ,
    \ces_6_0_io_ins_left[23] ,
    \ces_6_0_io_ins_left[22] ,
    \ces_6_0_io_ins_left[21] ,
    \ces_6_0_io_ins_left[20] ,
    \ces_6_0_io_ins_left[19] ,
    \ces_6_0_io_ins_left[18] ,
    \ces_6_0_io_ins_left[17] ,
    \ces_6_0_io_ins_left[16] ,
    \ces_6_0_io_ins_left[15] ,
    \ces_6_0_io_ins_left[14] ,
    \ces_6_0_io_ins_left[13] ,
    \ces_6_0_io_ins_left[12] ,
    \ces_6_0_io_ins_left[11] ,
    \ces_6_0_io_ins_left[10] ,
    \ces_6_0_io_ins_left[9] ,
    \ces_6_0_io_ins_left[8] ,
    \ces_6_0_io_ins_left[7] ,
    \ces_6_0_io_ins_left[6] ,
    \ces_6_0_io_ins_left[5] ,
    \ces_6_0_io_ins_left[4] ,
    \ces_6_0_io_ins_left[3] ,
    \ces_6_0_io_ins_left[2] ,
    \ces_6_0_io_ins_left[1] ,
    \ces_6_0_io_ins_left[0] }),
    .io_ins_right({net1468,
    net1467,
    net1466,
    net1465,
    net1463,
    net1462,
    net1461,
    net1460,
    net1459,
    net1458,
    net1457,
    net1456,
    net1455,
    net1454,
    net1452,
    net1451,
    net1450,
    net1449,
    net1448,
    net1447,
    net1446,
    net1445,
    net1444,
    net1443,
    net1441,
    net1440,
    net1439,
    net1438,
    net1437,
    net1436,
    net1435,
    net1434,
    net1433,
    net1432,
    net1430,
    net1429,
    net1428,
    net1427,
    net1426,
    net1425,
    net1424,
    net1423,
    net1422,
    net1421,
    net1419,
    net1418,
    net1417,
    net1416,
    net1415,
    net1414,
    net1413,
    net1412,
    net1411,
    net1410,
    net1472,
    net1471,
    net1470,
    net1469,
    net1464,
    net1453,
    net1442,
    net1431,
    net1420,
    net1409}),
    .io_ins_up({\ces_5_0_io_outs_up[63] ,
    \ces_5_0_io_outs_up[62] ,
    \ces_5_0_io_outs_up[61] ,
    \ces_5_0_io_outs_up[60] ,
    \ces_5_0_io_outs_up[59] ,
    \ces_5_0_io_outs_up[58] ,
    \ces_5_0_io_outs_up[57] ,
    \ces_5_0_io_outs_up[56] ,
    \ces_5_0_io_outs_up[55] ,
    \ces_5_0_io_outs_up[54] ,
    \ces_5_0_io_outs_up[53] ,
    \ces_5_0_io_outs_up[52] ,
    \ces_5_0_io_outs_up[51] ,
    \ces_5_0_io_outs_up[50] ,
    \ces_5_0_io_outs_up[49] ,
    \ces_5_0_io_outs_up[48] ,
    \ces_5_0_io_outs_up[47] ,
    \ces_5_0_io_outs_up[46] ,
    \ces_5_0_io_outs_up[45] ,
    \ces_5_0_io_outs_up[44] ,
    \ces_5_0_io_outs_up[43] ,
    \ces_5_0_io_outs_up[42] ,
    \ces_5_0_io_outs_up[41] ,
    \ces_5_0_io_outs_up[40] ,
    \ces_5_0_io_outs_up[39] ,
    \ces_5_0_io_outs_up[38] ,
    \ces_5_0_io_outs_up[37] ,
    \ces_5_0_io_outs_up[36] ,
    \ces_5_0_io_outs_up[35] ,
    \ces_5_0_io_outs_up[34] ,
    \ces_5_0_io_outs_up[33] ,
    \ces_5_0_io_outs_up[32] ,
    \ces_5_0_io_outs_up[31] ,
    \ces_5_0_io_outs_up[30] ,
    \ces_5_0_io_outs_up[29] ,
    \ces_5_0_io_outs_up[28] ,
    \ces_5_0_io_outs_up[27] ,
    \ces_5_0_io_outs_up[26] ,
    \ces_5_0_io_outs_up[25] ,
    \ces_5_0_io_outs_up[24] ,
    \ces_5_0_io_outs_up[23] ,
    \ces_5_0_io_outs_up[22] ,
    \ces_5_0_io_outs_up[21] ,
    \ces_5_0_io_outs_up[20] ,
    \ces_5_0_io_outs_up[19] ,
    \ces_5_0_io_outs_up[18] ,
    \ces_5_0_io_outs_up[17] ,
    \ces_5_0_io_outs_up[16] ,
    \ces_5_0_io_outs_up[15] ,
    \ces_5_0_io_outs_up[14] ,
    \ces_5_0_io_outs_up[13] ,
    \ces_5_0_io_outs_up[12] ,
    \ces_5_0_io_outs_up[11] ,
    \ces_5_0_io_outs_up[10] ,
    \ces_5_0_io_outs_up[9] ,
    \ces_5_0_io_outs_up[8] ,
    \ces_5_0_io_outs_up[7] ,
    \ces_5_0_io_outs_up[6] ,
    \ces_5_0_io_outs_up[5] ,
    \ces_5_0_io_outs_up[4] ,
    \ces_5_0_io_outs_up[3] ,
    \ces_5_0_io_outs_up[2] ,
    \ces_5_0_io_outs_up[1] ,
    \ces_5_0_io_outs_up[0] }),
    .io_outs_down({\ces_5_0_io_ins_down[63] ,
    \ces_5_0_io_ins_down[62] ,
    \ces_5_0_io_ins_down[61] ,
    \ces_5_0_io_ins_down[60] ,
    \ces_5_0_io_ins_down[59] ,
    \ces_5_0_io_ins_down[58] ,
    \ces_5_0_io_ins_down[57] ,
    \ces_5_0_io_ins_down[56] ,
    \ces_5_0_io_ins_down[55] ,
    \ces_5_0_io_ins_down[54] ,
    \ces_5_0_io_ins_down[53] ,
    \ces_5_0_io_ins_down[52] ,
    \ces_5_0_io_ins_down[51] ,
    \ces_5_0_io_ins_down[50] ,
    \ces_5_0_io_ins_down[49] ,
    \ces_5_0_io_ins_down[48] ,
    \ces_5_0_io_ins_down[47] ,
    \ces_5_0_io_ins_down[46] ,
    \ces_5_0_io_ins_down[45] ,
    \ces_5_0_io_ins_down[44] ,
    \ces_5_0_io_ins_down[43] ,
    \ces_5_0_io_ins_down[42] ,
    \ces_5_0_io_ins_down[41] ,
    \ces_5_0_io_ins_down[40] ,
    \ces_5_0_io_ins_down[39] ,
    \ces_5_0_io_ins_down[38] ,
    \ces_5_0_io_ins_down[37] ,
    \ces_5_0_io_ins_down[36] ,
    \ces_5_0_io_ins_down[35] ,
    \ces_5_0_io_ins_down[34] ,
    \ces_5_0_io_ins_down[33] ,
    \ces_5_0_io_ins_down[32] ,
    \ces_5_0_io_ins_down[31] ,
    \ces_5_0_io_ins_down[30] ,
    \ces_5_0_io_ins_down[29] ,
    \ces_5_0_io_ins_down[28] ,
    \ces_5_0_io_ins_down[27] ,
    \ces_5_0_io_ins_down[26] ,
    \ces_5_0_io_ins_down[25] ,
    \ces_5_0_io_ins_down[24] ,
    \ces_5_0_io_ins_down[23] ,
    \ces_5_0_io_ins_down[22] ,
    \ces_5_0_io_ins_down[21] ,
    \ces_5_0_io_ins_down[20] ,
    \ces_5_0_io_ins_down[19] ,
    \ces_5_0_io_ins_down[18] ,
    \ces_5_0_io_ins_down[17] ,
    \ces_5_0_io_ins_down[16] ,
    \ces_5_0_io_ins_down[15] ,
    \ces_5_0_io_ins_down[14] ,
    \ces_5_0_io_ins_down[13] ,
    \ces_5_0_io_ins_down[12] ,
    \ces_5_0_io_ins_down[11] ,
    \ces_5_0_io_ins_down[10] ,
    \ces_5_0_io_ins_down[9] ,
    \ces_5_0_io_ins_down[8] ,
    \ces_5_0_io_ins_down[7] ,
    \ces_5_0_io_ins_down[6] ,
    \ces_5_0_io_ins_down[5] ,
    \ces_5_0_io_ins_down[4] ,
    \ces_5_0_io_ins_down[3] ,
    \ces_5_0_io_ins_down[2] ,
    \ces_5_0_io_ins_down[1] ,
    \ces_5_0_io_ins_down[0] }),
    .io_outs_left({net3068,
    net3067,
    net3066,
    net3065,
    net3063,
    net3062,
    net3061,
    net3060,
    net3059,
    net3058,
    net3057,
    net3056,
    net3055,
    net3054,
    net3052,
    net3051,
    net3050,
    net3049,
    net3048,
    net3047,
    net3046,
    net3045,
    net3044,
    net3043,
    net3041,
    net3040,
    net3039,
    net3038,
    net3037,
    net3036,
    net3035,
    net3034,
    net3033,
    net3032,
    net3030,
    net3029,
    net3028,
    net3027,
    net3026,
    net3025,
    net3024,
    net3023,
    net3022,
    net3021,
    net3019,
    net3018,
    net3017,
    net3016,
    net3015,
    net3014,
    net3013,
    net3012,
    net3011,
    net3010,
    net3072,
    net3071,
    net3070,
    net3069,
    net3064,
    net3053,
    net3042,
    net3031,
    net3020,
    net3009}),
    .io_outs_right({\ces_6_0_io_outs_right[63] ,
    \ces_6_0_io_outs_right[62] ,
    \ces_6_0_io_outs_right[61] ,
    \ces_6_0_io_outs_right[60] ,
    \ces_6_0_io_outs_right[59] ,
    \ces_6_0_io_outs_right[58] ,
    \ces_6_0_io_outs_right[57] ,
    \ces_6_0_io_outs_right[56] ,
    \ces_6_0_io_outs_right[55] ,
    \ces_6_0_io_outs_right[54] ,
    \ces_6_0_io_outs_right[53] ,
    \ces_6_0_io_outs_right[52] ,
    \ces_6_0_io_outs_right[51] ,
    \ces_6_0_io_outs_right[50] ,
    \ces_6_0_io_outs_right[49] ,
    \ces_6_0_io_outs_right[48] ,
    \ces_6_0_io_outs_right[47] ,
    \ces_6_0_io_outs_right[46] ,
    \ces_6_0_io_outs_right[45] ,
    \ces_6_0_io_outs_right[44] ,
    \ces_6_0_io_outs_right[43] ,
    \ces_6_0_io_outs_right[42] ,
    \ces_6_0_io_outs_right[41] ,
    \ces_6_0_io_outs_right[40] ,
    \ces_6_0_io_outs_right[39] ,
    \ces_6_0_io_outs_right[38] ,
    \ces_6_0_io_outs_right[37] ,
    \ces_6_0_io_outs_right[36] ,
    \ces_6_0_io_outs_right[35] ,
    \ces_6_0_io_outs_right[34] ,
    \ces_6_0_io_outs_right[33] ,
    \ces_6_0_io_outs_right[32] ,
    \ces_6_0_io_outs_right[31] ,
    \ces_6_0_io_outs_right[30] ,
    \ces_6_0_io_outs_right[29] ,
    \ces_6_0_io_outs_right[28] ,
    \ces_6_0_io_outs_right[27] ,
    \ces_6_0_io_outs_right[26] ,
    \ces_6_0_io_outs_right[25] ,
    \ces_6_0_io_outs_right[24] ,
    \ces_6_0_io_outs_right[23] ,
    \ces_6_0_io_outs_right[22] ,
    \ces_6_0_io_outs_right[21] ,
    \ces_6_0_io_outs_right[20] ,
    \ces_6_0_io_outs_right[19] ,
    \ces_6_0_io_outs_right[18] ,
    \ces_6_0_io_outs_right[17] ,
    \ces_6_0_io_outs_right[16] ,
    \ces_6_0_io_outs_right[15] ,
    \ces_6_0_io_outs_right[14] ,
    \ces_6_0_io_outs_right[13] ,
    \ces_6_0_io_outs_right[12] ,
    \ces_6_0_io_outs_right[11] ,
    \ces_6_0_io_outs_right[10] ,
    \ces_6_0_io_outs_right[9] ,
    \ces_6_0_io_outs_right[8] ,
    \ces_6_0_io_outs_right[7] ,
    \ces_6_0_io_outs_right[6] ,
    \ces_6_0_io_outs_right[5] ,
    \ces_6_0_io_outs_right[4] ,
    \ces_6_0_io_outs_right[3] ,
    \ces_6_0_io_outs_right[2] ,
    \ces_6_0_io_outs_right[1] ,
    \ces_6_0_io_outs_right[0] }),
    .io_outs_up({\ces_6_0_io_outs_up[63] ,
    \ces_6_0_io_outs_up[62] ,
    \ces_6_0_io_outs_up[61] ,
    \ces_6_0_io_outs_up[60] ,
    \ces_6_0_io_outs_up[59] ,
    \ces_6_0_io_outs_up[58] ,
    \ces_6_0_io_outs_up[57] ,
    \ces_6_0_io_outs_up[56] ,
    \ces_6_0_io_outs_up[55] ,
    \ces_6_0_io_outs_up[54] ,
    \ces_6_0_io_outs_up[53] ,
    \ces_6_0_io_outs_up[52] ,
    \ces_6_0_io_outs_up[51] ,
    \ces_6_0_io_outs_up[50] ,
    \ces_6_0_io_outs_up[49] ,
    \ces_6_0_io_outs_up[48] ,
    \ces_6_0_io_outs_up[47] ,
    \ces_6_0_io_outs_up[46] ,
    \ces_6_0_io_outs_up[45] ,
    \ces_6_0_io_outs_up[44] ,
    \ces_6_0_io_outs_up[43] ,
    \ces_6_0_io_outs_up[42] ,
    \ces_6_0_io_outs_up[41] ,
    \ces_6_0_io_outs_up[40] ,
    \ces_6_0_io_outs_up[39] ,
    \ces_6_0_io_outs_up[38] ,
    \ces_6_0_io_outs_up[37] ,
    \ces_6_0_io_outs_up[36] ,
    \ces_6_0_io_outs_up[35] ,
    \ces_6_0_io_outs_up[34] ,
    \ces_6_0_io_outs_up[33] ,
    \ces_6_0_io_outs_up[32] ,
    \ces_6_0_io_outs_up[31] ,
    \ces_6_0_io_outs_up[30] ,
    \ces_6_0_io_outs_up[29] ,
    \ces_6_0_io_outs_up[28] ,
    \ces_6_0_io_outs_up[27] ,
    \ces_6_0_io_outs_up[26] ,
    \ces_6_0_io_outs_up[25] ,
    \ces_6_0_io_outs_up[24] ,
    \ces_6_0_io_outs_up[23] ,
    \ces_6_0_io_outs_up[22] ,
    \ces_6_0_io_outs_up[21] ,
    \ces_6_0_io_outs_up[20] ,
    \ces_6_0_io_outs_up[19] ,
    \ces_6_0_io_outs_up[18] ,
    \ces_6_0_io_outs_up[17] ,
    \ces_6_0_io_outs_up[16] ,
    \ces_6_0_io_outs_up[15] ,
    \ces_6_0_io_outs_up[14] ,
    \ces_6_0_io_outs_up[13] ,
    \ces_6_0_io_outs_up[12] ,
    \ces_6_0_io_outs_up[11] ,
    \ces_6_0_io_outs_up[10] ,
    \ces_6_0_io_outs_up[9] ,
    \ces_6_0_io_outs_up[8] ,
    \ces_6_0_io_outs_up[7] ,
    \ces_6_0_io_outs_up[6] ,
    \ces_6_0_io_outs_up[5] ,
    \ces_6_0_io_outs_up[4] ,
    \ces_6_0_io_outs_up[3] ,
    \ces_6_0_io_outs_up[2] ,
    \ces_6_0_io_outs_up[1] ,
    \ces_6_0_io_outs_up[0] }));
 Element ces_6_1 (.clock(clknet_3_5_0_clock),
    .io_lsbIns_1(ces_6_0_io_lsbOuts_1),
    .io_lsbIns_2(ces_6_0_io_lsbOuts_2),
    .io_lsbIns_3(ces_6_0_io_lsbOuts_3),
    .io_lsbIns_4(ces_6_0_io_lsbOuts_4),
    .io_lsbIns_5(ces_6_0_io_lsbOuts_5),
    .io_lsbIns_6(ces_6_0_io_lsbOuts_6),
    .io_lsbIns_7(ces_6_0_io_lsbOuts_7),
    .io_lsbOuts_0(ces_6_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_1_io_lsbOuts_7),
    .io_ins_down({\ces_6_1_io_ins_down[63] ,
    \ces_6_1_io_ins_down[62] ,
    \ces_6_1_io_ins_down[61] ,
    \ces_6_1_io_ins_down[60] ,
    \ces_6_1_io_ins_down[59] ,
    \ces_6_1_io_ins_down[58] ,
    \ces_6_1_io_ins_down[57] ,
    \ces_6_1_io_ins_down[56] ,
    \ces_6_1_io_ins_down[55] ,
    \ces_6_1_io_ins_down[54] ,
    \ces_6_1_io_ins_down[53] ,
    \ces_6_1_io_ins_down[52] ,
    \ces_6_1_io_ins_down[51] ,
    \ces_6_1_io_ins_down[50] ,
    \ces_6_1_io_ins_down[49] ,
    \ces_6_1_io_ins_down[48] ,
    \ces_6_1_io_ins_down[47] ,
    \ces_6_1_io_ins_down[46] ,
    \ces_6_1_io_ins_down[45] ,
    \ces_6_1_io_ins_down[44] ,
    \ces_6_1_io_ins_down[43] ,
    \ces_6_1_io_ins_down[42] ,
    \ces_6_1_io_ins_down[41] ,
    \ces_6_1_io_ins_down[40] ,
    \ces_6_1_io_ins_down[39] ,
    \ces_6_1_io_ins_down[38] ,
    \ces_6_1_io_ins_down[37] ,
    \ces_6_1_io_ins_down[36] ,
    \ces_6_1_io_ins_down[35] ,
    \ces_6_1_io_ins_down[34] ,
    \ces_6_1_io_ins_down[33] ,
    \ces_6_1_io_ins_down[32] ,
    \ces_6_1_io_ins_down[31] ,
    \ces_6_1_io_ins_down[30] ,
    \ces_6_1_io_ins_down[29] ,
    \ces_6_1_io_ins_down[28] ,
    \ces_6_1_io_ins_down[27] ,
    \ces_6_1_io_ins_down[26] ,
    \ces_6_1_io_ins_down[25] ,
    \ces_6_1_io_ins_down[24] ,
    \ces_6_1_io_ins_down[23] ,
    \ces_6_1_io_ins_down[22] ,
    \ces_6_1_io_ins_down[21] ,
    \ces_6_1_io_ins_down[20] ,
    \ces_6_1_io_ins_down[19] ,
    \ces_6_1_io_ins_down[18] ,
    \ces_6_1_io_ins_down[17] ,
    \ces_6_1_io_ins_down[16] ,
    \ces_6_1_io_ins_down[15] ,
    \ces_6_1_io_ins_down[14] ,
    \ces_6_1_io_ins_down[13] ,
    \ces_6_1_io_ins_down[12] ,
    \ces_6_1_io_ins_down[11] ,
    \ces_6_1_io_ins_down[10] ,
    \ces_6_1_io_ins_down[9] ,
    \ces_6_1_io_ins_down[8] ,
    \ces_6_1_io_ins_down[7] ,
    \ces_6_1_io_ins_down[6] ,
    \ces_6_1_io_ins_down[5] ,
    \ces_6_1_io_ins_down[4] ,
    \ces_6_1_io_ins_down[3] ,
    \ces_6_1_io_ins_down[2] ,
    \ces_6_1_io_ins_down[1] ,
    \ces_6_1_io_ins_down[0] }),
    .io_ins_left({\ces_6_1_io_ins_left[63] ,
    \ces_6_1_io_ins_left[62] ,
    \ces_6_1_io_ins_left[61] ,
    \ces_6_1_io_ins_left[60] ,
    \ces_6_1_io_ins_left[59] ,
    \ces_6_1_io_ins_left[58] ,
    \ces_6_1_io_ins_left[57] ,
    \ces_6_1_io_ins_left[56] ,
    \ces_6_1_io_ins_left[55] ,
    \ces_6_1_io_ins_left[54] ,
    \ces_6_1_io_ins_left[53] ,
    \ces_6_1_io_ins_left[52] ,
    \ces_6_1_io_ins_left[51] ,
    \ces_6_1_io_ins_left[50] ,
    \ces_6_1_io_ins_left[49] ,
    \ces_6_1_io_ins_left[48] ,
    \ces_6_1_io_ins_left[47] ,
    \ces_6_1_io_ins_left[46] ,
    \ces_6_1_io_ins_left[45] ,
    \ces_6_1_io_ins_left[44] ,
    \ces_6_1_io_ins_left[43] ,
    \ces_6_1_io_ins_left[42] ,
    \ces_6_1_io_ins_left[41] ,
    \ces_6_1_io_ins_left[40] ,
    \ces_6_1_io_ins_left[39] ,
    \ces_6_1_io_ins_left[38] ,
    \ces_6_1_io_ins_left[37] ,
    \ces_6_1_io_ins_left[36] ,
    \ces_6_1_io_ins_left[35] ,
    \ces_6_1_io_ins_left[34] ,
    \ces_6_1_io_ins_left[33] ,
    \ces_6_1_io_ins_left[32] ,
    \ces_6_1_io_ins_left[31] ,
    \ces_6_1_io_ins_left[30] ,
    \ces_6_1_io_ins_left[29] ,
    \ces_6_1_io_ins_left[28] ,
    \ces_6_1_io_ins_left[27] ,
    \ces_6_1_io_ins_left[26] ,
    \ces_6_1_io_ins_left[25] ,
    \ces_6_1_io_ins_left[24] ,
    \ces_6_1_io_ins_left[23] ,
    \ces_6_1_io_ins_left[22] ,
    \ces_6_1_io_ins_left[21] ,
    \ces_6_1_io_ins_left[20] ,
    \ces_6_1_io_ins_left[19] ,
    \ces_6_1_io_ins_left[18] ,
    \ces_6_1_io_ins_left[17] ,
    \ces_6_1_io_ins_left[16] ,
    \ces_6_1_io_ins_left[15] ,
    \ces_6_1_io_ins_left[14] ,
    \ces_6_1_io_ins_left[13] ,
    \ces_6_1_io_ins_left[12] ,
    \ces_6_1_io_ins_left[11] ,
    \ces_6_1_io_ins_left[10] ,
    \ces_6_1_io_ins_left[9] ,
    \ces_6_1_io_ins_left[8] ,
    \ces_6_1_io_ins_left[7] ,
    \ces_6_1_io_ins_left[6] ,
    \ces_6_1_io_ins_left[5] ,
    \ces_6_1_io_ins_left[4] ,
    \ces_6_1_io_ins_left[3] ,
    \ces_6_1_io_ins_left[2] ,
    \ces_6_1_io_ins_left[1] ,
    \ces_6_1_io_ins_left[0] }),
    .io_ins_right({\ces_6_0_io_outs_right[63] ,
    \ces_6_0_io_outs_right[62] ,
    \ces_6_0_io_outs_right[61] ,
    \ces_6_0_io_outs_right[60] ,
    \ces_6_0_io_outs_right[59] ,
    \ces_6_0_io_outs_right[58] ,
    \ces_6_0_io_outs_right[57] ,
    \ces_6_0_io_outs_right[56] ,
    \ces_6_0_io_outs_right[55] ,
    \ces_6_0_io_outs_right[54] ,
    \ces_6_0_io_outs_right[53] ,
    \ces_6_0_io_outs_right[52] ,
    \ces_6_0_io_outs_right[51] ,
    \ces_6_0_io_outs_right[50] ,
    \ces_6_0_io_outs_right[49] ,
    \ces_6_0_io_outs_right[48] ,
    \ces_6_0_io_outs_right[47] ,
    \ces_6_0_io_outs_right[46] ,
    \ces_6_0_io_outs_right[45] ,
    \ces_6_0_io_outs_right[44] ,
    \ces_6_0_io_outs_right[43] ,
    \ces_6_0_io_outs_right[42] ,
    \ces_6_0_io_outs_right[41] ,
    \ces_6_0_io_outs_right[40] ,
    \ces_6_0_io_outs_right[39] ,
    \ces_6_0_io_outs_right[38] ,
    \ces_6_0_io_outs_right[37] ,
    \ces_6_0_io_outs_right[36] ,
    \ces_6_0_io_outs_right[35] ,
    \ces_6_0_io_outs_right[34] ,
    \ces_6_0_io_outs_right[33] ,
    \ces_6_0_io_outs_right[32] ,
    \ces_6_0_io_outs_right[31] ,
    \ces_6_0_io_outs_right[30] ,
    \ces_6_0_io_outs_right[29] ,
    \ces_6_0_io_outs_right[28] ,
    \ces_6_0_io_outs_right[27] ,
    \ces_6_0_io_outs_right[26] ,
    \ces_6_0_io_outs_right[25] ,
    \ces_6_0_io_outs_right[24] ,
    \ces_6_0_io_outs_right[23] ,
    \ces_6_0_io_outs_right[22] ,
    \ces_6_0_io_outs_right[21] ,
    \ces_6_0_io_outs_right[20] ,
    \ces_6_0_io_outs_right[19] ,
    \ces_6_0_io_outs_right[18] ,
    \ces_6_0_io_outs_right[17] ,
    \ces_6_0_io_outs_right[16] ,
    \ces_6_0_io_outs_right[15] ,
    \ces_6_0_io_outs_right[14] ,
    \ces_6_0_io_outs_right[13] ,
    \ces_6_0_io_outs_right[12] ,
    \ces_6_0_io_outs_right[11] ,
    \ces_6_0_io_outs_right[10] ,
    \ces_6_0_io_outs_right[9] ,
    \ces_6_0_io_outs_right[8] ,
    \ces_6_0_io_outs_right[7] ,
    \ces_6_0_io_outs_right[6] ,
    \ces_6_0_io_outs_right[5] ,
    \ces_6_0_io_outs_right[4] ,
    \ces_6_0_io_outs_right[3] ,
    \ces_6_0_io_outs_right[2] ,
    \ces_6_0_io_outs_right[1] ,
    \ces_6_0_io_outs_right[0] }),
    .io_ins_up({\ces_5_1_io_outs_up[63] ,
    \ces_5_1_io_outs_up[62] ,
    \ces_5_1_io_outs_up[61] ,
    \ces_5_1_io_outs_up[60] ,
    \ces_5_1_io_outs_up[59] ,
    \ces_5_1_io_outs_up[58] ,
    \ces_5_1_io_outs_up[57] ,
    \ces_5_1_io_outs_up[56] ,
    \ces_5_1_io_outs_up[55] ,
    \ces_5_1_io_outs_up[54] ,
    \ces_5_1_io_outs_up[53] ,
    \ces_5_1_io_outs_up[52] ,
    \ces_5_1_io_outs_up[51] ,
    \ces_5_1_io_outs_up[50] ,
    \ces_5_1_io_outs_up[49] ,
    \ces_5_1_io_outs_up[48] ,
    \ces_5_1_io_outs_up[47] ,
    \ces_5_1_io_outs_up[46] ,
    \ces_5_1_io_outs_up[45] ,
    \ces_5_1_io_outs_up[44] ,
    \ces_5_1_io_outs_up[43] ,
    \ces_5_1_io_outs_up[42] ,
    \ces_5_1_io_outs_up[41] ,
    \ces_5_1_io_outs_up[40] ,
    \ces_5_1_io_outs_up[39] ,
    \ces_5_1_io_outs_up[38] ,
    \ces_5_1_io_outs_up[37] ,
    \ces_5_1_io_outs_up[36] ,
    \ces_5_1_io_outs_up[35] ,
    \ces_5_1_io_outs_up[34] ,
    \ces_5_1_io_outs_up[33] ,
    \ces_5_1_io_outs_up[32] ,
    \ces_5_1_io_outs_up[31] ,
    \ces_5_1_io_outs_up[30] ,
    \ces_5_1_io_outs_up[29] ,
    \ces_5_1_io_outs_up[28] ,
    \ces_5_1_io_outs_up[27] ,
    \ces_5_1_io_outs_up[26] ,
    \ces_5_1_io_outs_up[25] ,
    \ces_5_1_io_outs_up[24] ,
    \ces_5_1_io_outs_up[23] ,
    \ces_5_1_io_outs_up[22] ,
    \ces_5_1_io_outs_up[21] ,
    \ces_5_1_io_outs_up[20] ,
    \ces_5_1_io_outs_up[19] ,
    \ces_5_1_io_outs_up[18] ,
    \ces_5_1_io_outs_up[17] ,
    \ces_5_1_io_outs_up[16] ,
    \ces_5_1_io_outs_up[15] ,
    \ces_5_1_io_outs_up[14] ,
    \ces_5_1_io_outs_up[13] ,
    \ces_5_1_io_outs_up[12] ,
    \ces_5_1_io_outs_up[11] ,
    \ces_5_1_io_outs_up[10] ,
    \ces_5_1_io_outs_up[9] ,
    \ces_5_1_io_outs_up[8] ,
    \ces_5_1_io_outs_up[7] ,
    \ces_5_1_io_outs_up[6] ,
    \ces_5_1_io_outs_up[5] ,
    \ces_5_1_io_outs_up[4] ,
    \ces_5_1_io_outs_up[3] ,
    \ces_5_1_io_outs_up[2] ,
    \ces_5_1_io_outs_up[1] ,
    \ces_5_1_io_outs_up[0] }),
    .io_outs_down({\ces_5_1_io_ins_down[63] ,
    \ces_5_1_io_ins_down[62] ,
    \ces_5_1_io_ins_down[61] ,
    \ces_5_1_io_ins_down[60] ,
    \ces_5_1_io_ins_down[59] ,
    \ces_5_1_io_ins_down[58] ,
    \ces_5_1_io_ins_down[57] ,
    \ces_5_1_io_ins_down[56] ,
    \ces_5_1_io_ins_down[55] ,
    \ces_5_1_io_ins_down[54] ,
    \ces_5_1_io_ins_down[53] ,
    \ces_5_1_io_ins_down[52] ,
    \ces_5_1_io_ins_down[51] ,
    \ces_5_1_io_ins_down[50] ,
    \ces_5_1_io_ins_down[49] ,
    \ces_5_1_io_ins_down[48] ,
    \ces_5_1_io_ins_down[47] ,
    \ces_5_1_io_ins_down[46] ,
    \ces_5_1_io_ins_down[45] ,
    \ces_5_1_io_ins_down[44] ,
    \ces_5_1_io_ins_down[43] ,
    \ces_5_1_io_ins_down[42] ,
    \ces_5_1_io_ins_down[41] ,
    \ces_5_1_io_ins_down[40] ,
    \ces_5_1_io_ins_down[39] ,
    \ces_5_1_io_ins_down[38] ,
    \ces_5_1_io_ins_down[37] ,
    \ces_5_1_io_ins_down[36] ,
    \ces_5_1_io_ins_down[35] ,
    \ces_5_1_io_ins_down[34] ,
    \ces_5_1_io_ins_down[33] ,
    \ces_5_1_io_ins_down[32] ,
    \ces_5_1_io_ins_down[31] ,
    \ces_5_1_io_ins_down[30] ,
    \ces_5_1_io_ins_down[29] ,
    \ces_5_1_io_ins_down[28] ,
    \ces_5_1_io_ins_down[27] ,
    \ces_5_1_io_ins_down[26] ,
    \ces_5_1_io_ins_down[25] ,
    \ces_5_1_io_ins_down[24] ,
    \ces_5_1_io_ins_down[23] ,
    \ces_5_1_io_ins_down[22] ,
    \ces_5_1_io_ins_down[21] ,
    \ces_5_1_io_ins_down[20] ,
    \ces_5_1_io_ins_down[19] ,
    \ces_5_1_io_ins_down[18] ,
    \ces_5_1_io_ins_down[17] ,
    \ces_5_1_io_ins_down[16] ,
    \ces_5_1_io_ins_down[15] ,
    \ces_5_1_io_ins_down[14] ,
    \ces_5_1_io_ins_down[13] ,
    \ces_5_1_io_ins_down[12] ,
    \ces_5_1_io_ins_down[11] ,
    \ces_5_1_io_ins_down[10] ,
    \ces_5_1_io_ins_down[9] ,
    \ces_5_1_io_ins_down[8] ,
    \ces_5_1_io_ins_down[7] ,
    \ces_5_1_io_ins_down[6] ,
    \ces_5_1_io_ins_down[5] ,
    \ces_5_1_io_ins_down[4] ,
    \ces_5_1_io_ins_down[3] ,
    \ces_5_1_io_ins_down[2] ,
    \ces_5_1_io_ins_down[1] ,
    \ces_5_1_io_ins_down[0] }),
    .io_outs_left({\ces_6_0_io_ins_left[63] ,
    \ces_6_0_io_ins_left[62] ,
    \ces_6_0_io_ins_left[61] ,
    \ces_6_0_io_ins_left[60] ,
    \ces_6_0_io_ins_left[59] ,
    \ces_6_0_io_ins_left[58] ,
    \ces_6_0_io_ins_left[57] ,
    \ces_6_0_io_ins_left[56] ,
    \ces_6_0_io_ins_left[55] ,
    \ces_6_0_io_ins_left[54] ,
    \ces_6_0_io_ins_left[53] ,
    \ces_6_0_io_ins_left[52] ,
    \ces_6_0_io_ins_left[51] ,
    \ces_6_0_io_ins_left[50] ,
    \ces_6_0_io_ins_left[49] ,
    \ces_6_0_io_ins_left[48] ,
    \ces_6_0_io_ins_left[47] ,
    \ces_6_0_io_ins_left[46] ,
    \ces_6_0_io_ins_left[45] ,
    \ces_6_0_io_ins_left[44] ,
    \ces_6_0_io_ins_left[43] ,
    \ces_6_0_io_ins_left[42] ,
    \ces_6_0_io_ins_left[41] ,
    \ces_6_0_io_ins_left[40] ,
    \ces_6_0_io_ins_left[39] ,
    \ces_6_0_io_ins_left[38] ,
    \ces_6_0_io_ins_left[37] ,
    \ces_6_0_io_ins_left[36] ,
    \ces_6_0_io_ins_left[35] ,
    \ces_6_0_io_ins_left[34] ,
    \ces_6_0_io_ins_left[33] ,
    \ces_6_0_io_ins_left[32] ,
    \ces_6_0_io_ins_left[31] ,
    \ces_6_0_io_ins_left[30] ,
    \ces_6_0_io_ins_left[29] ,
    \ces_6_0_io_ins_left[28] ,
    \ces_6_0_io_ins_left[27] ,
    \ces_6_0_io_ins_left[26] ,
    \ces_6_0_io_ins_left[25] ,
    \ces_6_0_io_ins_left[24] ,
    \ces_6_0_io_ins_left[23] ,
    \ces_6_0_io_ins_left[22] ,
    \ces_6_0_io_ins_left[21] ,
    \ces_6_0_io_ins_left[20] ,
    \ces_6_0_io_ins_left[19] ,
    \ces_6_0_io_ins_left[18] ,
    \ces_6_0_io_ins_left[17] ,
    \ces_6_0_io_ins_left[16] ,
    \ces_6_0_io_ins_left[15] ,
    \ces_6_0_io_ins_left[14] ,
    \ces_6_0_io_ins_left[13] ,
    \ces_6_0_io_ins_left[12] ,
    \ces_6_0_io_ins_left[11] ,
    \ces_6_0_io_ins_left[10] ,
    \ces_6_0_io_ins_left[9] ,
    \ces_6_0_io_ins_left[8] ,
    \ces_6_0_io_ins_left[7] ,
    \ces_6_0_io_ins_left[6] ,
    \ces_6_0_io_ins_left[5] ,
    \ces_6_0_io_ins_left[4] ,
    \ces_6_0_io_ins_left[3] ,
    \ces_6_0_io_ins_left[2] ,
    \ces_6_0_io_ins_left[1] ,
    \ces_6_0_io_ins_left[0] }),
    .io_outs_right({\ces_6_1_io_outs_right[63] ,
    \ces_6_1_io_outs_right[62] ,
    \ces_6_1_io_outs_right[61] ,
    \ces_6_1_io_outs_right[60] ,
    \ces_6_1_io_outs_right[59] ,
    \ces_6_1_io_outs_right[58] ,
    \ces_6_1_io_outs_right[57] ,
    \ces_6_1_io_outs_right[56] ,
    \ces_6_1_io_outs_right[55] ,
    \ces_6_1_io_outs_right[54] ,
    \ces_6_1_io_outs_right[53] ,
    \ces_6_1_io_outs_right[52] ,
    \ces_6_1_io_outs_right[51] ,
    \ces_6_1_io_outs_right[50] ,
    \ces_6_1_io_outs_right[49] ,
    \ces_6_1_io_outs_right[48] ,
    \ces_6_1_io_outs_right[47] ,
    \ces_6_1_io_outs_right[46] ,
    \ces_6_1_io_outs_right[45] ,
    \ces_6_1_io_outs_right[44] ,
    \ces_6_1_io_outs_right[43] ,
    \ces_6_1_io_outs_right[42] ,
    \ces_6_1_io_outs_right[41] ,
    \ces_6_1_io_outs_right[40] ,
    \ces_6_1_io_outs_right[39] ,
    \ces_6_1_io_outs_right[38] ,
    \ces_6_1_io_outs_right[37] ,
    \ces_6_1_io_outs_right[36] ,
    \ces_6_1_io_outs_right[35] ,
    \ces_6_1_io_outs_right[34] ,
    \ces_6_1_io_outs_right[33] ,
    \ces_6_1_io_outs_right[32] ,
    \ces_6_1_io_outs_right[31] ,
    \ces_6_1_io_outs_right[30] ,
    \ces_6_1_io_outs_right[29] ,
    \ces_6_1_io_outs_right[28] ,
    \ces_6_1_io_outs_right[27] ,
    \ces_6_1_io_outs_right[26] ,
    \ces_6_1_io_outs_right[25] ,
    \ces_6_1_io_outs_right[24] ,
    \ces_6_1_io_outs_right[23] ,
    \ces_6_1_io_outs_right[22] ,
    \ces_6_1_io_outs_right[21] ,
    \ces_6_1_io_outs_right[20] ,
    \ces_6_1_io_outs_right[19] ,
    \ces_6_1_io_outs_right[18] ,
    \ces_6_1_io_outs_right[17] ,
    \ces_6_1_io_outs_right[16] ,
    \ces_6_1_io_outs_right[15] ,
    \ces_6_1_io_outs_right[14] ,
    \ces_6_1_io_outs_right[13] ,
    \ces_6_1_io_outs_right[12] ,
    \ces_6_1_io_outs_right[11] ,
    \ces_6_1_io_outs_right[10] ,
    \ces_6_1_io_outs_right[9] ,
    \ces_6_1_io_outs_right[8] ,
    \ces_6_1_io_outs_right[7] ,
    \ces_6_1_io_outs_right[6] ,
    \ces_6_1_io_outs_right[5] ,
    \ces_6_1_io_outs_right[4] ,
    \ces_6_1_io_outs_right[3] ,
    \ces_6_1_io_outs_right[2] ,
    \ces_6_1_io_outs_right[1] ,
    \ces_6_1_io_outs_right[0] }),
    .io_outs_up({\ces_6_1_io_outs_up[63] ,
    \ces_6_1_io_outs_up[62] ,
    \ces_6_1_io_outs_up[61] ,
    \ces_6_1_io_outs_up[60] ,
    \ces_6_1_io_outs_up[59] ,
    \ces_6_1_io_outs_up[58] ,
    \ces_6_1_io_outs_up[57] ,
    \ces_6_1_io_outs_up[56] ,
    \ces_6_1_io_outs_up[55] ,
    \ces_6_1_io_outs_up[54] ,
    \ces_6_1_io_outs_up[53] ,
    \ces_6_1_io_outs_up[52] ,
    \ces_6_1_io_outs_up[51] ,
    \ces_6_1_io_outs_up[50] ,
    \ces_6_1_io_outs_up[49] ,
    \ces_6_1_io_outs_up[48] ,
    \ces_6_1_io_outs_up[47] ,
    \ces_6_1_io_outs_up[46] ,
    \ces_6_1_io_outs_up[45] ,
    \ces_6_1_io_outs_up[44] ,
    \ces_6_1_io_outs_up[43] ,
    \ces_6_1_io_outs_up[42] ,
    \ces_6_1_io_outs_up[41] ,
    \ces_6_1_io_outs_up[40] ,
    \ces_6_1_io_outs_up[39] ,
    \ces_6_1_io_outs_up[38] ,
    \ces_6_1_io_outs_up[37] ,
    \ces_6_1_io_outs_up[36] ,
    \ces_6_1_io_outs_up[35] ,
    \ces_6_1_io_outs_up[34] ,
    \ces_6_1_io_outs_up[33] ,
    \ces_6_1_io_outs_up[32] ,
    \ces_6_1_io_outs_up[31] ,
    \ces_6_1_io_outs_up[30] ,
    \ces_6_1_io_outs_up[29] ,
    \ces_6_1_io_outs_up[28] ,
    \ces_6_1_io_outs_up[27] ,
    \ces_6_1_io_outs_up[26] ,
    \ces_6_1_io_outs_up[25] ,
    \ces_6_1_io_outs_up[24] ,
    \ces_6_1_io_outs_up[23] ,
    \ces_6_1_io_outs_up[22] ,
    \ces_6_1_io_outs_up[21] ,
    \ces_6_1_io_outs_up[20] ,
    \ces_6_1_io_outs_up[19] ,
    \ces_6_1_io_outs_up[18] ,
    \ces_6_1_io_outs_up[17] ,
    \ces_6_1_io_outs_up[16] ,
    \ces_6_1_io_outs_up[15] ,
    \ces_6_1_io_outs_up[14] ,
    \ces_6_1_io_outs_up[13] ,
    \ces_6_1_io_outs_up[12] ,
    \ces_6_1_io_outs_up[11] ,
    \ces_6_1_io_outs_up[10] ,
    \ces_6_1_io_outs_up[9] ,
    \ces_6_1_io_outs_up[8] ,
    \ces_6_1_io_outs_up[7] ,
    \ces_6_1_io_outs_up[6] ,
    \ces_6_1_io_outs_up[5] ,
    \ces_6_1_io_outs_up[4] ,
    \ces_6_1_io_outs_up[3] ,
    \ces_6_1_io_outs_up[2] ,
    \ces_6_1_io_outs_up[1] ,
    \ces_6_1_io_outs_up[0] }));
 Element ces_6_2 (.clock(clknet_3_5_0_clock),
    .io_lsbIns_1(ces_6_1_io_lsbOuts_1),
    .io_lsbIns_2(ces_6_1_io_lsbOuts_2),
    .io_lsbIns_3(ces_6_1_io_lsbOuts_3),
    .io_lsbIns_4(ces_6_1_io_lsbOuts_4),
    .io_lsbIns_5(ces_6_1_io_lsbOuts_5),
    .io_lsbIns_6(ces_6_1_io_lsbOuts_6),
    .io_lsbIns_7(ces_6_1_io_lsbOuts_7),
    .io_lsbOuts_0(ces_6_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_2_io_lsbOuts_7),
    .io_ins_down({\ces_6_2_io_ins_down[63] ,
    \ces_6_2_io_ins_down[62] ,
    \ces_6_2_io_ins_down[61] ,
    \ces_6_2_io_ins_down[60] ,
    \ces_6_2_io_ins_down[59] ,
    \ces_6_2_io_ins_down[58] ,
    \ces_6_2_io_ins_down[57] ,
    \ces_6_2_io_ins_down[56] ,
    \ces_6_2_io_ins_down[55] ,
    \ces_6_2_io_ins_down[54] ,
    \ces_6_2_io_ins_down[53] ,
    \ces_6_2_io_ins_down[52] ,
    \ces_6_2_io_ins_down[51] ,
    \ces_6_2_io_ins_down[50] ,
    \ces_6_2_io_ins_down[49] ,
    \ces_6_2_io_ins_down[48] ,
    \ces_6_2_io_ins_down[47] ,
    \ces_6_2_io_ins_down[46] ,
    \ces_6_2_io_ins_down[45] ,
    \ces_6_2_io_ins_down[44] ,
    \ces_6_2_io_ins_down[43] ,
    \ces_6_2_io_ins_down[42] ,
    \ces_6_2_io_ins_down[41] ,
    \ces_6_2_io_ins_down[40] ,
    \ces_6_2_io_ins_down[39] ,
    \ces_6_2_io_ins_down[38] ,
    \ces_6_2_io_ins_down[37] ,
    \ces_6_2_io_ins_down[36] ,
    \ces_6_2_io_ins_down[35] ,
    \ces_6_2_io_ins_down[34] ,
    \ces_6_2_io_ins_down[33] ,
    \ces_6_2_io_ins_down[32] ,
    \ces_6_2_io_ins_down[31] ,
    \ces_6_2_io_ins_down[30] ,
    \ces_6_2_io_ins_down[29] ,
    \ces_6_2_io_ins_down[28] ,
    \ces_6_2_io_ins_down[27] ,
    \ces_6_2_io_ins_down[26] ,
    \ces_6_2_io_ins_down[25] ,
    \ces_6_2_io_ins_down[24] ,
    \ces_6_2_io_ins_down[23] ,
    \ces_6_2_io_ins_down[22] ,
    \ces_6_2_io_ins_down[21] ,
    \ces_6_2_io_ins_down[20] ,
    \ces_6_2_io_ins_down[19] ,
    \ces_6_2_io_ins_down[18] ,
    \ces_6_2_io_ins_down[17] ,
    \ces_6_2_io_ins_down[16] ,
    \ces_6_2_io_ins_down[15] ,
    \ces_6_2_io_ins_down[14] ,
    \ces_6_2_io_ins_down[13] ,
    \ces_6_2_io_ins_down[12] ,
    \ces_6_2_io_ins_down[11] ,
    \ces_6_2_io_ins_down[10] ,
    \ces_6_2_io_ins_down[9] ,
    \ces_6_2_io_ins_down[8] ,
    \ces_6_2_io_ins_down[7] ,
    \ces_6_2_io_ins_down[6] ,
    \ces_6_2_io_ins_down[5] ,
    \ces_6_2_io_ins_down[4] ,
    \ces_6_2_io_ins_down[3] ,
    \ces_6_2_io_ins_down[2] ,
    \ces_6_2_io_ins_down[1] ,
    \ces_6_2_io_ins_down[0] }),
    .io_ins_left({\ces_6_2_io_ins_left[63] ,
    \ces_6_2_io_ins_left[62] ,
    \ces_6_2_io_ins_left[61] ,
    \ces_6_2_io_ins_left[60] ,
    \ces_6_2_io_ins_left[59] ,
    \ces_6_2_io_ins_left[58] ,
    \ces_6_2_io_ins_left[57] ,
    \ces_6_2_io_ins_left[56] ,
    \ces_6_2_io_ins_left[55] ,
    \ces_6_2_io_ins_left[54] ,
    \ces_6_2_io_ins_left[53] ,
    \ces_6_2_io_ins_left[52] ,
    \ces_6_2_io_ins_left[51] ,
    \ces_6_2_io_ins_left[50] ,
    \ces_6_2_io_ins_left[49] ,
    \ces_6_2_io_ins_left[48] ,
    \ces_6_2_io_ins_left[47] ,
    \ces_6_2_io_ins_left[46] ,
    \ces_6_2_io_ins_left[45] ,
    \ces_6_2_io_ins_left[44] ,
    \ces_6_2_io_ins_left[43] ,
    \ces_6_2_io_ins_left[42] ,
    \ces_6_2_io_ins_left[41] ,
    \ces_6_2_io_ins_left[40] ,
    \ces_6_2_io_ins_left[39] ,
    \ces_6_2_io_ins_left[38] ,
    \ces_6_2_io_ins_left[37] ,
    \ces_6_2_io_ins_left[36] ,
    \ces_6_2_io_ins_left[35] ,
    \ces_6_2_io_ins_left[34] ,
    \ces_6_2_io_ins_left[33] ,
    \ces_6_2_io_ins_left[32] ,
    \ces_6_2_io_ins_left[31] ,
    \ces_6_2_io_ins_left[30] ,
    \ces_6_2_io_ins_left[29] ,
    \ces_6_2_io_ins_left[28] ,
    \ces_6_2_io_ins_left[27] ,
    \ces_6_2_io_ins_left[26] ,
    \ces_6_2_io_ins_left[25] ,
    \ces_6_2_io_ins_left[24] ,
    \ces_6_2_io_ins_left[23] ,
    \ces_6_2_io_ins_left[22] ,
    \ces_6_2_io_ins_left[21] ,
    \ces_6_2_io_ins_left[20] ,
    \ces_6_2_io_ins_left[19] ,
    \ces_6_2_io_ins_left[18] ,
    \ces_6_2_io_ins_left[17] ,
    \ces_6_2_io_ins_left[16] ,
    \ces_6_2_io_ins_left[15] ,
    \ces_6_2_io_ins_left[14] ,
    \ces_6_2_io_ins_left[13] ,
    \ces_6_2_io_ins_left[12] ,
    \ces_6_2_io_ins_left[11] ,
    \ces_6_2_io_ins_left[10] ,
    \ces_6_2_io_ins_left[9] ,
    \ces_6_2_io_ins_left[8] ,
    \ces_6_2_io_ins_left[7] ,
    \ces_6_2_io_ins_left[6] ,
    \ces_6_2_io_ins_left[5] ,
    \ces_6_2_io_ins_left[4] ,
    \ces_6_2_io_ins_left[3] ,
    \ces_6_2_io_ins_left[2] ,
    \ces_6_2_io_ins_left[1] ,
    \ces_6_2_io_ins_left[0] }),
    .io_ins_right({\ces_6_1_io_outs_right[63] ,
    \ces_6_1_io_outs_right[62] ,
    \ces_6_1_io_outs_right[61] ,
    \ces_6_1_io_outs_right[60] ,
    \ces_6_1_io_outs_right[59] ,
    \ces_6_1_io_outs_right[58] ,
    \ces_6_1_io_outs_right[57] ,
    \ces_6_1_io_outs_right[56] ,
    \ces_6_1_io_outs_right[55] ,
    \ces_6_1_io_outs_right[54] ,
    \ces_6_1_io_outs_right[53] ,
    \ces_6_1_io_outs_right[52] ,
    \ces_6_1_io_outs_right[51] ,
    \ces_6_1_io_outs_right[50] ,
    \ces_6_1_io_outs_right[49] ,
    \ces_6_1_io_outs_right[48] ,
    \ces_6_1_io_outs_right[47] ,
    \ces_6_1_io_outs_right[46] ,
    \ces_6_1_io_outs_right[45] ,
    \ces_6_1_io_outs_right[44] ,
    \ces_6_1_io_outs_right[43] ,
    \ces_6_1_io_outs_right[42] ,
    \ces_6_1_io_outs_right[41] ,
    \ces_6_1_io_outs_right[40] ,
    \ces_6_1_io_outs_right[39] ,
    \ces_6_1_io_outs_right[38] ,
    \ces_6_1_io_outs_right[37] ,
    \ces_6_1_io_outs_right[36] ,
    \ces_6_1_io_outs_right[35] ,
    \ces_6_1_io_outs_right[34] ,
    \ces_6_1_io_outs_right[33] ,
    \ces_6_1_io_outs_right[32] ,
    \ces_6_1_io_outs_right[31] ,
    \ces_6_1_io_outs_right[30] ,
    \ces_6_1_io_outs_right[29] ,
    \ces_6_1_io_outs_right[28] ,
    \ces_6_1_io_outs_right[27] ,
    \ces_6_1_io_outs_right[26] ,
    \ces_6_1_io_outs_right[25] ,
    \ces_6_1_io_outs_right[24] ,
    \ces_6_1_io_outs_right[23] ,
    \ces_6_1_io_outs_right[22] ,
    \ces_6_1_io_outs_right[21] ,
    \ces_6_1_io_outs_right[20] ,
    \ces_6_1_io_outs_right[19] ,
    \ces_6_1_io_outs_right[18] ,
    \ces_6_1_io_outs_right[17] ,
    \ces_6_1_io_outs_right[16] ,
    \ces_6_1_io_outs_right[15] ,
    \ces_6_1_io_outs_right[14] ,
    \ces_6_1_io_outs_right[13] ,
    \ces_6_1_io_outs_right[12] ,
    \ces_6_1_io_outs_right[11] ,
    \ces_6_1_io_outs_right[10] ,
    \ces_6_1_io_outs_right[9] ,
    \ces_6_1_io_outs_right[8] ,
    \ces_6_1_io_outs_right[7] ,
    \ces_6_1_io_outs_right[6] ,
    \ces_6_1_io_outs_right[5] ,
    \ces_6_1_io_outs_right[4] ,
    \ces_6_1_io_outs_right[3] ,
    \ces_6_1_io_outs_right[2] ,
    \ces_6_1_io_outs_right[1] ,
    \ces_6_1_io_outs_right[0] }),
    .io_ins_up({\ces_5_2_io_outs_up[63] ,
    \ces_5_2_io_outs_up[62] ,
    \ces_5_2_io_outs_up[61] ,
    \ces_5_2_io_outs_up[60] ,
    \ces_5_2_io_outs_up[59] ,
    \ces_5_2_io_outs_up[58] ,
    \ces_5_2_io_outs_up[57] ,
    \ces_5_2_io_outs_up[56] ,
    \ces_5_2_io_outs_up[55] ,
    \ces_5_2_io_outs_up[54] ,
    \ces_5_2_io_outs_up[53] ,
    \ces_5_2_io_outs_up[52] ,
    \ces_5_2_io_outs_up[51] ,
    \ces_5_2_io_outs_up[50] ,
    \ces_5_2_io_outs_up[49] ,
    \ces_5_2_io_outs_up[48] ,
    \ces_5_2_io_outs_up[47] ,
    \ces_5_2_io_outs_up[46] ,
    \ces_5_2_io_outs_up[45] ,
    \ces_5_2_io_outs_up[44] ,
    \ces_5_2_io_outs_up[43] ,
    \ces_5_2_io_outs_up[42] ,
    \ces_5_2_io_outs_up[41] ,
    \ces_5_2_io_outs_up[40] ,
    \ces_5_2_io_outs_up[39] ,
    \ces_5_2_io_outs_up[38] ,
    \ces_5_2_io_outs_up[37] ,
    \ces_5_2_io_outs_up[36] ,
    \ces_5_2_io_outs_up[35] ,
    \ces_5_2_io_outs_up[34] ,
    \ces_5_2_io_outs_up[33] ,
    \ces_5_2_io_outs_up[32] ,
    \ces_5_2_io_outs_up[31] ,
    \ces_5_2_io_outs_up[30] ,
    \ces_5_2_io_outs_up[29] ,
    \ces_5_2_io_outs_up[28] ,
    \ces_5_2_io_outs_up[27] ,
    \ces_5_2_io_outs_up[26] ,
    \ces_5_2_io_outs_up[25] ,
    \ces_5_2_io_outs_up[24] ,
    \ces_5_2_io_outs_up[23] ,
    \ces_5_2_io_outs_up[22] ,
    \ces_5_2_io_outs_up[21] ,
    \ces_5_2_io_outs_up[20] ,
    \ces_5_2_io_outs_up[19] ,
    \ces_5_2_io_outs_up[18] ,
    \ces_5_2_io_outs_up[17] ,
    \ces_5_2_io_outs_up[16] ,
    \ces_5_2_io_outs_up[15] ,
    \ces_5_2_io_outs_up[14] ,
    \ces_5_2_io_outs_up[13] ,
    \ces_5_2_io_outs_up[12] ,
    \ces_5_2_io_outs_up[11] ,
    \ces_5_2_io_outs_up[10] ,
    \ces_5_2_io_outs_up[9] ,
    \ces_5_2_io_outs_up[8] ,
    \ces_5_2_io_outs_up[7] ,
    \ces_5_2_io_outs_up[6] ,
    \ces_5_2_io_outs_up[5] ,
    \ces_5_2_io_outs_up[4] ,
    \ces_5_2_io_outs_up[3] ,
    \ces_5_2_io_outs_up[2] ,
    \ces_5_2_io_outs_up[1] ,
    \ces_5_2_io_outs_up[0] }),
    .io_outs_down({\ces_5_2_io_ins_down[63] ,
    \ces_5_2_io_ins_down[62] ,
    \ces_5_2_io_ins_down[61] ,
    \ces_5_2_io_ins_down[60] ,
    \ces_5_2_io_ins_down[59] ,
    \ces_5_2_io_ins_down[58] ,
    \ces_5_2_io_ins_down[57] ,
    \ces_5_2_io_ins_down[56] ,
    \ces_5_2_io_ins_down[55] ,
    \ces_5_2_io_ins_down[54] ,
    \ces_5_2_io_ins_down[53] ,
    \ces_5_2_io_ins_down[52] ,
    \ces_5_2_io_ins_down[51] ,
    \ces_5_2_io_ins_down[50] ,
    \ces_5_2_io_ins_down[49] ,
    \ces_5_2_io_ins_down[48] ,
    \ces_5_2_io_ins_down[47] ,
    \ces_5_2_io_ins_down[46] ,
    \ces_5_2_io_ins_down[45] ,
    \ces_5_2_io_ins_down[44] ,
    \ces_5_2_io_ins_down[43] ,
    \ces_5_2_io_ins_down[42] ,
    \ces_5_2_io_ins_down[41] ,
    \ces_5_2_io_ins_down[40] ,
    \ces_5_2_io_ins_down[39] ,
    \ces_5_2_io_ins_down[38] ,
    \ces_5_2_io_ins_down[37] ,
    \ces_5_2_io_ins_down[36] ,
    \ces_5_2_io_ins_down[35] ,
    \ces_5_2_io_ins_down[34] ,
    \ces_5_2_io_ins_down[33] ,
    \ces_5_2_io_ins_down[32] ,
    \ces_5_2_io_ins_down[31] ,
    \ces_5_2_io_ins_down[30] ,
    \ces_5_2_io_ins_down[29] ,
    \ces_5_2_io_ins_down[28] ,
    \ces_5_2_io_ins_down[27] ,
    \ces_5_2_io_ins_down[26] ,
    \ces_5_2_io_ins_down[25] ,
    \ces_5_2_io_ins_down[24] ,
    \ces_5_2_io_ins_down[23] ,
    \ces_5_2_io_ins_down[22] ,
    \ces_5_2_io_ins_down[21] ,
    \ces_5_2_io_ins_down[20] ,
    \ces_5_2_io_ins_down[19] ,
    \ces_5_2_io_ins_down[18] ,
    \ces_5_2_io_ins_down[17] ,
    \ces_5_2_io_ins_down[16] ,
    \ces_5_2_io_ins_down[15] ,
    \ces_5_2_io_ins_down[14] ,
    \ces_5_2_io_ins_down[13] ,
    \ces_5_2_io_ins_down[12] ,
    \ces_5_2_io_ins_down[11] ,
    \ces_5_2_io_ins_down[10] ,
    \ces_5_2_io_ins_down[9] ,
    \ces_5_2_io_ins_down[8] ,
    \ces_5_2_io_ins_down[7] ,
    \ces_5_2_io_ins_down[6] ,
    \ces_5_2_io_ins_down[5] ,
    \ces_5_2_io_ins_down[4] ,
    \ces_5_2_io_ins_down[3] ,
    \ces_5_2_io_ins_down[2] ,
    \ces_5_2_io_ins_down[1] ,
    \ces_5_2_io_ins_down[0] }),
    .io_outs_left({\ces_6_1_io_ins_left[63] ,
    \ces_6_1_io_ins_left[62] ,
    \ces_6_1_io_ins_left[61] ,
    \ces_6_1_io_ins_left[60] ,
    \ces_6_1_io_ins_left[59] ,
    \ces_6_1_io_ins_left[58] ,
    \ces_6_1_io_ins_left[57] ,
    \ces_6_1_io_ins_left[56] ,
    \ces_6_1_io_ins_left[55] ,
    \ces_6_1_io_ins_left[54] ,
    \ces_6_1_io_ins_left[53] ,
    \ces_6_1_io_ins_left[52] ,
    \ces_6_1_io_ins_left[51] ,
    \ces_6_1_io_ins_left[50] ,
    \ces_6_1_io_ins_left[49] ,
    \ces_6_1_io_ins_left[48] ,
    \ces_6_1_io_ins_left[47] ,
    \ces_6_1_io_ins_left[46] ,
    \ces_6_1_io_ins_left[45] ,
    \ces_6_1_io_ins_left[44] ,
    \ces_6_1_io_ins_left[43] ,
    \ces_6_1_io_ins_left[42] ,
    \ces_6_1_io_ins_left[41] ,
    \ces_6_1_io_ins_left[40] ,
    \ces_6_1_io_ins_left[39] ,
    \ces_6_1_io_ins_left[38] ,
    \ces_6_1_io_ins_left[37] ,
    \ces_6_1_io_ins_left[36] ,
    \ces_6_1_io_ins_left[35] ,
    \ces_6_1_io_ins_left[34] ,
    \ces_6_1_io_ins_left[33] ,
    \ces_6_1_io_ins_left[32] ,
    \ces_6_1_io_ins_left[31] ,
    \ces_6_1_io_ins_left[30] ,
    \ces_6_1_io_ins_left[29] ,
    \ces_6_1_io_ins_left[28] ,
    \ces_6_1_io_ins_left[27] ,
    \ces_6_1_io_ins_left[26] ,
    \ces_6_1_io_ins_left[25] ,
    \ces_6_1_io_ins_left[24] ,
    \ces_6_1_io_ins_left[23] ,
    \ces_6_1_io_ins_left[22] ,
    \ces_6_1_io_ins_left[21] ,
    \ces_6_1_io_ins_left[20] ,
    \ces_6_1_io_ins_left[19] ,
    \ces_6_1_io_ins_left[18] ,
    \ces_6_1_io_ins_left[17] ,
    \ces_6_1_io_ins_left[16] ,
    \ces_6_1_io_ins_left[15] ,
    \ces_6_1_io_ins_left[14] ,
    \ces_6_1_io_ins_left[13] ,
    \ces_6_1_io_ins_left[12] ,
    \ces_6_1_io_ins_left[11] ,
    \ces_6_1_io_ins_left[10] ,
    \ces_6_1_io_ins_left[9] ,
    \ces_6_1_io_ins_left[8] ,
    \ces_6_1_io_ins_left[7] ,
    \ces_6_1_io_ins_left[6] ,
    \ces_6_1_io_ins_left[5] ,
    \ces_6_1_io_ins_left[4] ,
    \ces_6_1_io_ins_left[3] ,
    \ces_6_1_io_ins_left[2] ,
    \ces_6_1_io_ins_left[1] ,
    \ces_6_1_io_ins_left[0] }),
    .io_outs_right({\ces_6_2_io_outs_right[63] ,
    \ces_6_2_io_outs_right[62] ,
    \ces_6_2_io_outs_right[61] ,
    \ces_6_2_io_outs_right[60] ,
    \ces_6_2_io_outs_right[59] ,
    \ces_6_2_io_outs_right[58] ,
    \ces_6_2_io_outs_right[57] ,
    \ces_6_2_io_outs_right[56] ,
    \ces_6_2_io_outs_right[55] ,
    \ces_6_2_io_outs_right[54] ,
    \ces_6_2_io_outs_right[53] ,
    \ces_6_2_io_outs_right[52] ,
    \ces_6_2_io_outs_right[51] ,
    \ces_6_2_io_outs_right[50] ,
    \ces_6_2_io_outs_right[49] ,
    \ces_6_2_io_outs_right[48] ,
    \ces_6_2_io_outs_right[47] ,
    \ces_6_2_io_outs_right[46] ,
    \ces_6_2_io_outs_right[45] ,
    \ces_6_2_io_outs_right[44] ,
    \ces_6_2_io_outs_right[43] ,
    \ces_6_2_io_outs_right[42] ,
    \ces_6_2_io_outs_right[41] ,
    \ces_6_2_io_outs_right[40] ,
    \ces_6_2_io_outs_right[39] ,
    \ces_6_2_io_outs_right[38] ,
    \ces_6_2_io_outs_right[37] ,
    \ces_6_2_io_outs_right[36] ,
    \ces_6_2_io_outs_right[35] ,
    \ces_6_2_io_outs_right[34] ,
    \ces_6_2_io_outs_right[33] ,
    \ces_6_2_io_outs_right[32] ,
    \ces_6_2_io_outs_right[31] ,
    \ces_6_2_io_outs_right[30] ,
    \ces_6_2_io_outs_right[29] ,
    \ces_6_2_io_outs_right[28] ,
    \ces_6_2_io_outs_right[27] ,
    \ces_6_2_io_outs_right[26] ,
    \ces_6_2_io_outs_right[25] ,
    \ces_6_2_io_outs_right[24] ,
    \ces_6_2_io_outs_right[23] ,
    \ces_6_2_io_outs_right[22] ,
    \ces_6_2_io_outs_right[21] ,
    \ces_6_2_io_outs_right[20] ,
    \ces_6_2_io_outs_right[19] ,
    \ces_6_2_io_outs_right[18] ,
    \ces_6_2_io_outs_right[17] ,
    \ces_6_2_io_outs_right[16] ,
    \ces_6_2_io_outs_right[15] ,
    \ces_6_2_io_outs_right[14] ,
    \ces_6_2_io_outs_right[13] ,
    \ces_6_2_io_outs_right[12] ,
    \ces_6_2_io_outs_right[11] ,
    \ces_6_2_io_outs_right[10] ,
    \ces_6_2_io_outs_right[9] ,
    \ces_6_2_io_outs_right[8] ,
    \ces_6_2_io_outs_right[7] ,
    \ces_6_2_io_outs_right[6] ,
    \ces_6_2_io_outs_right[5] ,
    \ces_6_2_io_outs_right[4] ,
    \ces_6_2_io_outs_right[3] ,
    \ces_6_2_io_outs_right[2] ,
    \ces_6_2_io_outs_right[1] ,
    \ces_6_2_io_outs_right[0] }),
    .io_outs_up({\ces_6_2_io_outs_up[63] ,
    \ces_6_2_io_outs_up[62] ,
    \ces_6_2_io_outs_up[61] ,
    \ces_6_2_io_outs_up[60] ,
    \ces_6_2_io_outs_up[59] ,
    \ces_6_2_io_outs_up[58] ,
    \ces_6_2_io_outs_up[57] ,
    \ces_6_2_io_outs_up[56] ,
    \ces_6_2_io_outs_up[55] ,
    \ces_6_2_io_outs_up[54] ,
    \ces_6_2_io_outs_up[53] ,
    \ces_6_2_io_outs_up[52] ,
    \ces_6_2_io_outs_up[51] ,
    \ces_6_2_io_outs_up[50] ,
    \ces_6_2_io_outs_up[49] ,
    \ces_6_2_io_outs_up[48] ,
    \ces_6_2_io_outs_up[47] ,
    \ces_6_2_io_outs_up[46] ,
    \ces_6_2_io_outs_up[45] ,
    \ces_6_2_io_outs_up[44] ,
    \ces_6_2_io_outs_up[43] ,
    \ces_6_2_io_outs_up[42] ,
    \ces_6_2_io_outs_up[41] ,
    \ces_6_2_io_outs_up[40] ,
    \ces_6_2_io_outs_up[39] ,
    \ces_6_2_io_outs_up[38] ,
    \ces_6_2_io_outs_up[37] ,
    \ces_6_2_io_outs_up[36] ,
    \ces_6_2_io_outs_up[35] ,
    \ces_6_2_io_outs_up[34] ,
    \ces_6_2_io_outs_up[33] ,
    \ces_6_2_io_outs_up[32] ,
    \ces_6_2_io_outs_up[31] ,
    \ces_6_2_io_outs_up[30] ,
    \ces_6_2_io_outs_up[29] ,
    \ces_6_2_io_outs_up[28] ,
    \ces_6_2_io_outs_up[27] ,
    \ces_6_2_io_outs_up[26] ,
    \ces_6_2_io_outs_up[25] ,
    \ces_6_2_io_outs_up[24] ,
    \ces_6_2_io_outs_up[23] ,
    \ces_6_2_io_outs_up[22] ,
    \ces_6_2_io_outs_up[21] ,
    \ces_6_2_io_outs_up[20] ,
    \ces_6_2_io_outs_up[19] ,
    \ces_6_2_io_outs_up[18] ,
    \ces_6_2_io_outs_up[17] ,
    \ces_6_2_io_outs_up[16] ,
    \ces_6_2_io_outs_up[15] ,
    \ces_6_2_io_outs_up[14] ,
    \ces_6_2_io_outs_up[13] ,
    \ces_6_2_io_outs_up[12] ,
    \ces_6_2_io_outs_up[11] ,
    \ces_6_2_io_outs_up[10] ,
    \ces_6_2_io_outs_up[9] ,
    \ces_6_2_io_outs_up[8] ,
    \ces_6_2_io_outs_up[7] ,
    \ces_6_2_io_outs_up[6] ,
    \ces_6_2_io_outs_up[5] ,
    \ces_6_2_io_outs_up[4] ,
    \ces_6_2_io_outs_up[3] ,
    \ces_6_2_io_outs_up[2] ,
    \ces_6_2_io_outs_up[1] ,
    \ces_6_2_io_outs_up[0] }));
 Element ces_6_3 (.clock(clknet_3_5_0_clock),
    .io_lsbIns_1(ces_6_2_io_lsbOuts_1),
    .io_lsbIns_2(ces_6_2_io_lsbOuts_2),
    .io_lsbIns_3(ces_6_2_io_lsbOuts_3),
    .io_lsbIns_4(ces_6_2_io_lsbOuts_4),
    .io_lsbIns_5(ces_6_2_io_lsbOuts_5),
    .io_lsbIns_6(ces_6_2_io_lsbOuts_6),
    .io_lsbIns_7(ces_6_2_io_lsbOuts_7),
    .io_lsbOuts_0(ces_6_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_3_io_lsbOuts_7),
    .io_ins_down({\ces_6_3_io_ins_down[63] ,
    \ces_6_3_io_ins_down[62] ,
    \ces_6_3_io_ins_down[61] ,
    \ces_6_3_io_ins_down[60] ,
    \ces_6_3_io_ins_down[59] ,
    \ces_6_3_io_ins_down[58] ,
    \ces_6_3_io_ins_down[57] ,
    \ces_6_3_io_ins_down[56] ,
    \ces_6_3_io_ins_down[55] ,
    \ces_6_3_io_ins_down[54] ,
    \ces_6_3_io_ins_down[53] ,
    \ces_6_3_io_ins_down[52] ,
    \ces_6_3_io_ins_down[51] ,
    \ces_6_3_io_ins_down[50] ,
    \ces_6_3_io_ins_down[49] ,
    \ces_6_3_io_ins_down[48] ,
    \ces_6_3_io_ins_down[47] ,
    \ces_6_3_io_ins_down[46] ,
    \ces_6_3_io_ins_down[45] ,
    \ces_6_3_io_ins_down[44] ,
    \ces_6_3_io_ins_down[43] ,
    \ces_6_3_io_ins_down[42] ,
    \ces_6_3_io_ins_down[41] ,
    \ces_6_3_io_ins_down[40] ,
    \ces_6_3_io_ins_down[39] ,
    \ces_6_3_io_ins_down[38] ,
    \ces_6_3_io_ins_down[37] ,
    \ces_6_3_io_ins_down[36] ,
    \ces_6_3_io_ins_down[35] ,
    \ces_6_3_io_ins_down[34] ,
    \ces_6_3_io_ins_down[33] ,
    \ces_6_3_io_ins_down[32] ,
    \ces_6_3_io_ins_down[31] ,
    \ces_6_3_io_ins_down[30] ,
    \ces_6_3_io_ins_down[29] ,
    \ces_6_3_io_ins_down[28] ,
    \ces_6_3_io_ins_down[27] ,
    \ces_6_3_io_ins_down[26] ,
    \ces_6_3_io_ins_down[25] ,
    \ces_6_3_io_ins_down[24] ,
    \ces_6_3_io_ins_down[23] ,
    \ces_6_3_io_ins_down[22] ,
    \ces_6_3_io_ins_down[21] ,
    \ces_6_3_io_ins_down[20] ,
    \ces_6_3_io_ins_down[19] ,
    \ces_6_3_io_ins_down[18] ,
    \ces_6_3_io_ins_down[17] ,
    \ces_6_3_io_ins_down[16] ,
    \ces_6_3_io_ins_down[15] ,
    \ces_6_3_io_ins_down[14] ,
    \ces_6_3_io_ins_down[13] ,
    \ces_6_3_io_ins_down[12] ,
    \ces_6_3_io_ins_down[11] ,
    \ces_6_3_io_ins_down[10] ,
    \ces_6_3_io_ins_down[9] ,
    \ces_6_3_io_ins_down[8] ,
    \ces_6_3_io_ins_down[7] ,
    \ces_6_3_io_ins_down[6] ,
    \ces_6_3_io_ins_down[5] ,
    \ces_6_3_io_ins_down[4] ,
    \ces_6_3_io_ins_down[3] ,
    \ces_6_3_io_ins_down[2] ,
    \ces_6_3_io_ins_down[1] ,
    \ces_6_3_io_ins_down[0] }),
    .io_ins_left({\ces_6_3_io_ins_left[63] ,
    \ces_6_3_io_ins_left[62] ,
    \ces_6_3_io_ins_left[61] ,
    \ces_6_3_io_ins_left[60] ,
    \ces_6_3_io_ins_left[59] ,
    \ces_6_3_io_ins_left[58] ,
    \ces_6_3_io_ins_left[57] ,
    \ces_6_3_io_ins_left[56] ,
    \ces_6_3_io_ins_left[55] ,
    \ces_6_3_io_ins_left[54] ,
    \ces_6_3_io_ins_left[53] ,
    \ces_6_3_io_ins_left[52] ,
    \ces_6_3_io_ins_left[51] ,
    \ces_6_3_io_ins_left[50] ,
    \ces_6_3_io_ins_left[49] ,
    \ces_6_3_io_ins_left[48] ,
    \ces_6_3_io_ins_left[47] ,
    \ces_6_3_io_ins_left[46] ,
    \ces_6_3_io_ins_left[45] ,
    \ces_6_3_io_ins_left[44] ,
    \ces_6_3_io_ins_left[43] ,
    \ces_6_3_io_ins_left[42] ,
    \ces_6_3_io_ins_left[41] ,
    \ces_6_3_io_ins_left[40] ,
    \ces_6_3_io_ins_left[39] ,
    \ces_6_3_io_ins_left[38] ,
    \ces_6_3_io_ins_left[37] ,
    \ces_6_3_io_ins_left[36] ,
    \ces_6_3_io_ins_left[35] ,
    \ces_6_3_io_ins_left[34] ,
    \ces_6_3_io_ins_left[33] ,
    \ces_6_3_io_ins_left[32] ,
    \ces_6_3_io_ins_left[31] ,
    \ces_6_3_io_ins_left[30] ,
    \ces_6_3_io_ins_left[29] ,
    \ces_6_3_io_ins_left[28] ,
    \ces_6_3_io_ins_left[27] ,
    \ces_6_3_io_ins_left[26] ,
    \ces_6_3_io_ins_left[25] ,
    \ces_6_3_io_ins_left[24] ,
    \ces_6_3_io_ins_left[23] ,
    \ces_6_3_io_ins_left[22] ,
    \ces_6_3_io_ins_left[21] ,
    \ces_6_3_io_ins_left[20] ,
    \ces_6_3_io_ins_left[19] ,
    \ces_6_3_io_ins_left[18] ,
    \ces_6_3_io_ins_left[17] ,
    \ces_6_3_io_ins_left[16] ,
    \ces_6_3_io_ins_left[15] ,
    \ces_6_3_io_ins_left[14] ,
    \ces_6_3_io_ins_left[13] ,
    \ces_6_3_io_ins_left[12] ,
    \ces_6_3_io_ins_left[11] ,
    \ces_6_3_io_ins_left[10] ,
    \ces_6_3_io_ins_left[9] ,
    \ces_6_3_io_ins_left[8] ,
    \ces_6_3_io_ins_left[7] ,
    \ces_6_3_io_ins_left[6] ,
    \ces_6_3_io_ins_left[5] ,
    \ces_6_3_io_ins_left[4] ,
    \ces_6_3_io_ins_left[3] ,
    \ces_6_3_io_ins_left[2] ,
    \ces_6_3_io_ins_left[1] ,
    \ces_6_3_io_ins_left[0] }),
    .io_ins_right({\ces_6_2_io_outs_right[63] ,
    \ces_6_2_io_outs_right[62] ,
    \ces_6_2_io_outs_right[61] ,
    \ces_6_2_io_outs_right[60] ,
    \ces_6_2_io_outs_right[59] ,
    \ces_6_2_io_outs_right[58] ,
    \ces_6_2_io_outs_right[57] ,
    \ces_6_2_io_outs_right[56] ,
    \ces_6_2_io_outs_right[55] ,
    \ces_6_2_io_outs_right[54] ,
    \ces_6_2_io_outs_right[53] ,
    \ces_6_2_io_outs_right[52] ,
    \ces_6_2_io_outs_right[51] ,
    \ces_6_2_io_outs_right[50] ,
    \ces_6_2_io_outs_right[49] ,
    \ces_6_2_io_outs_right[48] ,
    \ces_6_2_io_outs_right[47] ,
    \ces_6_2_io_outs_right[46] ,
    \ces_6_2_io_outs_right[45] ,
    \ces_6_2_io_outs_right[44] ,
    \ces_6_2_io_outs_right[43] ,
    \ces_6_2_io_outs_right[42] ,
    \ces_6_2_io_outs_right[41] ,
    \ces_6_2_io_outs_right[40] ,
    \ces_6_2_io_outs_right[39] ,
    \ces_6_2_io_outs_right[38] ,
    \ces_6_2_io_outs_right[37] ,
    \ces_6_2_io_outs_right[36] ,
    \ces_6_2_io_outs_right[35] ,
    \ces_6_2_io_outs_right[34] ,
    \ces_6_2_io_outs_right[33] ,
    \ces_6_2_io_outs_right[32] ,
    \ces_6_2_io_outs_right[31] ,
    \ces_6_2_io_outs_right[30] ,
    \ces_6_2_io_outs_right[29] ,
    \ces_6_2_io_outs_right[28] ,
    \ces_6_2_io_outs_right[27] ,
    \ces_6_2_io_outs_right[26] ,
    \ces_6_2_io_outs_right[25] ,
    \ces_6_2_io_outs_right[24] ,
    \ces_6_2_io_outs_right[23] ,
    \ces_6_2_io_outs_right[22] ,
    \ces_6_2_io_outs_right[21] ,
    \ces_6_2_io_outs_right[20] ,
    \ces_6_2_io_outs_right[19] ,
    \ces_6_2_io_outs_right[18] ,
    \ces_6_2_io_outs_right[17] ,
    \ces_6_2_io_outs_right[16] ,
    \ces_6_2_io_outs_right[15] ,
    \ces_6_2_io_outs_right[14] ,
    \ces_6_2_io_outs_right[13] ,
    \ces_6_2_io_outs_right[12] ,
    \ces_6_2_io_outs_right[11] ,
    \ces_6_2_io_outs_right[10] ,
    \ces_6_2_io_outs_right[9] ,
    \ces_6_2_io_outs_right[8] ,
    \ces_6_2_io_outs_right[7] ,
    \ces_6_2_io_outs_right[6] ,
    \ces_6_2_io_outs_right[5] ,
    \ces_6_2_io_outs_right[4] ,
    \ces_6_2_io_outs_right[3] ,
    \ces_6_2_io_outs_right[2] ,
    \ces_6_2_io_outs_right[1] ,
    \ces_6_2_io_outs_right[0] }),
    .io_ins_up({\ces_5_3_io_outs_up[63] ,
    \ces_5_3_io_outs_up[62] ,
    \ces_5_3_io_outs_up[61] ,
    \ces_5_3_io_outs_up[60] ,
    \ces_5_3_io_outs_up[59] ,
    \ces_5_3_io_outs_up[58] ,
    \ces_5_3_io_outs_up[57] ,
    \ces_5_3_io_outs_up[56] ,
    \ces_5_3_io_outs_up[55] ,
    \ces_5_3_io_outs_up[54] ,
    \ces_5_3_io_outs_up[53] ,
    \ces_5_3_io_outs_up[52] ,
    \ces_5_3_io_outs_up[51] ,
    \ces_5_3_io_outs_up[50] ,
    \ces_5_3_io_outs_up[49] ,
    \ces_5_3_io_outs_up[48] ,
    \ces_5_3_io_outs_up[47] ,
    \ces_5_3_io_outs_up[46] ,
    \ces_5_3_io_outs_up[45] ,
    \ces_5_3_io_outs_up[44] ,
    \ces_5_3_io_outs_up[43] ,
    \ces_5_3_io_outs_up[42] ,
    \ces_5_3_io_outs_up[41] ,
    \ces_5_3_io_outs_up[40] ,
    \ces_5_3_io_outs_up[39] ,
    \ces_5_3_io_outs_up[38] ,
    \ces_5_3_io_outs_up[37] ,
    \ces_5_3_io_outs_up[36] ,
    \ces_5_3_io_outs_up[35] ,
    \ces_5_3_io_outs_up[34] ,
    \ces_5_3_io_outs_up[33] ,
    \ces_5_3_io_outs_up[32] ,
    \ces_5_3_io_outs_up[31] ,
    \ces_5_3_io_outs_up[30] ,
    \ces_5_3_io_outs_up[29] ,
    \ces_5_3_io_outs_up[28] ,
    \ces_5_3_io_outs_up[27] ,
    \ces_5_3_io_outs_up[26] ,
    \ces_5_3_io_outs_up[25] ,
    \ces_5_3_io_outs_up[24] ,
    \ces_5_3_io_outs_up[23] ,
    \ces_5_3_io_outs_up[22] ,
    \ces_5_3_io_outs_up[21] ,
    \ces_5_3_io_outs_up[20] ,
    \ces_5_3_io_outs_up[19] ,
    \ces_5_3_io_outs_up[18] ,
    \ces_5_3_io_outs_up[17] ,
    \ces_5_3_io_outs_up[16] ,
    \ces_5_3_io_outs_up[15] ,
    \ces_5_3_io_outs_up[14] ,
    \ces_5_3_io_outs_up[13] ,
    \ces_5_3_io_outs_up[12] ,
    \ces_5_3_io_outs_up[11] ,
    \ces_5_3_io_outs_up[10] ,
    \ces_5_3_io_outs_up[9] ,
    \ces_5_3_io_outs_up[8] ,
    \ces_5_3_io_outs_up[7] ,
    \ces_5_3_io_outs_up[6] ,
    \ces_5_3_io_outs_up[5] ,
    \ces_5_3_io_outs_up[4] ,
    \ces_5_3_io_outs_up[3] ,
    \ces_5_3_io_outs_up[2] ,
    \ces_5_3_io_outs_up[1] ,
    \ces_5_3_io_outs_up[0] }),
    .io_outs_down({\ces_5_3_io_ins_down[63] ,
    \ces_5_3_io_ins_down[62] ,
    \ces_5_3_io_ins_down[61] ,
    \ces_5_3_io_ins_down[60] ,
    \ces_5_3_io_ins_down[59] ,
    \ces_5_3_io_ins_down[58] ,
    \ces_5_3_io_ins_down[57] ,
    \ces_5_3_io_ins_down[56] ,
    \ces_5_3_io_ins_down[55] ,
    \ces_5_3_io_ins_down[54] ,
    \ces_5_3_io_ins_down[53] ,
    \ces_5_3_io_ins_down[52] ,
    \ces_5_3_io_ins_down[51] ,
    \ces_5_3_io_ins_down[50] ,
    \ces_5_3_io_ins_down[49] ,
    \ces_5_3_io_ins_down[48] ,
    \ces_5_3_io_ins_down[47] ,
    \ces_5_3_io_ins_down[46] ,
    \ces_5_3_io_ins_down[45] ,
    \ces_5_3_io_ins_down[44] ,
    \ces_5_3_io_ins_down[43] ,
    \ces_5_3_io_ins_down[42] ,
    \ces_5_3_io_ins_down[41] ,
    \ces_5_3_io_ins_down[40] ,
    \ces_5_3_io_ins_down[39] ,
    \ces_5_3_io_ins_down[38] ,
    \ces_5_3_io_ins_down[37] ,
    \ces_5_3_io_ins_down[36] ,
    \ces_5_3_io_ins_down[35] ,
    \ces_5_3_io_ins_down[34] ,
    \ces_5_3_io_ins_down[33] ,
    \ces_5_3_io_ins_down[32] ,
    \ces_5_3_io_ins_down[31] ,
    \ces_5_3_io_ins_down[30] ,
    \ces_5_3_io_ins_down[29] ,
    \ces_5_3_io_ins_down[28] ,
    \ces_5_3_io_ins_down[27] ,
    \ces_5_3_io_ins_down[26] ,
    \ces_5_3_io_ins_down[25] ,
    \ces_5_3_io_ins_down[24] ,
    \ces_5_3_io_ins_down[23] ,
    \ces_5_3_io_ins_down[22] ,
    \ces_5_3_io_ins_down[21] ,
    \ces_5_3_io_ins_down[20] ,
    \ces_5_3_io_ins_down[19] ,
    \ces_5_3_io_ins_down[18] ,
    \ces_5_3_io_ins_down[17] ,
    \ces_5_3_io_ins_down[16] ,
    \ces_5_3_io_ins_down[15] ,
    \ces_5_3_io_ins_down[14] ,
    \ces_5_3_io_ins_down[13] ,
    \ces_5_3_io_ins_down[12] ,
    \ces_5_3_io_ins_down[11] ,
    \ces_5_3_io_ins_down[10] ,
    \ces_5_3_io_ins_down[9] ,
    \ces_5_3_io_ins_down[8] ,
    \ces_5_3_io_ins_down[7] ,
    \ces_5_3_io_ins_down[6] ,
    \ces_5_3_io_ins_down[5] ,
    \ces_5_3_io_ins_down[4] ,
    \ces_5_3_io_ins_down[3] ,
    \ces_5_3_io_ins_down[2] ,
    \ces_5_3_io_ins_down[1] ,
    \ces_5_3_io_ins_down[0] }),
    .io_outs_left({\ces_6_2_io_ins_left[63] ,
    \ces_6_2_io_ins_left[62] ,
    \ces_6_2_io_ins_left[61] ,
    \ces_6_2_io_ins_left[60] ,
    \ces_6_2_io_ins_left[59] ,
    \ces_6_2_io_ins_left[58] ,
    \ces_6_2_io_ins_left[57] ,
    \ces_6_2_io_ins_left[56] ,
    \ces_6_2_io_ins_left[55] ,
    \ces_6_2_io_ins_left[54] ,
    \ces_6_2_io_ins_left[53] ,
    \ces_6_2_io_ins_left[52] ,
    \ces_6_2_io_ins_left[51] ,
    \ces_6_2_io_ins_left[50] ,
    \ces_6_2_io_ins_left[49] ,
    \ces_6_2_io_ins_left[48] ,
    \ces_6_2_io_ins_left[47] ,
    \ces_6_2_io_ins_left[46] ,
    \ces_6_2_io_ins_left[45] ,
    \ces_6_2_io_ins_left[44] ,
    \ces_6_2_io_ins_left[43] ,
    \ces_6_2_io_ins_left[42] ,
    \ces_6_2_io_ins_left[41] ,
    \ces_6_2_io_ins_left[40] ,
    \ces_6_2_io_ins_left[39] ,
    \ces_6_2_io_ins_left[38] ,
    \ces_6_2_io_ins_left[37] ,
    \ces_6_2_io_ins_left[36] ,
    \ces_6_2_io_ins_left[35] ,
    \ces_6_2_io_ins_left[34] ,
    \ces_6_2_io_ins_left[33] ,
    \ces_6_2_io_ins_left[32] ,
    \ces_6_2_io_ins_left[31] ,
    \ces_6_2_io_ins_left[30] ,
    \ces_6_2_io_ins_left[29] ,
    \ces_6_2_io_ins_left[28] ,
    \ces_6_2_io_ins_left[27] ,
    \ces_6_2_io_ins_left[26] ,
    \ces_6_2_io_ins_left[25] ,
    \ces_6_2_io_ins_left[24] ,
    \ces_6_2_io_ins_left[23] ,
    \ces_6_2_io_ins_left[22] ,
    \ces_6_2_io_ins_left[21] ,
    \ces_6_2_io_ins_left[20] ,
    \ces_6_2_io_ins_left[19] ,
    \ces_6_2_io_ins_left[18] ,
    \ces_6_2_io_ins_left[17] ,
    \ces_6_2_io_ins_left[16] ,
    \ces_6_2_io_ins_left[15] ,
    \ces_6_2_io_ins_left[14] ,
    \ces_6_2_io_ins_left[13] ,
    \ces_6_2_io_ins_left[12] ,
    \ces_6_2_io_ins_left[11] ,
    \ces_6_2_io_ins_left[10] ,
    \ces_6_2_io_ins_left[9] ,
    \ces_6_2_io_ins_left[8] ,
    \ces_6_2_io_ins_left[7] ,
    \ces_6_2_io_ins_left[6] ,
    \ces_6_2_io_ins_left[5] ,
    \ces_6_2_io_ins_left[4] ,
    \ces_6_2_io_ins_left[3] ,
    \ces_6_2_io_ins_left[2] ,
    \ces_6_2_io_ins_left[1] ,
    \ces_6_2_io_ins_left[0] }),
    .io_outs_right({\ces_6_3_io_outs_right[63] ,
    \ces_6_3_io_outs_right[62] ,
    \ces_6_3_io_outs_right[61] ,
    \ces_6_3_io_outs_right[60] ,
    \ces_6_3_io_outs_right[59] ,
    \ces_6_3_io_outs_right[58] ,
    \ces_6_3_io_outs_right[57] ,
    \ces_6_3_io_outs_right[56] ,
    \ces_6_3_io_outs_right[55] ,
    \ces_6_3_io_outs_right[54] ,
    \ces_6_3_io_outs_right[53] ,
    \ces_6_3_io_outs_right[52] ,
    \ces_6_3_io_outs_right[51] ,
    \ces_6_3_io_outs_right[50] ,
    \ces_6_3_io_outs_right[49] ,
    \ces_6_3_io_outs_right[48] ,
    \ces_6_3_io_outs_right[47] ,
    \ces_6_3_io_outs_right[46] ,
    \ces_6_3_io_outs_right[45] ,
    \ces_6_3_io_outs_right[44] ,
    \ces_6_3_io_outs_right[43] ,
    \ces_6_3_io_outs_right[42] ,
    \ces_6_3_io_outs_right[41] ,
    \ces_6_3_io_outs_right[40] ,
    \ces_6_3_io_outs_right[39] ,
    \ces_6_3_io_outs_right[38] ,
    \ces_6_3_io_outs_right[37] ,
    \ces_6_3_io_outs_right[36] ,
    \ces_6_3_io_outs_right[35] ,
    \ces_6_3_io_outs_right[34] ,
    \ces_6_3_io_outs_right[33] ,
    \ces_6_3_io_outs_right[32] ,
    \ces_6_3_io_outs_right[31] ,
    \ces_6_3_io_outs_right[30] ,
    \ces_6_3_io_outs_right[29] ,
    \ces_6_3_io_outs_right[28] ,
    \ces_6_3_io_outs_right[27] ,
    \ces_6_3_io_outs_right[26] ,
    \ces_6_3_io_outs_right[25] ,
    \ces_6_3_io_outs_right[24] ,
    \ces_6_3_io_outs_right[23] ,
    \ces_6_3_io_outs_right[22] ,
    \ces_6_3_io_outs_right[21] ,
    \ces_6_3_io_outs_right[20] ,
    \ces_6_3_io_outs_right[19] ,
    \ces_6_3_io_outs_right[18] ,
    \ces_6_3_io_outs_right[17] ,
    \ces_6_3_io_outs_right[16] ,
    \ces_6_3_io_outs_right[15] ,
    \ces_6_3_io_outs_right[14] ,
    \ces_6_3_io_outs_right[13] ,
    \ces_6_3_io_outs_right[12] ,
    \ces_6_3_io_outs_right[11] ,
    \ces_6_3_io_outs_right[10] ,
    \ces_6_3_io_outs_right[9] ,
    \ces_6_3_io_outs_right[8] ,
    \ces_6_3_io_outs_right[7] ,
    \ces_6_3_io_outs_right[6] ,
    \ces_6_3_io_outs_right[5] ,
    \ces_6_3_io_outs_right[4] ,
    \ces_6_3_io_outs_right[3] ,
    \ces_6_3_io_outs_right[2] ,
    \ces_6_3_io_outs_right[1] ,
    \ces_6_3_io_outs_right[0] }),
    .io_outs_up({\ces_6_3_io_outs_up[63] ,
    \ces_6_3_io_outs_up[62] ,
    \ces_6_3_io_outs_up[61] ,
    \ces_6_3_io_outs_up[60] ,
    \ces_6_3_io_outs_up[59] ,
    \ces_6_3_io_outs_up[58] ,
    \ces_6_3_io_outs_up[57] ,
    \ces_6_3_io_outs_up[56] ,
    \ces_6_3_io_outs_up[55] ,
    \ces_6_3_io_outs_up[54] ,
    \ces_6_3_io_outs_up[53] ,
    \ces_6_3_io_outs_up[52] ,
    \ces_6_3_io_outs_up[51] ,
    \ces_6_3_io_outs_up[50] ,
    \ces_6_3_io_outs_up[49] ,
    \ces_6_3_io_outs_up[48] ,
    \ces_6_3_io_outs_up[47] ,
    \ces_6_3_io_outs_up[46] ,
    \ces_6_3_io_outs_up[45] ,
    \ces_6_3_io_outs_up[44] ,
    \ces_6_3_io_outs_up[43] ,
    \ces_6_3_io_outs_up[42] ,
    \ces_6_3_io_outs_up[41] ,
    \ces_6_3_io_outs_up[40] ,
    \ces_6_3_io_outs_up[39] ,
    \ces_6_3_io_outs_up[38] ,
    \ces_6_3_io_outs_up[37] ,
    \ces_6_3_io_outs_up[36] ,
    \ces_6_3_io_outs_up[35] ,
    \ces_6_3_io_outs_up[34] ,
    \ces_6_3_io_outs_up[33] ,
    \ces_6_3_io_outs_up[32] ,
    \ces_6_3_io_outs_up[31] ,
    \ces_6_3_io_outs_up[30] ,
    \ces_6_3_io_outs_up[29] ,
    \ces_6_3_io_outs_up[28] ,
    \ces_6_3_io_outs_up[27] ,
    \ces_6_3_io_outs_up[26] ,
    \ces_6_3_io_outs_up[25] ,
    \ces_6_3_io_outs_up[24] ,
    \ces_6_3_io_outs_up[23] ,
    \ces_6_3_io_outs_up[22] ,
    \ces_6_3_io_outs_up[21] ,
    \ces_6_3_io_outs_up[20] ,
    \ces_6_3_io_outs_up[19] ,
    \ces_6_3_io_outs_up[18] ,
    \ces_6_3_io_outs_up[17] ,
    \ces_6_3_io_outs_up[16] ,
    \ces_6_3_io_outs_up[15] ,
    \ces_6_3_io_outs_up[14] ,
    \ces_6_3_io_outs_up[13] ,
    \ces_6_3_io_outs_up[12] ,
    \ces_6_3_io_outs_up[11] ,
    \ces_6_3_io_outs_up[10] ,
    \ces_6_3_io_outs_up[9] ,
    \ces_6_3_io_outs_up[8] ,
    \ces_6_3_io_outs_up[7] ,
    \ces_6_3_io_outs_up[6] ,
    \ces_6_3_io_outs_up[5] ,
    \ces_6_3_io_outs_up[4] ,
    \ces_6_3_io_outs_up[3] ,
    \ces_6_3_io_outs_up[2] ,
    \ces_6_3_io_outs_up[1] ,
    \ces_6_3_io_outs_up[0] }));
 Element ces_6_4 (.clock(clknet_3_7_0_clock),
    .io_lsbIns_1(ces_6_3_io_lsbOuts_1),
    .io_lsbIns_2(ces_6_3_io_lsbOuts_2),
    .io_lsbIns_3(ces_6_3_io_lsbOuts_3),
    .io_lsbIns_4(ces_6_3_io_lsbOuts_4),
    .io_lsbIns_5(ces_6_3_io_lsbOuts_5),
    .io_lsbIns_6(ces_6_3_io_lsbOuts_6),
    .io_lsbIns_7(ces_6_3_io_lsbOuts_7),
    .io_lsbOuts_0(ces_6_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_4_io_lsbOuts_7),
    .io_ins_down({\ces_6_4_io_ins_down[63] ,
    \ces_6_4_io_ins_down[62] ,
    \ces_6_4_io_ins_down[61] ,
    \ces_6_4_io_ins_down[60] ,
    \ces_6_4_io_ins_down[59] ,
    \ces_6_4_io_ins_down[58] ,
    \ces_6_4_io_ins_down[57] ,
    \ces_6_4_io_ins_down[56] ,
    \ces_6_4_io_ins_down[55] ,
    \ces_6_4_io_ins_down[54] ,
    \ces_6_4_io_ins_down[53] ,
    \ces_6_4_io_ins_down[52] ,
    \ces_6_4_io_ins_down[51] ,
    \ces_6_4_io_ins_down[50] ,
    \ces_6_4_io_ins_down[49] ,
    \ces_6_4_io_ins_down[48] ,
    \ces_6_4_io_ins_down[47] ,
    \ces_6_4_io_ins_down[46] ,
    \ces_6_4_io_ins_down[45] ,
    \ces_6_4_io_ins_down[44] ,
    \ces_6_4_io_ins_down[43] ,
    \ces_6_4_io_ins_down[42] ,
    \ces_6_4_io_ins_down[41] ,
    \ces_6_4_io_ins_down[40] ,
    \ces_6_4_io_ins_down[39] ,
    \ces_6_4_io_ins_down[38] ,
    \ces_6_4_io_ins_down[37] ,
    \ces_6_4_io_ins_down[36] ,
    \ces_6_4_io_ins_down[35] ,
    \ces_6_4_io_ins_down[34] ,
    \ces_6_4_io_ins_down[33] ,
    \ces_6_4_io_ins_down[32] ,
    \ces_6_4_io_ins_down[31] ,
    \ces_6_4_io_ins_down[30] ,
    \ces_6_4_io_ins_down[29] ,
    \ces_6_4_io_ins_down[28] ,
    \ces_6_4_io_ins_down[27] ,
    \ces_6_4_io_ins_down[26] ,
    \ces_6_4_io_ins_down[25] ,
    \ces_6_4_io_ins_down[24] ,
    \ces_6_4_io_ins_down[23] ,
    \ces_6_4_io_ins_down[22] ,
    \ces_6_4_io_ins_down[21] ,
    \ces_6_4_io_ins_down[20] ,
    \ces_6_4_io_ins_down[19] ,
    \ces_6_4_io_ins_down[18] ,
    \ces_6_4_io_ins_down[17] ,
    \ces_6_4_io_ins_down[16] ,
    \ces_6_4_io_ins_down[15] ,
    \ces_6_4_io_ins_down[14] ,
    \ces_6_4_io_ins_down[13] ,
    \ces_6_4_io_ins_down[12] ,
    \ces_6_4_io_ins_down[11] ,
    \ces_6_4_io_ins_down[10] ,
    \ces_6_4_io_ins_down[9] ,
    \ces_6_4_io_ins_down[8] ,
    \ces_6_4_io_ins_down[7] ,
    \ces_6_4_io_ins_down[6] ,
    \ces_6_4_io_ins_down[5] ,
    \ces_6_4_io_ins_down[4] ,
    \ces_6_4_io_ins_down[3] ,
    \ces_6_4_io_ins_down[2] ,
    \ces_6_4_io_ins_down[1] ,
    \ces_6_4_io_ins_down[0] }),
    .io_ins_left({\ces_6_4_io_ins_left[63] ,
    \ces_6_4_io_ins_left[62] ,
    \ces_6_4_io_ins_left[61] ,
    \ces_6_4_io_ins_left[60] ,
    \ces_6_4_io_ins_left[59] ,
    \ces_6_4_io_ins_left[58] ,
    \ces_6_4_io_ins_left[57] ,
    \ces_6_4_io_ins_left[56] ,
    \ces_6_4_io_ins_left[55] ,
    \ces_6_4_io_ins_left[54] ,
    \ces_6_4_io_ins_left[53] ,
    \ces_6_4_io_ins_left[52] ,
    \ces_6_4_io_ins_left[51] ,
    \ces_6_4_io_ins_left[50] ,
    \ces_6_4_io_ins_left[49] ,
    \ces_6_4_io_ins_left[48] ,
    \ces_6_4_io_ins_left[47] ,
    \ces_6_4_io_ins_left[46] ,
    \ces_6_4_io_ins_left[45] ,
    \ces_6_4_io_ins_left[44] ,
    \ces_6_4_io_ins_left[43] ,
    \ces_6_4_io_ins_left[42] ,
    \ces_6_4_io_ins_left[41] ,
    \ces_6_4_io_ins_left[40] ,
    \ces_6_4_io_ins_left[39] ,
    \ces_6_4_io_ins_left[38] ,
    \ces_6_4_io_ins_left[37] ,
    \ces_6_4_io_ins_left[36] ,
    \ces_6_4_io_ins_left[35] ,
    \ces_6_4_io_ins_left[34] ,
    \ces_6_4_io_ins_left[33] ,
    \ces_6_4_io_ins_left[32] ,
    \ces_6_4_io_ins_left[31] ,
    \ces_6_4_io_ins_left[30] ,
    \ces_6_4_io_ins_left[29] ,
    \ces_6_4_io_ins_left[28] ,
    \ces_6_4_io_ins_left[27] ,
    \ces_6_4_io_ins_left[26] ,
    \ces_6_4_io_ins_left[25] ,
    \ces_6_4_io_ins_left[24] ,
    \ces_6_4_io_ins_left[23] ,
    \ces_6_4_io_ins_left[22] ,
    \ces_6_4_io_ins_left[21] ,
    \ces_6_4_io_ins_left[20] ,
    \ces_6_4_io_ins_left[19] ,
    \ces_6_4_io_ins_left[18] ,
    \ces_6_4_io_ins_left[17] ,
    \ces_6_4_io_ins_left[16] ,
    \ces_6_4_io_ins_left[15] ,
    \ces_6_4_io_ins_left[14] ,
    \ces_6_4_io_ins_left[13] ,
    \ces_6_4_io_ins_left[12] ,
    \ces_6_4_io_ins_left[11] ,
    \ces_6_4_io_ins_left[10] ,
    \ces_6_4_io_ins_left[9] ,
    \ces_6_4_io_ins_left[8] ,
    \ces_6_4_io_ins_left[7] ,
    \ces_6_4_io_ins_left[6] ,
    \ces_6_4_io_ins_left[5] ,
    \ces_6_4_io_ins_left[4] ,
    \ces_6_4_io_ins_left[3] ,
    \ces_6_4_io_ins_left[2] ,
    \ces_6_4_io_ins_left[1] ,
    \ces_6_4_io_ins_left[0] }),
    .io_ins_right({\ces_6_3_io_outs_right[63] ,
    \ces_6_3_io_outs_right[62] ,
    \ces_6_3_io_outs_right[61] ,
    \ces_6_3_io_outs_right[60] ,
    \ces_6_3_io_outs_right[59] ,
    \ces_6_3_io_outs_right[58] ,
    \ces_6_3_io_outs_right[57] ,
    \ces_6_3_io_outs_right[56] ,
    \ces_6_3_io_outs_right[55] ,
    \ces_6_3_io_outs_right[54] ,
    \ces_6_3_io_outs_right[53] ,
    \ces_6_3_io_outs_right[52] ,
    \ces_6_3_io_outs_right[51] ,
    \ces_6_3_io_outs_right[50] ,
    \ces_6_3_io_outs_right[49] ,
    \ces_6_3_io_outs_right[48] ,
    \ces_6_3_io_outs_right[47] ,
    \ces_6_3_io_outs_right[46] ,
    \ces_6_3_io_outs_right[45] ,
    \ces_6_3_io_outs_right[44] ,
    \ces_6_3_io_outs_right[43] ,
    \ces_6_3_io_outs_right[42] ,
    \ces_6_3_io_outs_right[41] ,
    \ces_6_3_io_outs_right[40] ,
    \ces_6_3_io_outs_right[39] ,
    \ces_6_3_io_outs_right[38] ,
    \ces_6_3_io_outs_right[37] ,
    \ces_6_3_io_outs_right[36] ,
    \ces_6_3_io_outs_right[35] ,
    \ces_6_3_io_outs_right[34] ,
    \ces_6_3_io_outs_right[33] ,
    \ces_6_3_io_outs_right[32] ,
    \ces_6_3_io_outs_right[31] ,
    \ces_6_3_io_outs_right[30] ,
    \ces_6_3_io_outs_right[29] ,
    \ces_6_3_io_outs_right[28] ,
    \ces_6_3_io_outs_right[27] ,
    \ces_6_3_io_outs_right[26] ,
    \ces_6_3_io_outs_right[25] ,
    \ces_6_3_io_outs_right[24] ,
    \ces_6_3_io_outs_right[23] ,
    \ces_6_3_io_outs_right[22] ,
    \ces_6_3_io_outs_right[21] ,
    \ces_6_3_io_outs_right[20] ,
    \ces_6_3_io_outs_right[19] ,
    \ces_6_3_io_outs_right[18] ,
    \ces_6_3_io_outs_right[17] ,
    \ces_6_3_io_outs_right[16] ,
    \ces_6_3_io_outs_right[15] ,
    \ces_6_3_io_outs_right[14] ,
    \ces_6_3_io_outs_right[13] ,
    \ces_6_3_io_outs_right[12] ,
    \ces_6_3_io_outs_right[11] ,
    \ces_6_3_io_outs_right[10] ,
    \ces_6_3_io_outs_right[9] ,
    \ces_6_3_io_outs_right[8] ,
    \ces_6_3_io_outs_right[7] ,
    \ces_6_3_io_outs_right[6] ,
    \ces_6_3_io_outs_right[5] ,
    \ces_6_3_io_outs_right[4] ,
    \ces_6_3_io_outs_right[3] ,
    \ces_6_3_io_outs_right[2] ,
    \ces_6_3_io_outs_right[1] ,
    \ces_6_3_io_outs_right[0] }),
    .io_ins_up({\ces_5_4_io_outs_up[63] ,
    \ces_5_4_io_outs_up[62] ,
    \ces_5_4_io_outs_up[61] ,
    \ces_5_4_io_outs_up[60] ,
    \ces_5_4_io_outs_up[59] ,
    \ces_5_4_io_outs_up[58] ,
    \ces_5_4_io_outs_up[57] ,
    \ces_5_4_io_outs_up[56] ,
    \ces_5_4_io_outs_up[55] ,
    \ces_5_4_io_outs_up[54] ,
    \ces_5_4_io_outs_up[53] ,
    \ces_5_4_io_outs_up[52] ,
    \ces_5_4_io_outs_up[51] ,
    \ces_5_4_io_outs_up[50] ,
    \ces_5_4_io_outs_up[49] ,
    \ces_5_4_io_outs_up[48] ,
    \ces_5_4_io_outs_up[47] ,
    \ces_5_4_io_outs_up[46] ,
    \ces_5_4_io_outs_up[45] ,
    \ces_5_4_io_outs_up[44] ,
    \ces_5_4_io_outs_up[43] ,
    \ces_5_4_io_outs_up[42] ,
    \ces_5_4_io_outs_up[41] ,
    \ces_5_4_io_outs_up[40] ,
    \ces_5_4_io_outs_up[39] ,
    \ces_5_4_io_outs_up[38] ,
    \ces_5_4_io_outs_up[37] ,
    \ces_5_4_io_outs_up[36] ,
    \ces_5_4_io_outs_up[35] ,
    \ces_5_4_io_outs_up[34] ,
    \ces_5_4_io_outs_up[33] ,
    \ces_5_4_io_outs_up[32] ,
    \ces_5_4_io_outs_up[31] ,
    \ces_5_4_io_outs_up[30] ,
    \ces_5_4_io_outs_up[29] ,
    \ces_5_4_io_outs_up[28] ,
    \ces_5_4_io_outs_up[27] ,
    \ces_5_4_io_outs_up[26] ,
    \ces_5_4_io_outs_up[25] ,
    \ces_5_4_io_outs_up[24] ,
    \ces_5_4_io_outs_up[23] ,
    \ces_5_4_io_outs_up[22] ,
    \ces_5_4_io_outs_up[21] ,
    \ces_5_4_io_outs_up[20] ,
    \ces_5_4_io_outs_up[19] ,
    \ces_5_4_io_outs_up[18] ,
    \ces_5_4_io_outs_up[17] ,
    \ces_5_4_io_outs_up[16] ,
    \ces_5_4_io_outs_up[15] ,
    \ces_5_4_io_outs_up[14] ,
    \ces_5_4_io_outs_up[13] ,
    \ces_5_4_io_outs_up[12] ,
    \ces_5_4_io_outs_up[11] ,
    \ces_5_4_io_outs_up[10] ,
    \ces_5_4_io_outs_up[9] ,
    \ces_5_4_io_outs_up[8] ,
    \ces_5_4_io_outs_up[7] ,
    \ces_5_4_io_outs_up[6] ,
    \ces_5_4_io_outs_up[5] ,
    \ces_5_4_io_outs_up[4] ,
    \ces_5_4_io_outs_up[3] ,
    \ces_5_4_io_outs_up[2] ,
    \ces_5_4_io_outs_up[1] ,
    \ces_5_4_io_outs_up[0] }),
    .io_outs_down({\ces_5_4_io_ins_down[63] ,
    \ces_5_4_io_ins_down[62] ,
    \ces_5_4_io_ins_down[61] ,
    \ces_5_4_io_ins_down[60] ,
    \ces_5_4_io_ins_down[59] ,
    \ces_5_4_io_ins_down[58] ,
    \ces_5_4_io_ins_down[57] ,
    \ces_5_4_io_ins_down[56] ,
    \ces_5_4_io_ins_down[55] ,
    \ces_5_4_io_ins_down[54] ,
    \ces_5_4_io_ins_down[53] ,
    \ces_5_4_io_ins_down[52] ,
    \ces_5_4_io_ins_down[51] ,
    \ces_5_4_io_ins_down[50] ,
    \ces_5_4_io_ins_down[49] ,
    \ces_5_4_io_ins_down[48] ,
    \ces_5_4_io_ins_down[47] ,
    \ces_5_4_io_ins_down[46] ,
    \ces_5_4_io_ins_down[45] ,
    \ces_5_4_io_ins_down[44] ,
    \ces_5_4_io_ins_down[43] ,
    \ces_5_4_io_ins_down[42] ,
    \ces_5_4_io_ins_down[41] ,
    \ces_5_4_io_ins_down[40] ,
    \ces_5_4_io_ins_down[39] ,
    \ces_5_4_io_ins_down[38] ,
    \ces_5_4_io_ins_down[37] ,
    \ces_5_4_io_ins_down[36] ,
    \ces_5_4_io_ins_down[35] ,
    \ces_5_4_io_ins_down[34] ,
    \ces_5_4_io_ins_down[33] ,
    \ces_5_4_io_ins_down[32] ,
    \ces_5_4_io_ins_down[31] ,
    \ces_5_4_io_ins_down[30] ,
    \ces_5_4_io_ins_down[29] ,
    \ces_5_4_io_ins_down[28] ,
    \ces_5_4_io_ins_down[27] ,
    \ces_5_4_io_ins_down[26] ,
    \ces_5_4_io_ins_down[25] ,
    \ces_5_4_io_ins_down[24] ,
    \ces_5_4_io_ins_down[23] ,
    \ces_5_4_io_ins_down[22] ,
    \ces_5_4_io_ins_down[21] ,
    \ces_5_4_io_ins_down[20] ,
    \ces_5_4_io_ins_down[19] ,
    \ces_5_4_io_ins_down[18] ,
    \ces_5_4_io_ins_down[17] ,
    \ces_5_4_io_ins_down[16] ,
    \ces_5_4_io_ins_down[15] ,
    \ces_5_4_io_ins_down[14] ,
    \ces_5_4_io_ins_down[13] ,
    \ces_5_4_io_ins_down[12] ,
    \ces_5_4_io_ins_down[11] ,
    \ces_5_4_io_ins_down[10] ,
    \ces_5_4_io_ins_down[9] ,
    \ces_5_4_io_ins_down[8] ,
    \ces_5_4_io_ins_down[7] ,
    \ces_5_4_io_ins_down[6] ,
    \ces_5_4_io_ins_down[5] ,
    \ces_5_4_io_ins_down[4] ,
    \ces_5_4_io_ins_down[3] ,
    \ces_5_4_io_ins_down[2] ,
    \ces_5_4_io_ins_down[1] ,
    \ces_5_4_io_ins_down[0] }),
    .io_outs_left({\ces_6_3_io_ins_left[63] ,
    \ces_6_3_io_ins_left[62] ,
    \ces_6_3_io_ins_left[61] ,
    \ces_6_3_io_ins_left[60] ,
    \ces_6_3_io_ins_left[59] ,
    \ces_6_3_io_ins_left[58] ,
    \ces_6_3_io_ins_left[57] ,
    \ces_6_3_io_ins_left[56] ,
    \ces_6_3_io_ins_left[55] ,
    \ces_6_3_io_ins_left[54] ,
    \ces_6_3_io_ins_left[53] ,
    \ces_6_3_io_ins_left[52] ,
    \ces_6_3_io_ins_left[51] ,
    \ces_6_3_io_ins_left[50] ,
    \ces_6_3_io_ins_left[49] ,
    \ces_6_3_io_ins_left[48] ,
    \ces_6_3_io_ins_left[47] ,
    \ces_6_3_io_ins_left[46] ,
    \ces_6_3_io_ins_left[45] ,
    \ces_6_3_io_ins_left[44] ,
    \ces_6_3_io_ins_left[43] ,
    \ces_6_3_io_ins_left[42] ,
    \ces_6_3_io_ins_left[41] ,
    \ces_6_3_io_ins_left[40] ,
    \ces_6_3_io_ins_left[39] ,
    \ces_6_3_io_ins_left[38] ,
    \ces_6_3_io_ins_left[37] ,
    \ces_6_3_io_ins_left[36] ,
    \ces_6_3_io_ins_left[35] ,
    \ces_6_3_io_ins_left[34] ,
    \ces_6_3_io_ins_left[33] ,
    \ces_6_3_io_ins_left[32] ,
    \ces_6_3_io_ins_left[31] ,
    \ces_6_3_io_ins_left[30] ,
    \ces_6_3_io_ins_left[29] ,
    \ces_6_3_io_ins_left[28] ,
    \ces_6_3_io_ins_left[27] ,
    \ces_6_3_io_ins_left[26] ,
    \ces_6_3_io_ins_left[25] ,
    \ces_6_3_io_ins_left[24] ,
    \ces_6_3_io_ins_left[23] ,
    \ces_6_3_io_ins_left[22] ,
    \ces_6_3_io_ins_left[21] ,
    \ces_6_3_io_ins_left[20] ,
    \ces_6_3_io_ins_left[19] ,
    \ces_6_3_io_ins_left[18] ,
    \ces_6_3_io_ins_left[17] ,
    \ces_6_3_io_ins_left[16] ,
    \ces_6_3_io_ins_left[15] ,
    \ces_6_3_io_ins_left[14] ,
    \ces_6_3_io_ins_left[13] ,
    \ces_6_3_io_ins_left[12] ,
    \ces_6_3_io_ins_left[11] ,
    \ces_6_3_io_ins_left[10] ,
    \ces_6_3_io_ins_left[9] ,
    \ces_6_3_io_ins_left[8] ,
    \ces_6_3_io_ins_left[7] ,
    \ces_6_3_io_ins_left[6] ,
    \ces_6_3_io_ins_left[5] ,
    \ces_6_3_io_ins_left[4] ,
    \ces_6_3_io_ins_left[3] ,
    \ces_6_3_io_ins_left[2] ,
    \ces_6_3_io_ins_left[1] ,
    \ces_6_3_io_ins_left[0] }),
    .io_outs_right({\ces_6_4_io_outs_right[63] ,
    \ces_6_4_io_outs_right[62] ,
    \ces_6_4_io_outs_right[61] ,
    \ces_6_4_io_outs_right[60] ,
    \ces_6_4_io_outs_right[59] ,
    \ces_6_4_io_outs_right[58] ,
    \ces_6_4_io_outs_right[57] ,
    \ces_6_4_io_outs_right[56] ,
    \ces_6_4_io_outs_right[55] ,
    \ces_6_4_io_outs_right[54] ,
    \ces_6_4_io_outs_right[53] ,
    \ces_6_4_io_outs_right[52] ,
    \ces_6_4_io_outs_right[51] ,
    \ces_6_4_io_outs_right[50] ,
    \ces_6_4_io_outs_right[49] ,
    \ces_6_4_io_outs_right[48] ,
    \ces_6_4_io_outs_right[47] ,
    \ces_6_4_io_outs_right[46] ,
    \ces_6_4_io_outs_right[45] ,
    \ces_6_4_io_outs_right[44] ,
    \ces_6_4_io_outs_right[43] ,
    \ces_6_4_io_outs_right[42] ,
    \ces_6_4_io_outs_right[41] ,
    \ces_6_4_io_outs_right[40] ,
    \ces_6_4_io_outs_right[39] ,
    \ces_6_4_io_outs_right[38] ,
    \ces_6_4_io_outs_right[37] ,
    \ces_6_4_io_outs_right[36] ,
    \ces_6_4_io_outs_right[35] ,
    \ces_6_4_io_outs_right[34] ,
    \ces_6_4_io_outs_right[33] ,
    \ces_6_4_io_outs_right[32] ,
    \ces_6_4_io_outs_right[31] ,
    \ces_6_4_io_outs_right[30] ,
    \ces_6_4_io_outs_right[29] ,
    \ces_6_4_io_outs_right[28] ,
    \ces_6_4_io_outs_right[27] ,
    \ces_6_4_io_outs_right[26] ,
    \ces_6_4_io_outs_right[25] ,
    \ces_6_4_io_outs_right[24] ,
    \ces_6_4_io_outs_right[23] ,
    \ces_6_4_io_outs_right[22] ,
    \ces_6_4_io_outs_right[21] ,
    \ces_6_4_io_outs_right[20] ,
    \ces_6_4_io_outs_right[19] ,
    \ces_6_4_io_outs_right[18] ,
    \ces_6_4_io_outs_right[17] ,
    \ces_6_4_io_outs_right[16] ,
    \ces_6_4_io_outs_right[15] ,
    \ces_6_4_io_outs_right[14] ,
    \ces_6_4_io_outs_right[13] ,
    \ces_6_4_io_outs_right[12] ,
    \ces_6_4_io_outs_right[11] ,
    \ces_6_4_io_outs_right[10] ,
    \ces_6_4_io_outs_right[9] ,
    \ces_6_4_io_outs_right[8] ,
    \ces_6_4_io_outs_right[7] ,
    \ces_6_4_io_outs_right[6] ,
    \ces_6_4_io_outs_right[5] ,
    \ces_6_4_io_outs_right[4] ,
    \ces_6_4_io_outs_right[3] ,
    \ces_6_4_io_outs_right[2] ,
    \ces_6_4_io_outs_right[1] ,
    \ces_6_4_io_outs_right[0] }),
    .io_outs_up({\ces_6_4_io_outs_up[63] ,
    \ces_6_4_io_outs_up[62] ,
    \ces_6_4_io_outs_up[61] ,
    \ces_6_4_io_outs_up[60] ,
    \ces_6_4_io_outs_up[59] ,
    \ces_6_4_io_outs_up[58] ,
    \ces_6_4_io_outs_up[57] ,
    \ces_6_4_io_outs_up[56] ,
    \ces_6_4_io_outs_up[55] ,
    \ces_6_4_io_outs_up[54] ,
    \ces_6_4_io_outs_up[53] ,
    \ces_6_4_io_outs_up[52] ,
    \ces_6_4_io_outs_up[51] ,
    \ces_6_4_io_outs_up[50] ,
    \ces_6_4_io_outs_up[49] ,
    \ces_6_4_io_outs_up[48] ,
    \ces_6_4_io_outs_up[47] ,
    \ces_6_4_io_outs_up[46] ,
    \ces_6_4_io_outs_up[45] ,
    \ces_6_4_io_outs_up[44] ,
    \ces_6_4_io_outs_up[43] ,
    \ces_6_4_io_outs_up[42] ,
    \ces_6_4_io_outs_up[41] ,
    \ces_6_4_io_outs_up[40] ,
    \ces_6_4_io_outs_up[39] ,
    \ces_6_4_io_outs_up[38] ,
    \ces_6_4_io_outs_up[37] ,
    \ces_6_4_io_outs_up[36] ,
    \ces_6_4_io_outs_up[35] ,
    \ces_6_4_io_outs_up[34] ,
    \ces_6_4_io_outs_up[33] ,
    \ces_6_4_io_outs_up[32] ,
    \ces_6_4_io_outs_up[31] ,
    \ces_6_4_io_outs_up[30] ,
    \ces_6_4_io_outs_up[29] ,
    \ces_6_4_io_outs_up[28] ,
    \ces_6_4_io_outs_up[27] ,
    \ces_6_4_io_outs_up[26] ,
    \ces_6_4_io_outs_up[25] ,
    \ces_6_4_io_outs_up[24] ,
    \ces_6_4_io_outs_up[23] ,
    \ces_6_4_io_outs_up[22] ,
    \ces_6_4_io_outs_up[21] ,
    \ces_6_4_io_outs_up[20] ,
    \ces_6_4_io_outs_up[19] ,
    \ces_6_4_io_outs_up[18] ,
    \ces_6_4_io_outs_up[17] ,
    \ces_6_4_io_outs_up[16] ,
    \ces_6_4_io_outs_up[15] ,
    \ces_6_4_io_outs_up[14] ,
    \ces_6_4_io_outs_up[13] ,
    \ces_6_4_io_outs_up[12] ,
    \ces_6_4_io_outs_up[11] ,
    \ces_6_4_io_outs_up[10] ,
    \ces_6_4_io_outs_up[9] ,
    \ces_6_4_io_outs_up[8] ,
    \ces_6_4_io_outs_up[7] ,
    \ces_6_4_io_outs_up[6] ,
    \ces_6_4_io_outs_up[5] ,
    \ces_6_4_io_outs_up[4] ,
    \ces_6_4_io_outs_up[3] ,
    \ces_6_4_io_outs_up[2] ,
    \ces_6_4_io_outs_up[1] ,
    \ces_6_4_io_outs_up[0] }));
 Element ces_6_5 (.clock(clknet_3_7_0_clock),
    .io_lsbIns_1(ces_6_4_io_lsbOuts_1),
    .io_lsbIns_2(ces_6_4_io_lsbOuts_2),
    .io_lsbIns_3(ces_6_4_io_lsbOuts_3),
    .io_lsbIns_4(ces_6_4_io_lsbOuts_4),
    .io_lsbIns_5(ces_6_4_io_lsbOuts_5),
    .io_lsbIns_6(ces_6_4_io_lsbOuts_6),
    .io_lsbIns_7(ces_6_4_io_lsbOuts_7),
    .io_lsbOuts_0(ces_6_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_5_io_lsbOuts_7),
    .io_ins_down({\ces_6_5_io_ins_down[63] ,
    \ces_6_5_io_ins_down[62] ,
    \ces_6_5_io_ins_down[61] ,
    \ces_6_5_io_ins_down[60] ,
    \ces_6_5_io_ins_down[59] ,
    \ces_6_5_io_ins_down[58] ,
    \ces_6_5_io_ins_down[57] ,
    \ces_6_5_io_ins_down[56] ,
    \ces_6_5_io_ins_down[55] ,
    \ces_6_5_io_ins_down[54] ,
    \ces_6_5_io_ins_down[53] ,
    \ces_6_5_io_ins_down[52] ,
    \ces_6_5_io_ins_down[51] ,
    \ces_6_5_io_ins_down[50] ,
    \ces_6_5_io_ins_down[49] ,
    \ces_6_5_io_ins_down[48] ,
    \ces_6_5_io_ins_down[47] ,
    \ces_6_5_io_ins_down[46] ,
    \ces_6_5_io_ins_down[45] ,
    \ces_6_5_io_ins_down[44] ,
    \ces_6_5_io_ins_down[43] ,
    \ces_6_5_io_ins_down[42] ,
    \ces_6_5_io_ins_down[41] ,
    \ces_6_5_io_ins_down[40] ,
    \ces_6_5_io_ins_down[39] ,
    \ces_6_5_io_ins_down[38] ,
    \ces_6_5_io_ins_down[37] ,
    \ces_6_5_io_ins_down[36] ,
    \ces_6_5_io_ins_down[35] ,
    \ces_6_5_io_ins_down[34] ,
    \ces_6_5_io_ins_down[33] ,
    \ces_6_5_io_ins_down[32] ,
    \ces_6_5_io_ins_down[31] ,
    \ces_6_5_io_ins_down[30] ,
    \ces_6_5_io_ins_down[29] ,
    \ces_6_5_io_ins_down[28] ,
    \ces_6_5_io_ins_down[27] ,
    \ces_6_5_io_ins_down[26] ,
    \ces_6_5_io_ins_down[25] ,
    \ces_6_5_io_ins_down[24] ,
    \ces_6_5_io_ins_down[23] ,
    \ces_6_5_io_ins_down[22] ,
    \ces_6_5_io_ins_down[21] ,
    \ces_6_5_io_ins_down[20] ,
    \ces_6_5_io_ins_down[19] ,
    \ces_6_5_io_ins_down[18] ,
    \ces_6_5_io_ins_down[17] ,
    \ces_6_5_io_ins_down[16] ,
    \ces_6_5_io_ins_down[15] ,
    \ces_6_5_io_ins_down[14] ,
    \ces_6_5_io_ins_down[13] ,
    \ces_6_5_io_ins_down[12] ,
    \ces_6_5_io_ins_down[11] ,
    \ces_6_5_io_ins_down[10] ,
    \ces_6_5_io_ins_down[9] ,
    \ces_6_5_io_ins_down[8] ,
    \ces_6_5_io_ins_down[7] ,
    \ces_6_5_io_ins_down[6] ,
    \ces_6_5_io_ins_down[5] ,
    \ces_6_5_io_ins_down[4] ,
    \ces_6_5_io_ins_down[3] ,
    \ces_6_5_io_ins_down[2] ,
    \ces_6_5_io_ins_down[1] ,
    \ces_6_5_io_ins_down[0] }),
    .io_ins_left({\ces_6_5_io_ins_left[63] ,
    \ces_6_5_io_ins_left[62] ,
    \ces_6_5_io_ins_left[61] ,
    \ces_6_5_io_ins_left[60] ,
    \ces_6_5_io_ins_left[59] ,
    \ces_6_5_io_ins_left[58] ,
    \ces_6_5_io_ins_left[57] ,
    \ces_6_5_io_ins_left[56] ,
    \ces_6_5_io_ins_left[55] ,
    \ces_6_5_io_ins_left[54] ,
    \ces_6_5_io_ins_left[53] ,
    \ces_6_5_io_ins_left[52] ,
    \ces_6_5_io_ins_left[51] ,
    \ces_6_5_io_ins_left[50] ,
    \ces_6_5_io_ins_left[49] ,
    \ces_6_5_io_ins_left[48] ,
    \ces_6_5_io_ins_left[47] ,
    \ces_6_5_io_ins_left[46] ,
    \ces_6_5_io_ins_left[45] ,
    \ces_6_5_io_ins_left[44] ,
    \ces_6_5_io_ins_left[43] ,
    \ces_6_5_io_ins_left[42] ,
    \ces_6_5_io_ins_left[41] ,
    \ces_6_5_io_ins_left[40] ,
    \ces_6_5_io_ins_left[39] ,
    \ces_6_5_io_ins_left[38] ,
    \ces_6_5_io_ins_left[37] ,
    \ces_6_5_io_ins_left[36] ,
    \ces_6_5_io_ins_left[35] ,
    \ces_6_5_io_ins_left[34] ,
    \ces_6_5_io_ins_left[33] ,
    \ces_6_5_io_ins_left[32] ,
    \ces_6_5_io_ins_left[31] ,
    \ces_6_5_io_ins_left[30] ,
    \ces_6_5_io_ins_left[29] ,
    \ces_6_5_io_ins_left[28] ,
    \ces_6_5_io_ins_left[27] ,
    \ces_6_5_io_ins_left[26] ,
    \ces_6_5_io_ins_left[25] ,
    \ces_6_5_io_ins_left[24] ,
    \ces_6_5_io_ins_left[23] ,
    \ces_6_5_io_ins_left[22] ,
    \ces_6_5_io_ins_left[21] ,
    \ces_6_5_io_ins_left[20] ,
    \ces_6_5_io_ins_left[19] ,
    \ces_6_5_io_ins_left[18] ,
    \ces_6_5_io_ins_left[17] ,
    \ces_6_5_io_ins_left[16] ,
    \ces_6_5_io_ins_left[15] ,
    \ces_6_5_io_ins_left[14] ,
    \ces_6_5_io_ins_left[13] ,
    \ces_6_5_io_ins_left[12] ,
    \ces_6_5_io_ins_left[11] ,
    \ces_6_5_io_ins_left[10] ,
    \ces_6_5_io_ins_left[9] ,
    \ces_6_5_io_ins_left[8] ,
    \ces_6_5_io_ins_left[7] ,
    \ces_6_5_io_ins_left[6] ,
    \ces_6_5_io_ins_left[5] ,
    \ces_6_5_io_ins_left[4] ,
    \ces_6_5_io_ins_left[3] ,
    \ces_6_5_io_ins_left[2] ,
    \ces_6_5_io_ins_left[1] ,
    \ces_6_5_io_ins_left[0] }),
    .io_ins_right({\ces_6_4_io_outs_right[63] ,
    \ces_6_4_io_outs_right[62] ,
    \ces_6_4_io_outs_right[61] ,
    \ces_6_4_io_outs_right[60] ,
    \ces_6_4_io_outs_right[59] ,
    \ces_6_4_io_outs_right[58] ,
    \ces_6_4_io_outs_right[57] ,
    \ces_6_4_io_outs_right[56] ,
    \ces_6_4_io_outs_right[55] ,
    \ces_6_4_io_outs_right[54] ,
    \ces_6_4_io_outs_right[53] ,
    \ces_6_4_io_outs_right[52] ,
    \ces_6_4_io_outs_right[51] ,
    \ces_6_4_io_outs_right[50] ,
    \ces_6_4_io_outs_right[49] ,
    \ces_6_4_io_outs_right[48] ,
    \ces_6_4_io_outs_right[47] ,
    \ces_6_4_io_outs_right[46] ,
    \ces_6_4_io_outs_right[45] ,
    \ces_6_4_io_outs_right[44] ,
    \ces_6_4_io_outs_right[43] ,
    \ces_6_4_io_outs_right[42] ,
    \ces_6_4_io_outs_right[41] ,
    \ces_6_4_io_outs_right[40] ,
    \ces_6_4_io_outs_right[39] ,
    \ces_6_4_io_outs_right[38] ,
    \ces_6_4_io_outs_right[37] ,
    \ces_6_4_io_outs_right[36] ,
    \ces_6_4_io_outs_right[35] ,
    \ces_6_4_io_outs_right[34] ,
    \ces_6_4_io_outs_right[33] ,
    \ces_6_4_io_outs_right[32] ,
    \ces_6_4_io_outs_right[31] ,
    \ces_6_4_io_outs_right[30] ,
    \ces_6_4_io_outs_right[29] ,
    \ces_6_4_io_outs_right[28] ,
    \ces_6_4_io_outs_right[27] ,
    \ces_6_4_io_outs_right[26] ,
    \ces_6_4_io_outs_right[25] ,
    \ces_6_4_io_outs_right[24] ,
    \ces_6_4_io_outs_right[23] ,
    \ces_6_4_io_outs_right[22] ,
    \ces_6_4_io_outs_right[21] ,
    \ces_6_4_io_outs_right[20] ,
    \ces_6_4_io_outs_right[19] ,
    \ces_6_4_io_outs_right[18] ,
    \ces_6_4_io_outs_right[17] ,
    \ces_6_4_io_outs_right[16] ,
    \ces_6_4_io_outs_right[15] ,
    \ces_6_4_io_outs_right[14] ,
    \ces_6_4_io_outs_right[13] ,
    \ces_6_4_io_outs_right[12] ,
    \ces_6_4_io_outs_right[11] ,
    \ces_6_4_io_outs_right[10] ,
    \ces_6_4_io_outs_right[9] ,
    \ces_6_4_io_outs_right[8] ,
    \ces_6_4_io_outs_right[7] ,
    \ces_6_4_io_outs_right[6] ,
    \ces_6_4_io_outs_right[5] ,
    \ces_6_4_io_outs_right[4] ,
    \ces_6_4_io_outs_right[3] ,
    \ces_6_4_io_outs_right[2] ,
    \ces_6_4_io_outs_right[1] ,
    \ces_6_4_io_outs_right[0] }),
    .io_ins_up({\ces_5_5_io_outs_up[63] ,
    \ces_5_5_io_outs_up[62] ,
    \ces_5_5_io_outs_up[61] ,
    \ces_5_5_io_outs_up[60] ,
    \ces_5_5_io_outs_up[59] ,
    \ces_5_5_io_outs_up[58] ,
    \ces_5_5_io_outs_up[57] ,
    \ces_5_5_io_outs_up[56] ,
    \ces_5_5_io_outs_up[55] ,
    \ces_5_5_io_outs_up[54] ,
    \ces_5_5_io_outs_up[53] ,
    \ces_5_5_io_outs_up[52] ,
    \ces_5_5_io_outs_up[51] ,
    \ces_5_5_io_outs_up[50] ,
    \ces_5_5_io_outs_up[49] ,
    \ces_5_5_io_outs_up[48] ,
    \ces_5_5_io_outs_up[47] ,
    \ces_5_5_io_outs_up[46] ,
    \ces_5_5_io_outs_up[45] ,
    \ces_5_5_io_outs_up[44] ,
    \ces_5_5_io_outs_up[43] ,
    \ces_5_5_io_outs_up[42] ,
    \ces_5_5_io_outs_up[41] ,
    \ces_5_5_io_outs_up[40] ,
    \ces_5_5_io_outs_up[39] ,
    \ces_5_5_io_outs_up[38] ,
    \ces_5_5_io_outs_up[37] ,
    \ces_5_5_io_outs_up[36] ,
    \ces_5_5_io_outs_up[35] ,
    \ces_5_5_io_outs_up[34] ,
    \ces_5_5_io_outs_up[33] ,
    \ces_5_5_io_outs_up[32] ,
    \ces_5_5_io_outs_up[31] ,
    \ces_5_5_io_outs_up[30] ,
    \ces_5_5_io_outs_up[29] ,
    \ces_5_5_io_outs_up[28] ,
    \ces_5_5_io_outs_up[27] ,
    \ces_5_5_io_outs_up[26] ,
    \ces_5_5_io_outs_up[25] ,
    \ces_5_5_io_outs_up[24] ,
    \ces_5_5_io_outs_up[23] ,
    \ces_5_5_io_outs_up[22] ,
    \ces_5_5_io_outs_up[21] ,
    \ces_5_5_io_outs_up[20] ,
    \ces_5_5_io_outs_up[19] ,
    \ces_5_5_io_outs_up[18] ,
    \ces_5_5_io_outs_up[17] ,
    \ces_5_5_io_outs_up[16] ,
    \ces_5_5_io_outs_up[15] ,
    \ces_5_5_io_outs_up[14] ,
    \ces_5_5_io_outs_up[13] ,
    \ces_5_5_io_outs_up[12] ,
    \ces_5_5_io_outs_up[11] ,
    \ces_5_5_io_outs_up[10] ,
    \ces_5_5_io_outs_up[9] ,
    \ces_5_5_io_outs_up[8] ,
    \ces_5_5_io_outs_up[7] ,
    \ces_5_5_io_outs_up[6] ,
    \ces_5_5_io_outs_up[5] ,
    \ces_5_5_io_outs_up[4] ,
    \ces_5_5_io_outs_up[3] ,
    \ces_5_5_io_outs_up[2] ,
    \ces_5_5_io_outs_up[1] ,
    \ces_5_5_io_outs_up[0] }),
    .io_outs_down({\ces_5_5_io_ins_down[63] ,
    \ces_5_5_io_ins_down[62] ,
    \ces_5_5_io_ins_down[61] ,
    \ces_5_5_io_ins_down[60] ,
    \ces_5_5_io_ins_down[59] ,
    \ces_5_5_io_ins_down[58] ,
    \ces_5_5_io_ins_down[57] ,
    \ces_5_5_io_ins_down[56] ,
    \ces_5_5_io_ins_down[55] ,
    \ces_5_5_io_ins_down[54] ,
    \ces_5_5_io_ins_down[53] ,
    \ces_5_5_io_ins_down[52] ,
    \ces_5_5_io_ins_down[51] ,
    \ces_5_5_io_ins_down[50] ,
    \ces_5_5_io_ins_down[49] ,
    \ces_5_5_io_ins_down[48] ,
    \ces_5_5_io_ins_down[47] ,
    \ces_5_5_io_ins_down[46] ,
    \ces_5_5_io_ins_down[45] ,
    \ces_5_5_io_ins_down[44] ,
    \ces_5_5_io_ins_down[43] ,
    \ces_5_5_io_ins_down[42] ,
    \ces_5_5_io_ins_down[41] ,
    \ces_5_5_io_ins_down[40] ,
    \ces_5_5_io_ins_down[39] ,
    \ces_5_5_io_ins_down[38] ,
    \ces_5_5_io_ins_down[37] ,
    \ces_5_5_io_ins_down[36] ,
    \ces_5_5_io_ins_down[35] ,
    \ces_5_5_io_ins_down[34] ,
    \ces_5_5_io_ins_down[33] ,
    \ces_5_5_io_ins_down[32] ,
    \ces_5_5_io_ins_down[31] ,
    \ces_5_5_io_ins_down[30] ,
    \ces_5_5_io_ins_down[29] ,
    \ces_5_5_io_ins_down[28] ,
    \ces_5_5_io_ins_down[27] ,
    \ces_5_5_io_ins_down[26] ,
    \ces_5_5_io_ins_down[25] ,
    \ces_5_5_io_ins_down[24] ,
    \ces_5_5_io_ins_down[23] ,
    \ces_5_5_io_ins_down[22] ,
    \ces_5_5_io_ins_down[21] ,
    \ces_5_5_io_ins_down[20] ,
    \ces_5_5_io_ins_down[19] ,
    \ces_5_5_io_ins_down[18] ,
    \ces_5_5_io_ins_down[17] ,
    \ces_5_5_io_ins_down[16] ,
    \ces_5_5_io_ins_down[15] ,
    \ces_5_5_io_ins_down[14] ,
    \ces_5_5_io_ins_down[13] ,
    \ces_5_5_io_ins_down[12] ,
    \ces_5_5_io_ins_down[11] ,
    \ces_5_5_io_ins_down[10] ,
    \ces_5_5_io_ins_down[9] ,
    \ces_5_5_io_ins_down[8] ,
    \ces_5_5_io_ins_down[7] ,
    \ces_5_5_io_ins_down[6] ,
    \ces_5_5_io_ins_down[5] ,
    \ces_5_5_io_ins_down[4] ,
    \ces_5_5_io_ins_down[3] ,
    \ces_5_5_io_ins_down[2] ,
    \ces_5_5_io_ins_down[1] ,
    \ces_5_5_io_ins_down[0] }),
    .io_outs_left({\ces_6_4_io_ins_left[63] ,
    \ces_6_4_io_ins_left[62] ,
    \ces_6_4_io_ins_left[61] ,
    \ces_6_4_io_ins_left[60] ,
    \ces_6_4_io_ins_left[59] ,
    \ces_6_4_io_ins_left[58] ,
    \ces_6_4_io_ins_left[57] ,
    \ces_6_4_io_ins_left[56] ,
    \ces_6_4_io_ins_left[55] ,
    \ces_6_4_io_ins_left[54] ,
    \ces_6_4_io_ins_left[53] ,
    \ces_6_4_io_ins_left[52] ,
    \ces_6_4_io_ins_left[51] ,
    \ces_6_4_io_ins_left[50] ,
    \ces_6_4_io_ins_left[49] ,
    \ces_6_4_io_ins_left[48] ,
    \ces_6_4_io_ins_left[47] ,
    \ces_6_4_io_ins_left[46] ,
    \ces_6_4_io_ins_left[45] ,
    \ces_6_4_io_ins_left[44] ,
    \ces_6_4_io_ins_left[43] ,
    \ces_6_4_io_ins_left[42] ,
    \ces_6_4_io_ins_left[41] ,
    \ces_6_4_io_ins_left[40] ,
    \ces_6_4_io_ins_left[39] ,
    \ces_6_4_io_ins_left[38] ,
    \ces_6_4_io_ins_left[37] ,
    \ces_6_4_io_ins_left[36] ,
    \ces_6_4_io_ins_left[35] ,
    \ces_6_4_io_ins_left[34] ,
    \ces_6_4_io_ins_left[33] ,
    \ces_6_4_io_ins_left[32] ,
    \ces_6_4_io_ins_left[31] ,
    \ces_6_4_io_ins_left[30] ,
    \ces_6_4_io_ins_left[29] ,
    \ces_6_4_io_ins_left[28] ,
    \ces_6_4_io_ins_left[27] ,
    \ces_6_4_io_ins_left[26] ,
    \ces_6_4_io_ins_left[25] ,
    \ces_6_4_io_ins_left[24] ,
    \ces_6_4_io_ins_left[23] ,
    \ces_6_4_io_ins_left[22] ,
    \ces_6_4_io_ins_left[21] ,
    \ces_6_4_io_ins_left[20] ,
    \ces_6_4_io_ins_left[19] ,
    \ces_6_4_io_ins_left[18] ,
    \ces_6_4_io_ins_left[17] ,
    \ces_6_4_io_ins_left[16] ,
    \ces_6_4_io_ins_left[15] ,
    \ces_6_4_io_ins_left[14] ,
    \ces_6_4_io_ins_left[13] ,
    \ces_6_4_io_ins_left[12] ,
    \ces_6_4_io_ins_left[11] ,
    \ces_6_4_io_ins_left[10] ,
    \ces_6_4_io_ins_left[9] ,
    \ces_6_4_io_ins_left[8] ,
    \ces_6_4_io_ins_left[7] ,
    \ces_6_4_io_ins_left[6] ,
    \ces_6_4_io_ins_left[5] ,
    \ces_6_4_io_ins_left[4] ,
    \ces_6_4_io_ins_left[3] ,
    \ces_6_4_io_ins_left[2] ,
    \ces_6_4_io_ins_left[1] ,
    \ces_6_4_io_ins_left[0] }),
    .io_outs_right({\ces_6_5_io_outs_right[63] ,
    \ces_6_5_io_outs_right[62] ,
    \ces_6_5_io_outs_right[61] ,
    \ces_6_5_io_outs_right[60] ,
    \ces_6_5_io_outs_right[59] ,
    \ces_6_5_io_outs_right[58] ,
    \ces_6_5_io_outs_right[57] ,
    \ces_6_5_io_outs_right[56] ,
    \ces_6_5_io_outs_right[55] ,
    \ces_6_5_io_outs_right[54] ,
    \ces_6_5_io_outs_right[53] ,
    \ces_6_5_io_outs_right[52] ,
    \ces_6_5_io_outs_right[51] ,
    \ces_6_5_io_outs_right[50] ,
    \ces_6_5_io_outs_right[49] ,
    \ces_6_5_io_outs_right[48] ,
    \ces_6_5_io_outs_right[47] ,
    \ces_6_5_io_outs_right[46] ,
    \ces_6_5_io_outs_right[45] ,
    \ces_6_5_io_outs_right[44] ,
    \ces_6_5_io_outs_right[43] ,
    \ces_6_5_io_outs_right[42] ,
    \ces_6_5_io_outs_right[41] ,
    \ces_6_5_io_outs_right[40] ,
    \ces_6_5_io_outs_right[39] ,
    \ces_6_5_io_outs_right[38] ,
    \ces_6_5_io_outs_right[37] ,
    \ces_6_5_io_outs_right[36] ,
    \ces_6_5_io_outs_right[35] ,
    \ces_6_5_io_outs_right[34] ,
    \ces_6_5_io_outs_right[33] ,
    \ces_6_5_io_outs_right[32] ,
    \ces_6_5_io_outs_right[31] ,
    \ces_6_5_io_outs_right[30] ,
    \ces_6_5_io_outs_right[29] ,
    \ces_6_5_io_outs_right[28] ,
    \ces_6_5_io_outs_right[27] ,
    \ces_6_5_io_outs_right[26] ,
    \ces_6_5_io_outs_right[25] ,
    \ces_6_5_io_outs_right[24] ,
    \ces_6_5_io_outs_right[23] ,
    \ces_6_5_io_outs_right[22] ,
    \ces_6_5_io_outs_right[21] ,
    \ces_6_5_io_outs_right[20] ,
    \ces_6_5_io_outs_right[19] ,
    \ces_6_5_io_outs_right[18] ,
    \ces_6_5_io_outs_right[17] ,
    \ces_6_5_io_outs_right[16] ,
    \ces_6_5_io_outs_right[15] ,
    \ces_6_5_io_outs_right[14] ,
    \ces_6_5_io_outs_right[13] ,
    \ces_6_5_io_outs_right[12] ,
    \ces_6_5_io_outs_right[11] ,
    \ces_6_5_io_outs_right[10] ,
    \ces_6_5_io_outs_right[9] ,
    \ces_6_5_io_outs_right[8] ,
    \ces_6_5_io_outs_right[7] ,
    \ces_6_5_io_outs_right[6] ,
    \ces_6_5_io_outs_right[5] ,
    \ces_6_5_io_outs_right[4] ,
    \ces_6_5_io_outs_right[3] ,
    \ces_6_5_io_outs_right[2] ,
    \ces_6_5_io_outs_right[1] ,
    \ces_6_5_io_outs_right[0] }),
    .io_outs_up({\ces_6_5_io_outs_up[63] ,
    \ces_6_5_io_outs_up[62] ,
    \ces_6_5_io_outs_up[61] ,
    \ces_6_5_io_outs_up[60] ,
    \ces_6_5_io_outs_up[59] ,
    \ces_6_5_io_outs_up[58] ,
    \ces_6_5_io_outs_up[57] ,
    \ces_6_5_io_outs_up[56] ,
    \ces_6_5_io_outs_up[55] ,
    \ces_6_5_io_outs_up[54] ,
    \ces_6_5_io_outs_up[53] ,
    \ces_6_5_io_outs_up[52] ,
    \ces_6_5_io_outs_up[51] ,
    \ces_6_5_io_outs_up[50] ,
    \ces_6_5_io_outs_up[49] ,
    \ces_6_5_io_outs_up[48] ,
    \ces_6_5_io_outs_up[47] ,
    \ces_6_5_io_outs_up[46] ,
    \ces_6_5_io_outs_up[45] ,
    \ces_6_5_io_outs_up[44] ,
    \ces_6_5_io_outs_up[43] ,
    \ces_6_5_io_outs_up[42] ,
    \ces_6_5_io_outs_up[41] ,
    \ces_6_5_io_outs_up[40] ,
    \ces_6_5_io_outs_up[39] ,
    \ces_6_5_io_outs_up[38] ,
    \ces_6_5_io_outs_up[37] ,
    \ces_6_5_io_outs_up[36] ,
    \ces_6_5_io_outs_up[35] ,
    \ces_6_5_io_outs_up[34] ,
    \ces_6_5_io_outs_up[33] ,
    \ces_6_5_io_outs_up[32] ,
    \ces_6_5_io_outs_up[31] ,
    \ces_6_5_io_outs_up[30] ,
    \ces_6_5_io_outs_up[29] ,
    \ces_6_5_io_outs_up[28] ,
    \ces_6_5_io_outs_up[27] ,
    \ces_6_5_io_outs_up[26] ,
    \ces_6_5_io_outs_up[25] ,
    \ces_6_5_io_outs_up[24] ,
    \ces_6_5_io_outs_up[23] ,
    \ces_6_5_io_outs_up[22] ,
    \ces_6_5_io_outs_up[21] ,
    \ces_6_5_io_outs_up[20] ,
    \ces_6_5_io_outs_up[19] ,
    \ces_6_5_io_outs_up[18] ,
    \ces_6_5_io_outs_up[17] ,
    \ces_6_5_io_outs_up[16] ,
    \ces_6_5_io_outs_up[15] ,
    \ces_6_5_io_outs_up[14] ,
    \ces_6_5_io_outs_up[13] ,
    \ces_6_5_io_outs_up[12] ,
    \ces_6_5_io_outs_up[11] ,
    \ces_6_5_io_outs_up[10] ,
    \ces_6_5_io_outs_up[9] ,
    \ces_6_5_io_outs_up[8] ,
    \ces_6_5_io_outs_up[7] ,
    \ces_6_5_io_outs_up[6] ,
    \ces_6_5_io_outs_up[5] ,
    \ces_6_5_io_outs_up[4] ,
    \ces_6_5_io_outs_up[3] ,
    \ces_6_5_io_outs_up[2] ,
    \ces_6_5_io_outs_up[1] ,
    \ces_6_5_io_outs_up[0] }));
 Element ces_6_6 (.clock(clknet_3_7_0_clock),
    .io_lsbIns_1(ces_6_5_io_lsbOuts_1),
    .io_lsbIns_2(ces_6_5_io_lsbOuts_2),
    .io_lsbIns_3(ces_6_5_io_lsbOuts_3),
    .io_lsbIns_4(ces_6_5_io_lsbOuts_4),
    .io_lsbIns_5(ces_6_5_io_lsbOuts_5),
    .io_lsbIns_6(ces_6_5_io_lsbOuts_6),
    .io_lsbIns_7(ces_6_5_io_lsbOuts_7),
    .io_lsbOuts_0(ces_6_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_6_io_lsbOuts_7),
    .io_ins_down({\ces_6_6_io_ins_down[63] ,
    \ces_6_6_io_ins_down[62] ,
    \ces_6_6_io_ins_down[61] ,
    \ces_6_6_io_ins_down[60] ,
    \ces_6_6_io_ins_down[59] ,
    \ces_6_6_io_ins_down[58] ,
    \ces_6_6_io_ins_down[57] ,
    \ces_6_6_io_ins_down[56] ,
    \ces_6_6_io_ins_down[55] ,
    \ces_6_6_io_ins_down[54] ,
    \ces_6_6_io_ins_down[53] ,
    \ces_6_6_io_ins_down[52] ,
    \ces_6_6_io_ins_down[51] ,
    \ces_6_6_io_ins_down[50] ,
    \ces_6_6_io_ins_down[49] ,
    \ces_6_6_io_ins_down[48] ,
    \ces_6_6_io_ins_down[47] ,
    \ces_6_6_io_ins_down[46] ,
    \ces_6_6_io_ins_down[45] ,
    \ces_6_6_io_ins_down[44] ,
    \ces_6_6_io_ins_down[43] ,
    \ces_6_6_io_ins_down[42] ,
    \ces_6_6_io_ins_down[41] ,
    \ces_6_6_io_ins_down[40] ,
    \ces_6_6_io_ins_down[39] ,
    \ces_6_6_io_ins_down[38] ,
    \ces_6_6_io_ins_down[37] ,
    \ces_6_6_io_ins_down[36] ,
    \ces_6_6_io_ins_down[35] ,
    \ces_6_6_io_ins_down[34] ,
    \ces_6_6_io_ins_down[33] ,
    \ces_6_6_io_ins_down[32] ,
    \ces_6_6_io_ins_down[31] ,
    \ces_6_6_io_ins_down[30] ,
    \ces_6_6_io_ins_down[29] ,
    \ces_6_6_io_ins_down[28] ,
    \ces_6_6_io_ins_down[27] ,
    \ces_6_6_io_ins_down[26] ,
    \ces_6_6_io_ins_down[25] ,
    \ces_6_6_io_ins_down[24] ,
    \ces_6_6_io_ins_down[23] ,
    \ces_6_6_io_ins_down[22] ,
    \ces_6_6_io_ins_down[21] ,
    \ces_6_6_io_ins_down[20] ,
    \ces_6_6_io_ins_down[19] ,
    \ces_6_6_io_ins_down[18] ,
    \ces_6_6_io_ins_down[17] ,
    \ces_6_6_io_ins_down[16] ,
    \ces_6_6_io_ins_down[15] ,
    \ces_6_6_io_ins_down[14] ,
    \ces_6_6_io_ins_down[13] ,
    \ces_6_6_io_ins_down[12] ,
    \ces_6_6_io_ins_down[11] ,
    \ces_6_6_io_ins_down[10] ,
    \ces_6_6_io_ins_down[9] ,
    \ces_6_6_io_ins_down[8] ,
    \ces_6_6_io_ins_down[7] ,
    \ces_6_6_io_ins_down[6] ,
    \ces_6_6_io_ins_down[5] ,
    \ces_6_6_io_ins_down[4] ,
    \ces_6_6_io_ins_down[3] ,
    \ces_6_6_io_ins_down[2] ,
    \ces_6_6_io_ins_down[1] ,
    \ces_6_6_io_ins_down[0] }),
    .io_ins_left({\ces_6_6_io_ins_left[63] ,
    \ces_6_6_io_ins_left[62] ,
    \ces_6_6_io_ins_left[61] ,
    \ces_6_6_io_ins_left[60] ,
    \ces_6_6_io_ins_left[59] ,
    \ces_6_6_io_ins_left[58] ,
    \ces_6_6_io_ins_left[57] ,
    \ces_6_6_io_ins_left[56] ,
    \ces_6_6_io_ins_left[55] ,
    \ces_6_6_io_ins_left[54] ,
    \ces_6_6_io_ins_left[53] ,
    \ces_6_6_io_ins_left[52] ,
    \ces_6_6_io_ins_left[51] ,
    \ces_6_6_io_ins_left[50] ,
    \ces_6_6_io_ins_left[49] ,
    \ces_6_6_io_ins_left[48] ,
    \ces_6_6_io_ins_left[47] ,
    \ces_6_6_io_ins_left[46] ,
    \ces_6_6_io_ins_left[45] ,
    \ces_6_6_io_ins_left[44] ,
    \ces_6_6_io_ins_left[43] ,
    \ces_6_6_io_ins_left[42] ,
    \ces_6_6_io_ins_left[41] ,
    \ces_6_6_io_ins_left[40] ,
    \ces_6_6_io_ins_left[39] ,
    \ces_6_6_io_ins_left[38] ,
    \ces_6_6_io_ins_left[37] ,
    \ces_6_6_io_ins_left[36] ,
    \ces_6_6_io_ins_left[35] ,
    \ces_6_6_io_ins_left[34] ,
    \ces_6_6_io_ins_left[33] ,
    \ces_6_6_io_ins_left[32] ,
    \ces_6_6_io_ins_left[31] ,
    \ces_6_6_io_ins_left[30] ,
    \ces_6_6_io_ins_left[29] ,
    \ces_6_6_io_ins_left[28] ,
    \ces_6_6_io_ins_left[27] ,
    \ces_6_6_io_ins_left[26] ,
    \ces_6_6_io_ins_left[25] ,
    \ces_6_6_io_ins_left[24] ,
    \ces_6_6_io_ins_left[23] ,
    \ces_6_6_io_ins_left[22] ,
    \ces_6_6_io_ins_left[21] ,
    \ces_6_6_io_ins_left[20] ,
    \ces_6_6_io_ins_left[19] ,
    \ces_6_6_io_ins_left[18] ,
    \ces_6_6_io_ins_left[17] ,
    \ces_6_6_io_ins_left[16] ,
    \ces_6_6_io_ins_left[15] ,
    \ces_6_6_io_ins_left[14] ,
    \ces_6_6_io_ins_left[13] ,
    \ces_6_6_io_ins_left[12] ,
    \ces_6_6_io_ins_left[11] ,
    \ces_6_6_io_ins_left[10] ,
    \ces_6_6_io_ins_left[9] ,
    \ces_6_6_io_ins_left[8] ,
    \ces_6_6_io_ins_left[7] ,
    \ces_6_6_io_ins_left[6] ,
    \ces_6_6_io_ins_left[5] ,
    \ces_6_6_io_ins_left[4] ,
    \ces_6_6_io_ins_left[3] ,
    \ces_6_6_io_ins_left[2] ,
    \ces_6_6_io_ins_left[1] ,
    \ces_6_6_io_ins_left[0] }),
    .io_ins_right({\ces_6_5_io_outs_right[63] ,
    \ces_6_5_io_outs_right[62] ,
    \ces_6_5_io_outs_right[61] ,
    \ces_6_5_io_outs_right[60] ,
    \ces_6_5_io_outs_right[59] ,
    \ces_6_5_io_outs_right[58] ,
    \ces_6_5_io_outs_right[57] ,
    \ces_6_5_io_outs_right[56] ,
    \ces_6_5_io_outs_right[55] ,
    \ces_6_5_io_outs_right[54] ,
    \ces_6_5_io_outs_right[53] ,
    \ces_6_5_io_outs_right[52] ,
    \ces_6_5_io_outs_right[51] ,
    \ces_6_5_io_outs_right[50] ,
    \ces_6_5_io_outs_right[49] ,
    \ces_6_5_io_outs_right[48] ,
    \ces_6_5_io_outs_right[47] ,
    \ces_6_5_io_outs_right[46] ,
    \ces_6_5_io_outs_right[45] ,
    \ces_6_5_io_outs_right[44] ,
    \ces_6_5_io_outs_right[43] ,
    \ces_6_5_io_outs_right[42] ,
    \ces_6_5_io_outs_right[41] ,
    \ces_6_5_io_outs_right[40] ,
    \ces_6_5_io_outs_right[39] ,
    \ces_6_5_io_outs_right[38] ,
    \ces_6_5_io_outs_right[37] ,
    \ces_6_5_io_outs_right[36] ,
    \ces_6_5_io_outs_right[35] ,
    \ces_6_5_io_outs_right[34] ,
    \ces_6_5_io_outs_right[33] ,
    \ces_6_5_io_outs_right[32] ,
    \ces_6_5_io_outs_right[31] ,
    \ces_6_5_io_outs_right[30] ,
    \ces_6_5_io_outs_right[29] ,
    \ces_6_5_io_outs_right[28] ,
    \ces_6_5_io_outs_right[27] ,
    \ces_6_5_io_outs_right[26] ,
    \ces_6_5_io_outs_right[25] ,
    \ces_6_5_io_outs_right[24] ,
    \ces_6_5_io_outs_right[23] ,
    \ces_6_5_io_outs_right[22] ,
    \ces_6_5_io_outs_right[21] ,
    \ces_6_5_io_outs_right[20] ,
    \ces_6_5_io_outs_right[19] ,
    \ces_6_5_io_outs_right[18] ,
    \ces_6_5_io_outs_right[17] ,
    \ces_6_5_io_outs_right[16] ,
    \ces_6_5_io_outs_right[15] ,
    \ces_6_5_io_outs_right[14] ,
    \ces_6_5_io_outs_right[13] ,
    \ces_6_5_io_outs_right[12] ,
    \ces_6_5_io_outs_right[11] ,
    \ces_6_5_io_outs_right[10] ,
    \ces_6_5_io_outs_right[9] ,
    \ces_6_5_io_outs_right[8] ,
    \ces_6_5_io_outs_right[7] ,
    \ces_6_5_io_outs_right[6] ,
    \ces_6_5_io_outs_right[5] ,
    \ces_6_5_io_outs_right[4] ,
    \ces_6_5_io_outs_right[3] ,
    \ces_6_5_io_outs_right[2] ,
    \ces_6_5_io_outs_right[1] ,
    \ces_6_5_io_outs_right[0] }),
    .io_ins_up({\ces_5_6_io_outs_up[63] ,
    \ces_5_6_io_outs_up[62] ,
    \ces_5_6_io_outs_up[61] ,
    \ces_5_6_io_outs_up[60] ,
    \ces_5_6_io_outs_up[59] ,
    \ces_5_6_io_outs_up[58] ,
    \ces_5_6_io_outs_up[57] ,
    \ces_5_6_io_outs_up[56] ,
    \ces_5_6_io_outs_up[55] ,
    \ces_5_6_io_outs_up[54] ,
    \ces_5_6_io_outs_up[53] ,
    \ces_5_6_io_outs_up[52] ,
    \ces_5_6_io_outs_up[51] ,
    \ces_5_6_io_outs_up[50] ,
    \ces_5_6_io_outs_up[49] ,
    \ces_5_6_io_outs_up[48] ,
    \ces_5_6_io_outs_up[47] ,
    \ces_5_6_io_outs_up[46] ,
    \ces_5_6_io_outs_up[45] ,
    \ces_5_6_io_outs_up[44] ,
    \ces_5_6_io_outs_up[43] ,
    \ces_5_6_io_outs_up[42] ,
    \ces_5_6_io_outs_up[41] ,
    \ces_5_6_io_outs_up[40] ,
    \ces_5_6_io_outs_up[39] ,
    \ces_5_6_io_outs_up[38] ,
    \ces_5_6_io_outs_up[37] ,
    \ces_5_6_io_outs_up[36] ,
    \ces_5_6_io_outs_up[35] ,
    \ces_5_6_io_outs_up[34] ,
    \ces_5_6_io_outs_up[33] ,
    \ces_5_6_io_outs_up[32] ,
    \ces_5_6_io_outs_up[31] ,
    \ces_5_6_io_outs_up[30] ,
    \ces_5_6_io_outs_up[29] ,
    \ces_5_6_io_outs_up[28] ,
    \ces_5_6_io_outs_up[27] ,
    \ces_5_6_io_outs_up[26] ,
    \ces_5_6_io_outs_up[25] ,
    \ces_5_6_io_outs_up[24] ,
    \ces_5_6_io_outs_up[23] ,
    \ces_5_6_io_outs_up[22] ,
    \ces_5_6_io_outs_up[21] ,
    \ces_5_6_io_outs_up[20] ,
    \ces_5_6_io_outs_up[19] ,
    \ces_5_6_io_outs_up[18] ,
    \ces_5_6_io_outs_up[17] ,
    \ces_5_6_io_outs_up[16] ,
    \ces_5_6_io_outs_up[15] ,
    \ces_5_6_io_outs_up[14] ,
    \ces_5_6_io_outs_up[13] ,
    \ces_5_6_io_outs_up[12] ,
    \ces_5_6_io_outs_up[11] ,
    \ces_5_6_io_outs_up[10] ,
    \ces_5_6_io_outs_up[9] ,
    \ces_5_6_io_outs_up[8] ,
    \ces_5_6_io_outs_up[7] ,
    \ces_5_6_io_outs_up[6] ,
    \ces_5_6_io_outs_up[5] ,
    \ces_5_6_io_outs_up[4] ,
    \ces_5_6_io_outs_up[3] ,
    \ces_5_6_io_outs_up[2] ,
    \ces_5_6_io_outs_up[1] ,
    \ces_5_6_io_outs_up[0] }),
    .io_outs_down({\ces_5_6_io_ins_down[63] ,
    \ces_5_6_io_ins_down[62] ,
    \ces_5_6_io_ins_down[61] ,
    \ces_5_6_io_ins_down[60] ,
    \ces_5_6_io_ins_down[59] ,
    \ces_5_6_io_ins_down[58] ,
    \ces_5_6_io_ins_down[57] ,
    \ces_5_6_io_ins_down[56] ,
    \ces_5_6_io_ins_down[55] ,
    \ces_5_6_io_ins_down[54] ,
    \ces_5_6_io_ins_down[53] ,
    \ces_5_6_io_ins_down[52] ,
    \ces_5_6_io_ins_down[51] ,
    \ces_5_6_io_ins_down[50] ,
    \ces_5_6_io_ins_down[49] ,
    \ces_5_6_io_ins_down[48] ,
    \ces_5_6_io_ins_down[47] ,
    \ces_5_6_io_ins_down[46] ,
    \ces_5_6_io_ins_down[45] ,
    \ces_5_6_io_ins_down[44] ,
    \ces_5_6_io_ins_down[43] ,
    \ces_5_6_io_ins_down[42] ,
    \ces_5_6_io_ins_down[41] ,
    \ces_5_6_io_ins_down[40] ,
    \ces_5_6_io_ins_down[39] ,
    \ces_5_6_io_ins_down[38] ,
    \ces_5_6_io_ins_down[37] ,
    \ces_5_6_io_ins_down[36] ,
    \ces_5_6_io_ins_down[35] ,
    \ces_5_6_io_ins_down[34] ,
    \ces_5_6_io_ins_down[33] ,
    \ces_5_6_io_ins_down[32] ,
    \ces_5_6_io_ins_down[31] ,
    \ces_5_6_io_ins_down[30] ,
    \ces_5_6_io_ins_down[29] ,
    \ces_5_6_io_ins_down[28] ,
    \ces_5_6_io_ins_down[27] ,
    \ces_5_6_io_ins_down[26] ,
    \ces_5_6_io_ins_down[25] ,
    \ces_5_6_io_ins_down[24] ,
    \ces_5_6_io_ins_down[23] ,
    \ces_5_6_io_ins_down[22] ,
    \ces_5_6_io_ins_down[21] ,
    \ces_5_6_io_ins_down[20] ,
    \ces_5_6_io_ins_down[19] ,
    \ces_5_6_io_ins_down[18] ,
    \ces_5_6_io_ins_down[17] ,
    \ces_5_6_io_ins_down[16] ,
    \ces_5_6_io_ins_down[15] ,
    \ces_5_6_io_ins_down[14] ,
    \ces_5_6_io_ins_down[13] ,
    \ces_5_6_io_ins_down[12] ,
    \ces_5_6_io_ins_down[11] ,
    \ces_5_6_io_ins_down[10] ,
    \ces_5_6_io_ins_down[9] ,
    \ces_5_6_io_ins_down[8] ,
    \ces_5_6_io_ins_down[7] ,
    \ces_5_6_io_ins_down[6] ,
    \ces_5_6_io_ins_down[5] ,
    \ces_5_6_io_ins_down[4] ,
    \ces_5_6_io_ins_down[3] ,
    \ces_5_6_io_ins_down[2] ,
    \ces_5_6_io_ins_down[1] ,
    \ces_5_6_io_ins_down[0] }),
    .io_outs_left({\ces_6_5_io_ins_left[63] ,
    \ces_6_5_io_ins_left[62] ,
    \ces_6_5_io_ins_left[61] ,
    \ces_6_5_io_ins_left[60] ,
    \ces_6_5_io_ins_left[59] ,
    \ces_6_5_io_ins_left[58] ,
    \ces_6_5_io_ins_left[57] ,
    \ces_6_5_io_ins_left[56] ,
    \ces_6_5_io_ins_left[55] ,
    \ces_6_5_io_ins_left[54] ,
    \ces_6_5_io_ins_left[53] ,
    \ces_6_5_io_ins_left[52] ,
    \ces_6_5_io_ins_left[51] ,
    \ces_6_5_io_ins_left[50] ,
    \ces_6_5_io_ins_left[49] ,
    \ces_6_5_io_ins_left[48] ,
    \ces_6_5_io_ins_left[47] ,
    \ces_6_5_io_ins_left[46] ,
    \ces_6_5_io_ins_left[45] ,
    \ces_6_5_io_ins_left[44] ,
    \ces_6_5_io_ins_left[43] ,
    \ces_6_5_io_ins_left[42] ,
    \ces_6_5_io_ins_left[41] ,
    \ces_6_5_io_ins_left[40] ,
    \ces_6_5_io_ins_left[39] ,
    \ces_6_5_io_ins_left[38] ,
    \ces_6_5_io_ins_left[37] ,
    \ces_6_5_io_ins_left[36] ,
    \ces_6_5_io_ins_left[35] ,
    \ces_6_5_io_ins_left[34] ,
    \ces_6_5_io_ins_left[33] ,
    \ces_6_5_io_ins_left[32] ,
    \ces_6_5_io_ins_left[31] ,
    \ces_6_5_io_ins_left[30] ,
    \ces_6_5_io_ins_left[29] ,
    \ces_6_5_io_ins_left[28] ,
    \ces_6_5_io_ins_left[27] ,
    \ces_6_5_io_ins_left[26] ,
    \ces_6_5_io_ins_left[25] ,
    \ces_6_5_io_ins_left[24] ,
    \ces_6_5_io_ins_left[23] ,
    \ces_6_5_io_ins_left[22] ,
    \ces_6_5_io_ins_left[21] ,
    \ces_6_5_io_ins_left[20] ,
    \ces_6_5_io_ins_left[19] ,
    \ces_6_5_io_ins_left[18] ,
    \ces_6_5_io_ins_left[17] ,
    \ces_6_5_io_ins_left[16] ,
    \ces_6_5_io_ins_left[15] ,
    \ces_6_5_io_ins_left[14] ,
    \ces_6_5_io_ins_left[13] ,
    \ces_6_5_io_ins_left[12] ,
    \ces_6_5_io_ins_left[11] ,
    \ces_6_5_io_ins_left[10] ,
    \ces_6_5_io_ins_left[9] ,
    \ces_6_5_io_ins_left[8] ,
    \ces_6_5_io_ins_left[7] ,
    \ces_6_5_io_ins_left[6] ,
    \ces_6_5_io_ins_left[5] ,
    \ces_6_5_io_ins_left[4] ,
    \ces_6_5_io_ins_left[3] ,
    \ces_6_5_io_ins_left[2] ,
    \ces_6_5_io_ins_left[1] ,
    \ces_6_5_io_ins_left[0] }),
    .io_outs_right({\ces_6_6_io_outs_right[63] ,
    \ces_6_6_io_outs_right[62] ,
    \ces_6_6_io_outs_right[61] ,
    \ces_6_6_io_outs_right[60] ,
    \ces_6_6_io_outs_right[59] ,
    \ces_6_6_io_outs_right[58] ,
    \ces_6_6_io_outs_right[57] ,
    \ces_6_6_io_outs_right[56] ,
    \ces_6_6_io_outs_right[55] ,
    \ces_6_6_io_outs_right[54] ,
    \ces_6_6_io_outs_right[53] ,
    \ces_6_6_io_outs_right[52] ,
    \ces_6_6_io_outs_right[51] ,
    \ces_6_6_io_outs_right[50] ,
    \ces_6_6_io_outs_right[49] ,
    \ces_6_6_io_outs_right[48] ,
    \ces_6_6_io_outs_right[47] ,
    \ces_6_6_io_outs_right[46] ,
    \ces_6_6_io_outs_right[45] ,
    \ces_6_6_io_outs_right[44] ,
    \ces_6_6_io_outs_right[43] ,
    \ces_6_6_io_outs_right[42] ,
    \ces_6_6_io_outs_right[41] ,
    \ces_6_6_io_outs_right[40] ,
    \ces_6_6_io_outs_right[39] ,
    \ces_6_6_io_outs_right[38] ,
    \ces_6_6_io_outs_right[37] ,
    \ces_6_6_io_outs_right[36] ,
    \ces_6_6_io_outs_right[35] ,
    \ces_6_6_io_outs_right[34] ,
    \ces_6_6_io_outs_right[33] ,
    \ces_6_6_io_outs_right[32] ,
    \ces_6_6_io_outs_right[31] ,
    \ces_6_6_io_outs_right[30] ,
    \ces_6_6_io_outs_right[29] ,
    \ces_6_6_io_outs_right[28] ,
    \ces_6_6_io_outs_right[27] ,
    \ces_6_6_io_outs_right[26] ,
    \ces_6_6_io_outs_right[25] ,
    \ces_6_6_io_outs_right[24] ,
    \ces_6_6_io_outs_right[23] ,
    \ces_6_6_io_outs_right[22] ,
    \ces_6_6_io_outs_right[21] ,
    \ces_6_6_io_outs_right[20] ,
    \ces_6_6_io_outs_right[19] ,
    \ces_6_6_io_outs_right[18] ,
    \ces_6_6_io_outs_right[17] ,
    \ces_6_6_io_outs_right[16] ,
    \ces_6_6_io_outs_right[15] ,
    \ces_6_6_io_outs_right[14] ,
    \ces_6_6_io_outs_right[13] ,
    \ces_6_6_io_outs_right[12] ,
    \ces_6_6_io_outs_right[11] ,
    \ces_6_6_io_outs_right[10] ,
    \ces_6_6_io_outs_right[9] ,
    \ces_6_6_io_outs_right[8] ,
    \ces_6_6_io_outs_right[7] ,
    \ces_6_6_io_outs_right[6] ,
    \ces_6_6_io_outs_right[5] ,
    \ces_6_6_io_outs_right[4] ,
    \ces_6_6_io_outs_right[3] ,
    \ces_6_6_io_outs_right[2] ,
    \ces_6_6_io_outs_right[1] ,
    \ces_6_6_io_outs_right[0] }),
    .io_outs_up({\ces_6_6_io_outs_up[63] ,
    \ces_6_6_io_outs_up[62] ,
    \ces_6_6_io_outs_up[61] ,
    \ces_6_6_io_outs_up[60] ,
    \ces_6_6_io_outs_up[59] ,
    \ces_6_6_io_outs_up[58] ,
    \ces_6_6_io_outs_up[57] ,
    \ces_6_6_io_outs_up[56] ,
    \ces_6_6_io_outs_up[55] ,
    \ces_6_6_io_outs_up[54] ,
    \ces_6_6_io_outs_up[53] ,
    \ces_6_6_io_outs_up[52] ,
    \ces_6_6_io_outs_up[51] ,
    \ces_6_6_io_outs_up[50] ,
    \ces_6_6_io_outs_up[49] ,
    \ces_6_6_io_outs_up[48] ,
    \ces_6_6_io_outs_up[47] ,
    \ces_6_6_io_outs_up[46] ,
    \ces_6_6_io_outs_up[45] ,
    \ces_6_6_io_outs_up[44] ,
    \ces_6_6_io_outs_up[43] ,
    \ces_6_6_io_outs_up[42] ,
    \ces_6_6_io_outs_up[41] ,
    \ces_6_6_io_outs_up[40] ,
    \ces_6_6_io_outs_up[39] ,
    \ces_6_6_io_outs_up[38] ,
    \ces_6_6_io_outs_up[37] ,
    \ces_6_6_io_outs_up[36] ,
    \ces_6_6_io_outs_up[35] ,
    \ces_6_6_io_outs_up[34] ,
    \ces_6_6_io_outs_up[33] ,
    \ces_6_6_io_outs_up[32] ,
    \ces_6_6_io_outs_up[31] ,
    \ces_6_6_io_outs_up[30] ,
    \ces_6_6_io_outs_up[29] ,
    \ces_6_6_io_outs_up[28] ,
    \ces_6_6_io_outs_up[27] ,
    \ces_6_6_io_outs_up[26] ,
    \ces_6_6_io_outs_up[25] ,
    \ces_6_6_io_outs_up[24] ,
    \ces_6_6_io_outs_up[23] ,
    \ces_6_6_io_outs_up[22] ,
    \ces_6_6_io_outs_up[21] ,
    \ces_6_6_io_outs_up[20] ,
    \ces_6_6_io_outs_up[19] ,
    \ces_6_6_io_outs_up[18] ,
    \ces_6_6_io_outs_up[17] ,
    \ces_6_6_io_outs_up[16] ,
    \ces_6_6_io_outs_up[15] ,
    \ces_6_6_io_outs_up[14] ,
    \ces_6_6_io_outs_up[13] ,
    \ces_6_6_io_outs_up[12] ,
    \ces_6_6_io_outs_up[11] ,
    \ces_6_6_io_outs_up[10] ,
    \ces_6_6_io_outs_up[9] ,
    \ces_6_6_io_outs_up[8] ,
    \ces_6_6_io_outs_up[7] ,
    \ces_6_6_io_outs_up[6] ,
    \ces_6_6_io_outs_up[5] ,
    \ces_6_6_io_outs_up[4] ,
    \ces_6_6_io_outs_up[3] ,
    \ces_6_6_io_outs_up[2] ,
    \ces_6_6_io_outs_up[1] ,
    \ces_6_6_io_outs_up[0] }));
 Element ces_6_7 (.clock(clknet_3_7_0_clock),
    .io_lsbIns_1(ces_6_6_io_lsbOuts_1),
    .io_lsbIns_2(ces_6_6_io_lsbOuts_2),
    .io_lsbIns_3(ces_6_6_io_lsbOuts_3),
    .io_lsbIns_4(ces_6_6_io_lsbOuts_4),
    .io_lsbIns_5(ces_6_6_io_lsbOuts_5),
    .io_lsbIns_6(ces_6_6_io_lsbOuts_6),
    .io_lsbIns_7(ces_6_6_io_lsbOuts_7),
    .io_lsbOuts_0(ces_6_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_6_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_6_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_6_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_6_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_6_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_6_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_6_7_io_lsbOuts_7),
    .io_ins_down({\ces_6_7_io_ins_down[63] ,
    \ces_6_7_io_ins_down[62] ,
    \ces_6_7_io_ins_down[61] ,
    \ces_6_7_io_ins_down[60] ,
    \ces_6_7_io_ins_down[59] ,
    \ces_6_7_io_ins_down[58] ,
    \ces_6_7_io_ins_down[57] ,
    \ces_6_7_io_ins_down[56] ,
    \ces_6_7_io_ins_down[55] ,
    \ces_6_7_io_ins_down[54] ,
    \ces_6_7_io_ins_down[53] ,
    \ces_6_7_io_ins_down[52] ,
    \ces_6_7_io_ins_down[51] ,
    \ces_6_7_io_ins_down[50] ,
    \ces_6_7_io_ins_down[49] ,
    \ces_6_7_io_ins_down[48] ,
    \ces_6_7_io_ins_down[47] ,
    \ces_6_7_io_ins_down[46] ,
    \ces_6_7_io_ins_down[45] ,
    \ces_6_7_io_ins_down[44] ,
    \ces_6_7_io_ins_down[43] ,
    \ces_6_7_io_ins_down[42] ,
    \ces_6_7_io_ins_down[41] ,
    \ces_6_7_io_ins_down[40] ,
    \ces_6_7_io_ins_down[39] ,
    \ces_6_7_io_ins_down[38] ,
    \ces_6_7_io_ins_down[37] ,
    \ces_6_7_io_ins_down[36] ,
    \ces_6_7_io_ins_down[35] ,
    \ces_6_7_io_ins_down[34] ,
    \ces_6_7_io_ins_down[33] ,
    \ces_6_7_io_ins_down[32] ,
    \ces_6_7_io_ins_down[31] ,
    \ces_6_7_io_ins_down[30] ,
    \ces_6_7_io_ins_down[29] ,
    \ces_6_7_io_ins_down[28] ,
    \ces_6_7_io_ins_down[27] ,
    \ces_6_7_io_ins_down[26] ,
    \ces_6_7_io_ins_down[25] ,
    \ces_6_7_io_ins_down[24] ,
    \ces_6_7_io_ins_down[23] ,
    \ces_6_7_io_ins_down[22] ,
    \ces_6_7_io_ins_down[21] ,
    \ces_6_7_io_ins_down[20] ,
    \ces_6_7_io_ins_down[19] ,
    \ces_6_7_io_ins_down[18] ,
    \ces_6_7_io_ins_down[17] ,
    \ces_6_7_io_ins_down[16] ,
    \ces_6_7_io_ins_down[15] ,
    \ces_6_7_io_ins_down[14] ,
    \ces_6_7_io_ins_down[13] ,
    \ces_6_7_io_ins_down[12] ,
    \ces_6_7_io_ins_down[11] ,
    \ces_6_7_io_ins_down[10] ,
    \ces_6_7_io_ins_down[9] ,
    \ces_6_7_io_ins_down[8] ,
    \ces_6_7_io_ins_down[7] ,
    \ces_6_7_io_ins_down[6] ,
    \ces_6_7_io_ins_down[5] ,
    \ces_6_7_io_ins_down[4] ,
    \ces_6_7_io_ins_down[3] ,
    \ces_6_7_io_ins_down[2] ,
    \ces_6_7_io_ins_down[1] ,
    \ces_6_7_io_ins_down[0] }),
    .io_ins_left({net956,
    net955,
    net954,
    net953,
    net951,
    net950,
    net949,
    net948,
    net947,
    net946,
    net945,
    net944,
    net943,
    net942,
    net940,
    net939,
    net938,
    net937,
    net936,
    net935,
    net934,
    net933,
    net932,
    net931,
    net929,
    net928,
    net927,
    net926,
    net925,
    net924,
    net923,
    net922,
    net921,
    net920,
    net918,
    net917,
    net916,
    net915,
    net914,
    net913,
    net912,
    net911,
    net910,
    net909,
    net907,
    net906,
    net905,
    net904,
    net903,
    net902,
    net901,
    net900,
    net899,
    net898,
    net960,
    net959,
    net958,
    net957,
    net952,
    net941,
    net930,
    net919,
    net908,
    net897}),
    .io_ins_right({\ces_6_6_io_outs_right[63] ,
    \ces_6_6_io_outs_right[62] ,
    \ces_6_6_io_outs_right[61] ,
    \ces_6_6_io_outs_right[60] ,
    \ces_6_6_io_outs_right[59] ,
    \ces_6_6_io_outs_right[58] ,
    \ces_6_6_io_outs_right[57] ,
    \ces_6_6_io_outs_right[56] ,
    \ces_6_6_io_outs_right[55] ,
    \ces_6_6_io_outs_right[54] ,
    \ces_6_6_io_outs_right[53] ,
    \ces_6_6_io_outs_right[52] ,
    \ces_6_6_io_outs_right[51] ,
    \ces_6_6_io_outs_right[50] ,
    \ces_6_6_io_outs_right[49] ,
    \ces_6_6_io_outs_right[48] ,
    \ces_6_6_io_outs_right[47] ,
    \ces_6_6_io_outs_right[46] ,
    \ces_6_6_io_outs_right[45] ,
    \ces_6_6_io_outs_right[44] ,
    \ces_6_6_io_outs_right[43] ,
    \ces_6_6_io_outs_right[42] ,
    \ces_6_6_io_outs_right[41] ,
    \ces_6_6_io_outs_right[40] ,
    \ces_6_6_io_outs_right[39] ,
    \ces_6_6_io_outs_right[38] ,
    \ces_6_6_io_outs_right[37] ,
    \ces_6_6_io_outs_right[36] ,
    \ces_6_6_io_outs_right[35] ,
    \ces_6_6_io_outs_right[34] ,
    \ces_6_6_io_outs_right[33] ,
    \ces_6_6_io_outs_right[32] ,
    \ces_6_6_io_outs_right[31] ,
    \ces_6_6_io_outs_right[30] ,
    \ces_6_6_io_outs_right[29] ,
    \ces_6_6_io_outs_right[28] ,
    \ces_6_6_io_outs_right[27] ,
    \ces_6_6_io_outs_right[26] ,
    \ces_6_6_io_outs_right[25] ,
    \ces_6_6_io_outs_right[24] ,
    \ces_6_6_io_outs_right[23] ,
    \ces_6_6_io_outs_right[22] ,
    \ces_6_6_io_outs_right[21] ,
    \ces_6_6_io_outs_right[20] ,
    \ces_6_6_io_outs_right[19] ,
    \ces_6_6_io_outs_right[18] ,
    \ces_6_6_io_outs_right[17] ,
    \ces_6_6_io_outs_right[16] ,
    \ces_6_6_io_outs_right[15] ,
    \ces_6_6_io_outs_right[14] ,
    \ces_6_6_io_outs_right[13] ,
    \ces_6_6_io_outs_right[12] ,
    \ces_6_6_io_outs_right[11] ,
    \ces_6_6_io_outs_right[10] ,
    \ces_6_6_io_outs_right[9] ,
    \ces_6_6_io_outs_right[8] ,
    \ces_6_6_io_outs_right[7] ,
    \ces_6_6_io_outs_right[6] ,
    \ces_6_6_io_outs_right[5] ,
    \ces_6_6_io_outs_right[4] ,
    \ces_6_6_io_outs_right[3] ,
    \ces_6_6_io_outs_right[2] ,
    \ces_6_6_io_outs_right[1] ,
    \ces_6_6_io_outs_right[0] }),
    .io_ins_up({\ces_5_7_io_outs_up[63] ,
    \ces_5_7_io_outs_up[62] ,
    \ces_5_7_io_outs_up[61] ,
    \ces_5_7_io_outs_up[60] ,
    \ces_5_7_io_outs_up[59] ,
    \ces_5_7_io_outs_up[58] ,
    \ces_5_7_io_outs_up[57] ,
    \ces_5_7_io_outs_up[56] ,
    \ces_5_7_io_outs_up[55] ,
    \ces_5_7_io_outs_up[54] ,
    \ces_5_7_io_outs_up[53] ,
    \ces_5_7_io_outs_up[52] ,
    \ces_5_7_io_outs_up[51] ,
    \ces_5_7_io_outs_up[50] ,
    \ces_5_7_io_outs_up[49] ,
    \ces_5_7_io_outs_up[48] ,
    \ces_5_7_io_outs_up[47] ,
    \ces_5_7_io_outs_up[46] ,
    \ces_5_7_io_outs_up[45] ,
    \ces_5_7_io_outs_up[44] ,
    \ces_5_7_io_outs_up[43] ,
    \ces_5_7_io_outs_up[42] ,
    \ces_5_7_io_outs_up[41] ,
    \ces_5_7_io_outs_up[40] ,
    \ces_5_7_io_outs_up[39] ,
    \ces_5_7_io_outs_up[38] ,
    \ces_5_7_io_outs_up[37] ,
    \ces_5_7_io_outs_up[36] ,
    \ces_5_7_io_outs_up[35] ,
    \ces_5_7_io_outs_up[34] ,
    \ces_5_7_io_outs_up[33] ,
    \ces_5_7_io_outs_up[32] ,
    \ces_5_7_io_outs_up[31] ,
    \ces_5_7_io_outs_up[30] ,
    \ces_5_7_io_outs_up[29] ,
    \ces_5_7_io_outs_up[28] ,
    \ces_5_7_io_outs_up[27] ,
    \ces_5_7_io_outs_up[26] ,
    \ces_5_7_io_outs_up[25] ,
    \ces_5_7_io_outs_up[24] ,
    \ces_5_7_io_outs_up[23] ,
    \ces_5_7_io_outs_up[22] ,
    \ces_5_7_io_outs_up[21] ,
    \ces_5_7_io_outs_up[20] ,
    \ces_5_7_io_outs_up[19] ,
    \ces_5_7_io_outs_up[18] ,
    \ces_5_7_io_outs_up[17] ,
    \ces_5_7_io_outs_up[16] ,
    \ces_5_7_io_outs_up[15] ,
    \ces_5_7_io_outs_up[14] ,
    \ces_5_7_io_outs_up[13] ,
    \ces_5_7_io_outs_up[12] ,
    \ces_5_7_io_outs_up[11] ,
    \ces_5_7_io_outs_up[10] ,
    \ces_5_7_io_outs_up[9] ,
    \ces_5_7_io_outs_up[8] ,
    \ces_5_7_io_outs_up[7] ,
    \ces_5_7_io_outs_up[6] ,
    \ces_5_7_io_outs_up[5] ,
    \ces_5_7_io_outs_up[4] ,
    \ces_5_7_io_outs_up[3] ,
    \ces_5_7_io_outs_up[2] ,
    \ces_5_7_io_outs_up[1] ,
    \ces_5_7_io_outs_up[0] }),
    .io_outs_down({\ces_5_7_io_ins_down[63] ,
    \ces_5_7_io_ins_down[62] ,
    \ces_5_7_io_ins_down[61] ,
    \ces_5_7_io_ins_down[60] ,
    \ces_5_7_io_ins_down[59] ,
    \ces_5_7_io_ins_down[58] ,
    \ces_5_7_io_ins_down[57] ,
    \ces_5_7_io_ins_down[56] ,
    \ces_5_7_io_ins_down[55] ,
    \ces_5_7_io_ins_down[54] ,
    \ces_5_7_io_ins_down[53] ,
    \ces_5_7_io_ins_down[52] ,
    \ces_5_7_io_ins_down[51] ,
    \ces_5_7_io_ins_down[50] ,
    \ces_5_7_io_ins_down[49] ,
    \ces_5_7_io_ins_down[48] ,
    \ces_5_7_io_ins_down[47] ,
    \ces_5_7_io_ins_down[46] ,
    \ces_5_7_io_ins_down[45] ,
    \ces_5_7_io_ins_down[44] ,
    \ces_5_7_io_ins_down[43] ,
    \ces_5_7_io_ins_down[42] ,
    \ces_5_7_io_ins_down[41] ,
    \ces_5_7_io_ins_down[40] ,
    \ces_5_7_io_ins_down[39] ,
    \ces_5_7_io_ins_down[38] ,
    \ces_5_7_io_ins_down[37] ,
    \ces_5_7_io_ins_down[36] ,
    \ces_5_7_io_ins_down[35] ,
    \ces_5_7_io_ins_down[34] ,
    \ces_5_7_io_ins_down[33] ,
    \ces_5_7_io_ins_down[32] ,
    \ces_5_7_io_ins_down[31] ,
    \ces_5_7_io_ins_down[30] ,
    \ces_5_7_io_ins_down[29] ,
    \ces_5_7_io_ins_down[28] ,
    \ces_5_7_io_ins_down[27] ,
    \ces_5_7_io_ins_down[26] ,
    \ces_5_7_io_ins_down[25] ,
    \ces_5_7_io_ins_down[24] ,
    \ces_5_7_io_ins_down[23] ,
    \ces_5_7_io_ins_down[22] ,
    \ces_5_7_io_ins_down[21] ,
    \ces_5_7_io_ins_down[20] ,
    \ces_5_7_io_ins_down[19] ,
    \ces_5_7_io_ins_down[18] ,
    \ces_5_7_io_ins_down[17] ,
    \ces_5_7_io_ins_down[16] ,
    \ces_5_7_io_ins_down[15] ,
    \ces_5_7_io_ins_down[14] ,
    \ces_5_7_io_ins_down[13] ,
    \ces_5_7_io_ins_down[12] ,
    \ces_5_7_io_ins_down[11] ,
    \ces_5_7_io_ins_down[10] ,
    \ces_5_7_io_ins_down[9] ,
    \ces_5_7_io_ins_down[8] ,
    \ces_5_7_io_ins_down[7] ,
    \ces_5_7_io_ins_down[6] ,
    \ces_5_7_io_ins_down[5] ,
    \ces_5_7_io_ins_down[4] ,
    \ces_5_7_io_ins_down[3] ,
    \ces_5_7_io_ins_down[2] ,
    \ces_5_7_io_ins_down[1] ,
    \ces_5_7_io_ins_down[0] }),
    .io_outs_left({\ces_6_6_io_ins_left[63] ,
    \ces_6_6_io_ins_left[62] ,
    \ces_6_6_io_ins_left[61] ,
    \ces_6_6_io_ins_left[60] ,
    \ces_6_6_io_ins_left[59] ,
    \ces_6_6_io_ins_left[58] ,
    \ces_6_6_io_ins_left[57] ,
    \ces_6_6_io_ins_left[56] ,
    \ces_6_6_io_ins_left[55] ,
    \ces_6_6_io_ins_left[54] ,
    \ces_6_6_io_ins_left[53] ,
    \ces_6_6_io_ins_left[52] ,
    \ces_6_6_io_ins_left[51] ,
    \ces_6_6_io_ins_left[50] ,
    \ces_6_6_io_ins_left[49] ,
    \ces_6_6_io_ins_left[48] ,
    \ces_6_6_io_ins_left[47] ,
    \ces_6_6_io_ins_left[46] ,
    \ces_6_6_io_ins_left[45] ,
    \ces_6_6_io_ins_left[44] ,
    \ces_6_6_io_ins_left[43] ,
    \ces_6_6_io_ins_left[42] ,
    \ces_6_6_io_ins_left[41] ,
    \ces_6_6_io_ins_left[40] ,
    \ces_6_6_io_ins_left[39] ,
    \ces_6_6_io_ins_left[38] ,
    \ces_6_6_io_ins_left[37] ,
    \ces_6_6_io_ins_left[36] ,
    \ces_6_6_io_ins_left[35] ,
    \ces_6_6_io_ins_left[34] ,
    \ces_6_6_io_ins_left[33] ,
    \ces_6_6_io_ins_left[32] ,
    \ces_6_6_io_ins_left[31] ,
    \ces_6_6_io_ins_left[30] ,
    \ces_6_6_io_ins_left[29] ,
    \ces_6_6_io_ins_left[28] ,
    \ces_6_6_io_ins_left[27] ,
    \ces_6_6_io_ins_left[26] ,
    \ces_6_6_io_ins_left[25] ,
    \ces_6_6_io_ins_left[24] ,
    \ces_6_6_io_ins_left[23] ,
    \ces_6_6_io_ins_left[22] ,
    \ces_6_6_io_ins_left[21] ,
    \ces_6_6_io_ins_left[20] ,
    \ces_6_6_io_ins_left[19] ,
    \ces_6_6_io_ins_left[18] ,
    \ces_6_6_io_ins_left[17] ,
    \ces_6_6_io_ins_left[16] ,
    \ces_6_6_io_ins_left[15] ,
    \ces_6_6_io_ins_left[14] ,
    \ces_6_6_io_ins_left[13] ,
    \ces_6_6_io_ins_left[12] ,
    \ces_6_6_io_ins_left[11] ,
    \ces_6_6_io_ins_left[10] ,
    \ces_6_6_io_ins_left[9] ,
    \ces_6_6_io_ins_left[8] ,
    \ces_6_6_io_ins_left[7] ,
    \ces_6_6_io_ins_left[6] ,
    \ces_6_6_io_ins_left[5] ,
    \ces_6_6_io_ins_left[4] ,
    \ces_6_6_io_ins_left[3] ,
    \ces_6_6_io_ins_left[2] ,
    \ces_6_6_io_ins_left[1] ,
    \ces_6_6_io_ins_left[0] }),
    .io_outs_right({net3580,
    net3579,
    net3578,
    net3577,
    net3575,
    net3574,
    net3573,
    net3572,
    net3571,
    net3570,
    net3569,
    net3568,
    net3567,
    net3566,
    net3564,
    net3563,
    net3562,
    net3561,
    net3560,
    net3559,
    net3558,
    net3557,
    net3556,
    net3555,
    net3553,
    net3552,
    net3551,
    net3550,
    net3549,
    net3548,
    net3547,
    net3546,
    net3545,
    net3544,
    net3542,
    net3541,
    net3540,
    net3539,
    net3538,
    net3537,
    net3536,
    net3535,
    net3534,
    net3533,
    net3531,
    net3530,
    net3529,
    net3528,
    net3527,
    net3526,
    net3525,
    net3524,
    net3523,
    net3522,
    net3584,
    net3583,
    net3582,
    net3581,
    net3576,
    net3565,
    net3554,
    net3543,
    net3532,
    net3521}),
    .io_outs_up({\ces_6_7_io_outs_up[63] ,
    \ces_6_7_io_outs_up[62] ,
    \ces_6_7_io_outs_up[61] ,
    \ces_6_7_io_outs_up[60] ,
    \ces_6_7_io_outs_up[59] ,
    \ces_6_7_io_outs_up[58] ,
    \ces_6_7_io_outs_up[57] ,
    \ces_6_7_io_outs_up[56] ,
    \ces_6_7_io_outs_up[55] ,
    \ces_6_7_io_outs_up[54] ,
    \ces_6_7_io_outs_up[53] ,
    \ces_6_7_io_outs_up[52] ,
    \ces_6_7_io_outs_up[51] ,
    \ces_6_7_io_outs_up[50] ,
    \ces_6_7_io_outs_up[49] ,
    \ces_6_7_io_outs_up[48] ,
    \ces_6_7_io_outs_up[47] ,
    \ces_6_7_io_outs_up[46] ,
    \ces_6_7_io_outs_up[45] ,
    \ces_6_7_io_outs_up[44] ,
    \ces_6_7_io_outs_up[43] ,
    \ces_6_7_io_outs_up[42] ,
    \ces_6_7_io_outs_up[41] ,
    \ces_6_7_io_outs_up[40] ,
    \ces_6_7_io_outs_up[39] ,
    \ces_6_7_io_outs_up[38] ,
    \ces_6_7_io_outs_up[37] ,
    \ces_6_7_io_outs_up[36] ,
    \ces_6_7_io_outs_up[35] ,
    \ces_6_7_io_outs_up[34] ,
    \ces_6_7_io_outs_up[33] ,
    \ces_6_7_io_outs_up[32] ,
    \ces_6_7_io_outs_up[31] ,
    \ces_6_7_io_outs_up[30] ,
    \ces_6_7_io_outs_up[29] ,
    \ces_6_7_io_outs_up[28] ,
    \ces_6_7_io_outs_up[27] ,
    \ces_6_7_io_outs_up[26] ,
    \ces_6_7_io_outs_up[25] ,
    \ces_6_7_io_outs_up[24] ,
    \ces_6_7_io_outs_up[23] ,
    \ces_6_7_io_outs_up[22] ,
    \ces_6_7_io_outs_up[21] ,
    \ces_6_7_io_outs_up[20] ,
    \ces_6_7_io_outs_up[19] ,
    \ces_6_7_io_outs_up[18] ,
    \ces_6_7_io_outs_up[17] ,
    \ces_6_7_io_outs_up[16] ,
    \ces_6_7_io_outs_up[15] ,
    \ces_6_7_io_outs_up[14] ,
    \ces_6_7_io_outs_up[13] ,
    \ces_6_7_io_outs_up[12] ,
    \ces_6_7_io_outs_up[11] ,
    \ces_6_7_io_outs_up[10] ,
    \ces_6_7_io_outs_up[9] ,
    \ces_6_7_io_outs_up[8] ,
    \ces_6_7_io_outs_up[7] ,
    \ces_6_7_io_outs_up[6] ,
    \ces_6_7_io_outs_up[5] ,
    \ces_6_7_io_outs_up[4] ,
    \ces_6_7_io_outs_up[3] ,
    \ces_6_7_io_outs_up[2] ,
    \ces_6_7_io_outs_up[1] ,
    \ces_6_7_io_outs_up[0] }));
 Element ces_7_0 (.clock(clknet_3_5_0_clock),
    .io_lsbIns_1(net4210),
    .io_lsbIns_2(net4211),
    .io_lsbIns_3(net4212),
    .io_lsbIns_4(net4213),
    .io_lsbIns_5(net4214),
    .io_lsbIns_6(net4215),
    .io_lsbIns_7(net4216),
    .io_lsbOuts_0(ces_7_0_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_0_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_0_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_0_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_0_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_0_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_0_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_0_io_lsbOuts_7),
    .io_ins_down({net60,
    net59,
    net58,
    net57,
    net55,
    net54,
    net53,
    net52,
    net51,
    net50,
    net49,
    net48,
    net47,
    net46,
    net44,
    net43,
    net42,
    net41,
    net40,
    net39,
    net38,
    net37,
    net36,
    net35,
    net33,
    net32,
    net31,
    net30,
    net29,
    net28,
    net27,
    net26,
    net25,
    net24,
    net22,
    net21,
    net20,
    net19,
    net18,
    net17,
    net16,
    net15,
    net14,
    net13,
    net11,
    net10,
    net9,
    net8,
    net7,
    net6,
    net5,
    net4,
    net3,
    net2,
    net64,
    net63,
    net62,
    net61,
    net56,
    net45,
    net34,
    net23,
    net12,
    net1}),
    .io_ins_left({\ces_7_0_io_ins_left[63] ,
    \ces_7_0_io_ins_left[62] ,
    \ces_7_0_io_ins_left[61] ,
    \ces_7_0_io_ins_left[60] ,
    \ces_7_0_io_ins_left[59] ,
    \ces_7_0_io_ins_left[58] ,
    \ces_7_0_io_ins_left[57] ,
    \ces_7_0_io_ins_left[56] ,
    \ces_7_0_io_ins_left[55] ,
    \ces_7_0_io_ins_left[54] ,
    \ces_7_0_io_ins_left[53] ,
    \ces_7_0_io_ins_left[52] ,
    \ces_7_0_io_ins_left[51] ,
    \ces_7_0_io_ins_left[50] ,
    \ces_7_0_io_ins_left[49] ,
    \ces_7_0_io_ins_left[48] ,
    \ces_7_0_io_ins_left[47] ,
    \ces_7_0_io_ins_left[46] ,
    \ces_7_0_io_ins_left[45] ,
    \ces_7_0_io_ins_left[44] ,
    \ces_7_0_io_ins_left[43] ,
    \ces_7_0_io_ins_left[42] ,
    \ces_7_0_io_ins_left[41] ,
    \ces_7_0_io_ins_left[40] ,
    \ces_7_0_io_ins_left[39] ,
    \ces_7_0_io_ins_left[38] ,
    \ces_7_0_io_ins_left[37] ,
    \ces_7_0_io_ins_left[36] ,
    \ces_7_0_io_ins_left[35] ,
    \ces_7_0_io_ins_left[34] ,
    \ces_7_0_io_ins_left[33] ,
    \ces_7_0_io_ins_left[32] ,
    \ces_7_0_io_ins_left[31] ,
    \ces_7_0_io_ins_left[30] ,
    \ces_7_0_io_ins_left[29] ,
    \ces_7_0_io_ins_left[28] ,
    \ces_7_0_io_ins_left[27] ,
    \ces_7_0_io_ins_left[26] ,
    \ces_7_0_io_ins_left[25] ,
    \ces_7_0_io_ins_left[24] ,
    \ces_7_0_io_ins_left[23] ,
    \ces_7_0_io_ins_left[22] ,
    \ces_7_0_io_ins_left[21] ,
    \ces_7_0_io_ins_left[20] ,
    \ces_7_0_io_ins_left[19] ,
    \ces_7_0_io_ins_left[18] ,
    \ces_7_0_io_ins_left[17] ,
    \ces_7_0_io_ins_left[16] ,
    \ces_7_0_io_ins_left[15] ,
    \ces_7_0_io_ins_left[14] ,
    \ces_7_0_io_ins_left[13] ,
    \ces_7_0_io_ins_left[12] ,
    \ces_7_0_io_ins_left[11] ,
    \ces_7_0_io_ins_left[10] ,
    \ces_7_0_io_ins_left[9] ,
    \ces_7_0_io_ins_left[8] ,
    \ces_7_0_io_ins_left[7] ,
    \ces_7_0_io_ins_left[6] ,
    \ces_7_0_io_ins_left[5] ,
    \ces_7_0_io_ins_left[4] ,
    \ces_7_0_io_ins_left[3] ,
    \ces_7_0_io_ins_left[2] ,
    \ces_7_0_io_ins_left[1] ,
    \ces_7_0_io_ins_left[0] }),
    .io_ins_right({net1532,
    net1531,
    net1530,
    net1529,
    net1527,
    net1526,
    net1525,
    net1524,
    net1523,
    net1522,
    net1521,
    net1520,
    net1519,
    net1518,
    net1516,
    net1515,
    net1514,
    net1513,
    net1512,
    net1511,
    net1510,
    net1509,
    net1508,
    net1507,
    net1505,
    net1504,
    net1503,
    net1502,
    net1501,
    net1500,
    net1499,
    net1498,
    net1497,
    net1496,
    net1494,
    net1493,
    net1492,
    net1491,
    net1490,
    net1489,
    net1488,
    net1487,
    net1486,
    net1485,
    net1483,
    net1482,
    net1481,
    net1480,
    net1479,
    net1478,
    net1477,
    net1476,
    net1475,
    net1474,
    net1536,
    net1535,
    net1534,
    net1533,
    net1528,
    net1517,
    net1506,
    net1495,
    net1484,
    net1473}),
    .io_ins_up({\ces_6_0_io_outs_up[63] ,
    \ces_6_0_io_outs_up[62] ,
    \ces_6_0_io_outs_up[61] ,
    \ces_6_0_io_outs_up[60] ,
    \ces_6_0_io_outs_up[59] ,
    \ces_6_0_io_outs_up[58] ,
    \ces_6_0_io_outs_up[57] ,
    \ces_6_0_io_outs_up[56] ,
    \ces_6_0_io_outs_up[55] ,
    \ces_6_0_io_outs_up[54] ,
    \ces_6_0_io_outs_up[53] ,
    \ces_6_0_io_outs_up[52] ,
    \ces_6_0_io_outs_up[51] ,
    \ces_6_0_io_outs_up[50] ,
    \ces_6_0_io_outs_up[49] ,
    \ces_6_0_io_outs_up[48] ,
    \ces_6_0_io_outs_up[47] ,
    \ces_6_0_io_outs_up[46] ,
    \ces_6_0_io_outs_up[45] ,
    \ces_6_0_io_outs_up[44] ,
    \ces_6_0_io_outs_up[43] ,
    \ces_6_0_io_outs_up[42] ,
    \ces_6_0_io_outs_up[41] ,
    \ces_6_0_io_outs_up[40] ,
    \ces_6_0_io_outs_up[39] ,
    \ces_6_0_io_outs_up[38] ,
    \ces_6_0_io_outs_up[37] ,
    \ces_6_0_io_outs_up[36] ,
    \ces_6_0_io_outs_up[35] ,
    \ces_6_0_io_outs_up[34] ,
    \ces_6_0_io_outs_up[33] ,
    \ces_6_0_io_outs_up[32] ,
    \ces_6_0_io_outs_up[31] ,
    \ces_6_0_io_outs_up[30] ,
    \ces_6_0_io_outs_up[29] ,
    \ces_6_0_io_outs_up[28] ,
    \ces_6_0_io_outs_up[27] ,
    \ces_6_0_io_outs_up[26] ,
    \ces_6_0_io_outs_up[25] ,
    \ces_6_0_io_outs_up[24] ,
    \ces_6_0_io_outs_up[23] ,
    \ces_6_0_io_outs_up[22] ,
    \ces_6_0_io_outs_up[21] ,
    \ces_6_0_io_outs_up[20] ,
    \ces_6_0_io_outs_up[19] ,
    \ces_6_0_io_outs_up[18] ,
    \ces_6_0_io_outs_up[17] ,
    \ces_6_0_io_outs_up[16] ,
    \ces_6_0_io_outs_up[15] ,
    \ces_6_0_io_outs_up[14] ,
    \ces_6_0_io_outs_up[13] ,
    \ces_6_0_io_outs_up[12] ,
    \ces_6_0_io_outs_up[11] ,
    \ces_6_0_io_outs_up[10] ,
    \ces_6_0_io_outs_up[9] ,
    \ces_6_0_io_outs_up[8] ,
    \ces_6_0_io_outs_up[7] ,
    \ces_6_0_io_outs_up[6] ,
    \ces_6_0_io_outs_up[5] ,
    \ces_6_0_io_outs_up[4] ,
    \ces_6_0_io_outs_up[3] ,
    \ces_6_0_io_outs_up[2] ,
    \ces_6_0_io_outs_up[1] ,
    \ces_6_0_io_outs_up[0] }),
    .io_outs_down({\ces_6_0_io_ins_down[63] ,
    \ces_6_0_io_ins_down[62] ,
    \ces_6_0_io_ins_down[61] ,
    \ces_6_0_io_ins_down[60] ,
    \ces_6_0_io_ins_down[59] ,
    \ces_6_0_io_ins_down[58] ,
    \ces_6_0_io_ins_down[57] ,
    \ces_6_0_io_ins_down[56] ,
    \ces_6_0_io_ins_down[55] ,
    \ces_6_0_io_ins_down[54] ,
    \ces_6_0_io_ins_down[53] ,
    \ces_6_0_io_ins_down[52] ,
    \ces_6_0_io_ins_down[51] ,
    \ces_6_0_io_ins_down[50] ,
    \ces_6_0_io_ins_down[49] ,
    \ces_6_0_io_ins_down[48] ,
    \ces_6_0_io_ins_down[47] ,
    \ces_6_0_io_ins_down[46] ,
    \ces_6_0_io_ins_down[45] ,
    \ces_6_0_io_ins_down[44] ,
    \ces_6_0_io_ins_down[43] ,
    \ces_6_0_io_ins_down[42] ,
    \ces_6_0_io_ins_down[41] ,
    \ces_6_0_io_ins_down[40] ,
    \ces_6_0_io_ins_down[39] ,
    \ces_6_0_io_ins_down[38] ,
    \ces_6_0_io_ins_down[37] ,
    \ces_6_0_io_ins_down[36] ,
    \ces_6_0_io_ins_down[35] ,
    \ces_6_0_io_ins_down[34] ,
    \ces_6_0_io_ins_down[33] ,
    \ces_6_0_io_ins_down[32] ,
    \ces_6_0_io_ins_down[31] ,
    \ces_6_0_io_ins_down[30] ,
    \ces_6_0_io_ins_down[29] ,
    \ces_6_0_io_ins_down[28] ,
    \ces_6_0_io_ins_down[27] ,
    \ces_6_0_io_ins_down[26] ,
    \ces_6_0_io_ins_down[25] ,
    \ces_6_0_io_ins_down[24] ,
    \ces_6_0_io_ins_down[23] ,
    \ces_6_0_io_ins_down[22] ,
    \ces_6_0_io_ins_down[21] ,
    \ces_6_0_io_ins_down[20] ,
    \ces_6_0_io_ins_down[19] ,
    \ces_6_0_io_ins_down[18] ,
    \ces_6_0_io_ins_down[17] ,
    \ces_6_0_io_ins_down[16] ,
    \ces_6_0_io_ins_down[15] ,
    \ces_6_0_io_ins_down[14] ,
    \ces_6_0_io_ins_down[13] ,
    \ces_6_0_io_ins_down[12] ,
    \ces_6_0_io_ins_down[11] ,
    \ces_6_0_io_ins_down[10] ,
    \ces_6_0_io_ins_down[9] ,
    \ces_6_0_io_ins_down[8] ,
    \ces_6_0_io_ins_down[7] ,
    \ces_6_0_io_ins_down[6] ,
    \ces_6_0_io_ins_down[5] ,
    \ces_6_0_io_ins_down[4] ,
    \ces_6_0_io_ins_down[3] ,
    \ces_6_0_io_ins_down[2] ,
    \ces_6_0_io_ins_down[1] ,
    \ces_6_0_io_ins_down[0] }),
    .io_outs_left({net3132,
    net3131,
    net3130,
    net3129,
    net3127,
    net3126,
    net3125,
    net3124,
    net3123,
    net3122,
    net3121,
    net3120,
    net3119,
    net3118,
    net3116,
    net3115,
    net3114,
    net3113,
    net3112,
    net3111,
    net3110,
    net3109,
    net3108,
    net3107,
    net3105,
    net3104,
    net3103,
    net3102,
    net3101,
    net3100,
    net3099,
    net3098,
    net3097,
    net3096,
    net3094,
    net3093,
    net3092,
    net3091,
    net3090,
    net3089,
    net3088,
    net3087,
    net3086,
    net3085,
    net3083,
    net3082,
    net3081,
    net3080,
    net3079,
    net3078,
    net3077,
    net3076,
    net3075,
    net3074,
    net3136,
    net3135,
    net3134,
    net3133,
    net3128,
    net3117,
    net3106,
    net3095,
    net3084,
    net3073}),
    .io_outs_right({\ces_7_0_io_outs_right[63] ,
    \ces_7_0_io_outs_right[62] ,
    \ces_7_0_io_outs_right[61] ,
    \ces_7_0_io_outs_right[60] ,
    \ces_7_0_io_outs_right[59] ,
    \ces_7_0_io_outs_right[58] ,
    \ces_7_0_io_outs_right[57] ,
    \ces_7_0_io_outs_right[56] ,
    \ces_7_0_io_outs_right[55] ,
    \ces_7_0_io_outs_right[54] ,
    \ces_7_0_io_outs_right[53] ,
    \ces_7_0_io_outs_right[52] ,
    \ces_7_0_io_outs_right[51] ,
    \ces_7_0_io_outs_right[50] ,
    \ces_7_0_io_outs_right[49] ,
    \ces_7_0_io_outs_right[48] ,
    \ces_7_0_io_outs_right[47] ,
    \ces_7_0_io_outs_right[46] ,
    \ces_7_0_io_outs_right[45] ,
    \ces_7_0_io_outs_right[44] ,
    \ces_7_0_io_outs_right[43] ,
    \ces_7_0_io_outs_right[42] ,
    \ces_7_0_io_outs_right[41] ,
    \ces_7_0_io_outs_right[40] ,
    \ces_7_0_io_outs_right[39] ,
    \ces_7_0_io_outs_right[38] ,
    \ces_7_0_io_outs_right[37] ,
    \ces_7_0_io_outs_right[36] ,
    \ces_7_0_io_outs_right[35] ,
    \ces_7_0_io_outs_right[34] ,
    \ces_7_0_io_outs_right[33] ,
    \ces_7_0_io_outs_right[32] ,
    \ces_7_0_io_outs_right[31] ,
    \ces_7_0_io_outs_right[30] ,
    \ces_7_0_io_outs_right[29] ,
    \ces_7_0_io_outs_right[28] ,
    \ces_7_0_io_outs_right[27] ,
    \ces_7_0_io_outs_right[26] ,
    \ces_7_0_io_outs_right[25] ,
    \ces_7_0_io_outs_right[24] ,
    \ces_7_0_io_outs_right[23] ,
    \ces_7_0_io_outs_right[22] ,
    \ces_7_0_io_outs_right[21] ,
    \ces_7_0_io_outs_right[20] ,
    \ces_7_0_io_outs_right[19] ,
    \ces_7_0_io_outs_right[18] ,
    \ces_7_0_io_outs_right[17] ,
    \ces_7_0_io_outs_right[16] ,
    \ces_7_0_io_outs_right[15] ,
    \ces_7_0_io_outs_right[14] ,
    \ces_7_0_io_outs_right[13] ,
    \ces_7_0_io_outs_right[12] ,
    \ces_7_0_io_outs_right[11] ,
    \ces_7_0_io_outs_right[10] ,
    \ces_7_0_io_outs_right[9] ,
    \ces_7_0_io_outs_right[8] ,
    \ces_7_0_io_outs_right[7] ,
    \ces_7_0_io_outs_right[6] ,
    \ces_7_0_io_outs_right[5] ,
    \ces_7_0_io_outs_right[4] ,
    \ces_7_0_io_outs_right[3] ,
    \ces_7_0_io_outs_right[2] ,
    \ces_7_0_io_outs_right[1] ,
    \ces_7_0_io_outs_right[0] }),
    .io_outs_up({net3708,
    net3707,
    net3706,
    net3705,
    net3703,
    net3702,
    net3701,
    net3700,
    net3699,
    net3698,
    net3697,
    net3696,
    net3695,
    net3694,
    net3692,
    net3691,
    net3690,
    net3689,
    net3688,
    net3687,
    net3686,
    net3685,
    net3684,
    net3683,
    net3681,
    net3680,
    net3679,
    net3678,
    net3677,
    net3676,
    net3675,
    net3674,
    net3673,
    net3672,
    net3670,
    net3669,
    net3668,
    net3667,
    net3666,
    net3665,
    net3664,
    net3663,
    net3662,
    net3661,
    net3659,
    net3658,
    net3657,
    net3656,
    net3655,
    net3654,
    net3653,
    net3652,
    net3651,
    net3650,
    net3712,
    net3711,
    net3710,
    net3709,
    net3704,
    net3693,
    net3682,
    net3671,
    net3660,
    net3649}));
 Element ces_7_1 (.clock(clknet_3_5_0_clock),
    .io_lsbIns_1(ces_7_0_io_lsbOuts_1),
    .io_lsbIns_2(ces_7_0_io_lsbOuts_2),
    .io_lsbIns_3(ces_7_0_io_lsbOuts_3),
    .io_lsbIns_4(ces_7_0_io_lsbOuts_4),
    .io_lsbIns_5(ces_7_0_io_lsbOuts_5),
    .io_lsbIns_6(ces_7_0_io_lsbOuts_6),
    .io_lsbIns_7(ces_7_0_io_lsbOuts_7),
    .io_lsbOuts_0(ces_7_1_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_1_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_1_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_1_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_1_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_1_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_1_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_1_io_lsbOuts_7),
    .io_ins_down({net124,
    net123,
    net122,
    net121,
    net119,
    net118,
    net117,
    net116,
    net115,
    net114,
    net113,
    net112,
    net111,
    net110,
    net108,
    net107,
    net106,
    net105,
    net104,
    net103,
    net102,
    net101,
    net100,
    net99,
    net97,
    net96,
    net95,
    net94,
    net93,
    net92,
    net91,
    net90,
    net89,
    net88,
    net86,
    net85,
    net84,
    net83,
    net82,
    net81,
    net80,
    net79,
    net78,
    net77,
    net75,
    net74,
    net73,
    net72,
    net71,
    net70,
    net69,
    net68,
    net67,
    net66,
    net128,
    net127,
    net126,
    net125,
    net120,
    net109,
    net98,
    net87,
    net76,
    net65}),
    .io_ins_left({\ces_7_1_io_ins_left[63] ,
    \ces_7_1_io_ins_left[62] ,
    \ces_7_1_io_ins_left[61] ,
    \ces_7_1_io_ins_left[60] ,
    \ces_7_1_io_ins_left[59] ,
    \ces_7_1_io_ins_left[58] ,
    \ces_7_1_io_ins_left[57] ,
    \ces_7_1_io_ins_left[56] ,
    \ces_7_1_io_ins_left[55] ,
    \ces_7_1_io_ins_left[54] ,
    \ces_7_1_io_ins_left[53] ,
    \ces_7_1_io_ins_left[52] ,
    \ces_7_1_io_ins_left[51] ,
    \ces_7_1_io_ins_left[50] ,
    \ces_7_1_io_ins_left[49] ,
    \ces_7_1_io_ins_left[48] ,
    \ces_7_1_io_ins_left[47] ,
    \ces_7_1_io_ins_left[46] ,
    \ces_7_1_io_ins_left[45] ,
    \ces_7_1_io_ins_left[44] ,
    \ces_7_1_io_ins_left[43] ,
    \ces_7_1_io_ins_left[42] ,
    \ces_7_1_io_ins_left[41] ,
    \ces_7_1_io_ins_left[40] ,
    \ces_7_1_io_ins_left[39] ,
    \ces_7_1_io_ins_left[38] ,
    \ces_7_1_io_ins_left[37] ,
    \ces_7_1_io_ins_left[36] ,
    \ces_7_1_io_ins_left[35] ,
    \ces_7_1_io_ins_left[34] ,
    \ces_7_1_io_ins_left[33] ,
    \ces_7_1_io_ins_left[32] ,
    \ces_7_1_io_ins_left[31] ,
    \ces_7_1_io_ins_left[30] ,
    \ces_7_1_io_ins_left[29] ,
    \ces_7_1_io_ins_left[28] ,
    \ces_7_1_io_ins_left[27] ,
    \ces_7_1_io_ins_left[26] ,
    \ces_7_1_io_ins_left[25] ,
    \ces_7_1_io_ins_left[24] ,
    \ces_7_1_io_ins_left[23] ,
    \ces_7_1_io_ins_left[22] ,
    \ces_7_1_io_ins_left[21] ,
    \ces_7_1_io_ins_left[20] ,
    \ces_7_1_io_ins_left[19] ,
    \ces_7_1_io_ins_left[18] ,
    \ces_7_1_io_ins_left[17] ,
    \ces_7_1_io_ins_left[16] ,
    \ces_7_1_io_ins_left[15] ,
    \ces_7_1_io_ins_left[14] ,
    \ces_7_1_io_ins_left[13] ,
    \ces_7_1_io_ins_left[12] ,
    \ces_7_1_io_ins_left[11] ,
    \ces_7_1_io_ins_left[10] ,
    \ces_7_1_io_ins_left[9] ,
    \ces_7_1_io_ins_left[8] ,
    \ces_7_1_io_ins_left[7] ,
    \ces_7_1_io_ins_left[6] ,
    \ces_7_1_io_ins_left[5] ,
    \ces_7_1_io_ins_left[4] ,
    \ces_7_1_io_ins_left[3] ,
    \ces_7_1_io_ins_left[2] ,
    \ces_7_1_io_ins_left[1] ,
    \ces_7_1_io_ins_left[0] }),
    .io_ins_right({\ces_7_0_io_outs_right[63] ,
    \ces_7_0_io_outs_right[62] ,
    \ces_7_0_io_outs_right[61] ,
    \ces_7_0_io_outs_right[60] ,
    \ces_7_0_io_outs_right[59] ,
    \ces_7_0_io_outs_right[58] ,
    \ces_7_0_io_outs_right[57] ,
    \ces_7_0_io_outs_right[56] ,
    \ces_7_0_io_outs_right[55] ,
    \ces_7_0_io_outs_right[54] ,
    \ces_7_0_io_outs_right[53] ,
    \ces_7_0_io_outs_right[52] ,
    \ces_7_0_io_outs_right[51] ,
    \ces_7_0_io_outs_right[50] ,
    \ces_7_0_io_outs_right[49] ,
    \ces_7_0_io_outs_right[48] ,
    \ces_7_0_io_outs_right[47] ,
    \ces_7_0_io_outs_right[46] ,
    \ces_7_0_io_outs_right[45] ,
    \ces_7_0_io_outs_right[44] ,
    \ces_7_0_io_outs_right[43] ,
    \ces_7_0_io_outs_right[42] ,
    \ces_7_0_io_outs_right[41] ,
    \ces_7_0_io_outs_right[40] ,
    \ces_7_0_io_outs_right[39] ,
    \ces_7_0_io_outs_right[38] ,
    \ces_7_0_io_outs_right[37] ,
    \ces_7_0_io_outs_right[36] ,
    \ces_7_0_io_outs_right[35] ,
    \ces_7_0_io_outs_right[34] ,
    \ces_7_0_io_outs_right[33] ,
    \ces_7_0_io_outs_right[32] ,
    \ces_7_0_io_outs_right[31] ,
    \ces_7_0_io_outs_right[30] ,
    \ces_7_0_io_outs_right[29] ,
    \ces_7_0_io_outs_right[28] ,
    \ces_7_0_io_outs_right[27] ,
    \ces_7_0_io_outs_right[26] ,
    \ces_7_0_io_outs_right[25] ,
    \ces_7_0_io_outs_right[24] ,
    \ces_7_0_io_outs_right[23] ,
    \ces_7_0_io_outs_right[22] ,
    \ces_7_0_io_outs_right[21] ,
    \ces_7_0_io_outs_right[20] ,
    \ces_7_0_io_outs_right[19] ,
    \ces_7_0_io_outs_right[18] ,
    \ces_7_0_io_outs_right[17] ,
    \ces_7_0_io_outs_right[16] ,
    \ces_7_0_io_outs_right[15] ,
    \ces_7_0_io_outs_right[14] ,
    \ces_7_0_io_outs_right[13] ,
    \ces_7_0_io_outs_right[12] ,
    \ces_7_0_io_outs_right[11] ,
    \ces_7_0_io_outs_right[10] ,
    \ces_7_0_io_outs_right[9] ,
    \ces_7_0_io_outs_right[8] ,
    \ces_7_0_io_outs_right[7] ,
    \ces_7_0_io_outs_right[6] ,
    \ces_7_0_io_outs_right[5] ,
    \ces_7_0_io_outs_right[4] ,
    \ces_7_0_io_outs_right[3] ,
    \ces_7_0_io_outs_right[2] ,
    \ces_7_0_io_outs_right[1] ,
    \ces_7_0_io_outs_right[0] }),
    .io_ins_up({\ces_6_1_io_outs_up[63] ,
    \ces_6_1_io_outs_up[62] ,
    \ces_6_1_io_outs_up[61] ,
    \ces_6_1_io_outs_up[60] ,
    \ces_6_1_io_outs_up[59] ,
    \ces_6_1_io_outs_up[58] ,
    \ces_6_1_io_outs_up[57] ,
    \ces_6_1_io_outs_up[56] ,
    \ces_6_1_io_outs_up[55] ,
    \ces_6_1_io_outs_up[54] ,
    \ces_6_1_io_outs_up[53] ,
    \ces_6_1_io_outs_up[52] ,
    \ces_6_1_io_outs_up[51] ,
    \ces_6_1_io_outs_up[50] ,
    \ces_6_1_io_outs_up[49] ,
    \ces_6_1_io_outs_up[48] ,
    \ces_6_1_io_outs_up[47] ,
    \ces_6_1_io_outs_up[46] ,
    \ces_6_1_io_outs_up[45] ,
    \ces_6_1_io_outs_up[44] ,
    \ces_6_1_io_outs_up[43] ,
    \ces_6_1_io_outs_up[42] ,
    \ces_6_1_io_outs_up[41] ,
    \ces_6_1_io_outs_up[40] ,
    \ces_6_1_io_outs_up[39] ,
    \ces_6_1_io_outs_up[38] ,
    \ces_6_1_io_outs_up[37] ,
    \ces_6_1_io_outs_up[36] ,
    \ces_6_1_io_outs_up[35] ,
    \ces_6_1_io_outs_up[34] ,
    \ces_6_1_io_outs_up[33] ,
    \ces_6_1_io_outs_up[32] ,
    \ces_6_1_io_outs_up[31] ,
    \ces_6_1_io_outs_up[30] ,
    \ces_6_1_io_outs_up[29] ,
    \ces_6_1_io_outs_up[28] ,
    \ces_6_1_io_outs_up[27] ,
    \ces_6_1_io_outs_up[26] ,
    \ces_6_1_io_outs_up[25] ,
    \ces_6_1_io_outs_up[24] ,
    \ces_6_1_io_outs_up[23] ,
    \ces_6_1_io_outs_up[22] ,
    \ces_6_1_io_outs_up[21] ,
    \ces_6_1_io_outs_up[20] ,
    \ces_6_1_io_outs_up[19] ,
    \ces_6_1_io_outs_up[18] ,
    \ces_6_1_io_outs_up[17] ,
    \ces_6_1_io_outs_up[16] ,
    \ces_6_1_io_outs_up[15] ,
    \ces_6_1_io_outs_up[14] ,
    \ces_6_1_io_outs_up[13] ,
    \ces_6_1_io_outs_up[12] ,
    \ces_6_1_io_outs_up[11] ,
    \ces_6_1_io_outs_up[10] ,
    \ces_6_1_io_outs_up[9] ,
    \ces_6_1_io_outs_up[8] ,
    \ces_6_1_io_outs_up[7] ,
    \ces_6_1_io_outs_up[6] ,
    \ces_6_1_io_outs_up[5] ,
    \ces_6_1_io_outs_up[4] ,
    \ces_6_1_io_outs_up[3] ,
    \ces_6_1_io_outs_up[2] ,
    \ces_6_1_io_outs_up[1] ,
    \ces_6_1_io_outs_up[0] }),
    .io_outs_down({\ces_6_1_io_ins_down[63] ,
    \ces_6_1_io_ins_down[62] ,
    \ces_6_1_io_ins_down[61] ,
    \ces_6_1_io_ins_down[60] ,
    \ces_6_1_io_ins_down[59] ,
    \ces_6_1_io_ins_down[58] ,
    \ces_6_1_io_ins_down[57] ,
    \ces_6_1_io_ins_down[56] ,
    \ces_6_1_io_ins_down[55] ,
    \ces_6_1_io_ins_down[54] ,
    \ces_6_1_io_ins_down[53] ,
    \ces_6_1_io_ins_down[52] ,
    \ces_6_1_io_ins_down[51] ,
    \ces_6_1_io_ins_down[50] ,
    \ces_6_1_io_ins_down[49] ,
    \ces_6_1_io_ins_down[48] ,
    \ces_6_1_io_ins_down[47] ,
    \ces_6_1_io_ins_down[46] ,
    \ces_6_1_io_ins_down[45] ,
    \ces_6_1_io_ins_down[44] ,
    \ces_6_1_io_ins_down[43] ,
    \ces_6_1_io_ins_down[42] ,
    \ces_6_1_io_ins_down[41] ,
    \ces_6_1_io_ins_down[40] ,
    \ces_6_1_io_ins_down[39] ,
    \ces_6_1_io_ins_down[38] ,
    \ces_6_1_io_ins_down[37] ,
    \ces_6_1_io_ins_down[36] ,
    \ces_6_1_io_ins_down[35] ,
    \ces_6_1_io_ins_down[34] ,
    \ces_6_1_io_ins_down[33] ,
    \ces_6_1_io_ins_down[32] ,
    \ces_6_1_io_ins_down[31] ,
    \ces_6_1_io_ins_down[30] ,
    \ces_6_1_io_ins_down[29] ,
    \ces_6_1_io_ins_down[28] ,
    \ces_6_1_io_ins_down[27] ,
    \ces_6_1_io_ins_down[26] ,
    \ces_6_1_io_ins_down[25] ,
    \ces_6_1_io_ins_down[24] ,
    \ces_6_1_io_ins_down[23] ,
    \ces_6_1_io_ins_down[22] ,
    \ces_6_1_io_ins_down[21] ,
    \ces_6_1_io_ins_down[20] ,
    \ces_6_1_io_ins_down[19] ,
    \ces_6_1_io_ins_down[18] ,
    \ces_6_1_io_ins_down[17] ,
    \ces_6_1_io_ins_down[16] ,
    \ces_6_1_io_ins_down[15] ,
    \ces_6_1_io_ins_down[14] ,
    \ces_6_1_io_ins_down[13] ,
    \ces_6_1_io_ins_down[12] ,
    \ces_6_1_io_ins_down[11] ,
    \ces_6_1_io_ins_down[10] ,
    \ces_6_1_io_ins_down[9] ,
    \ces_6_1_io_ins_down[8] ,
    \ces_6_1_io_ins_down[7] ,
    \ces_6_1_io_ins_down[6] ,
    \ces_6_1_io_ins_down[5] ,
    \ces_6_1_io_ins_down[4] ,
    \ces_6_1_io_ins_down[3] ,
    \ces_6_1_io_ins_down[2] ,
    \ces_6_1_io_ins_down[1] ,
    \ces_6_1_io_ins_down[0] }),
    .io_outs_left({\ces_7_0_io_ins_left[63] ,
    \ces_7_0_io_ins_left[62] ,
    \ces_7_0_io_ins_left[61] ,
    \ces_7_0_io_ins_left[60] ,
    \ces_7_0_io_ins_left[59] ,
    \ces_7_0_io_ins_left[58] ,
    \ces_7_0_io_ins_left[57] ,
    \ces_7_0_io_ins_left[56] ,
    \ces_7_0_io_ins_left[55] ,
    \ces_7_0_io_ins_left[54] ,
    \ces_7_0_io_ins_left[53] ,
    \ces_7_0_io_ins_left[52] ,
    \ces_7_0_io_ins_left[51] ,
    \ces_7_0_io_ins_left[50] ,
    \ces_7_0_io_ins_left[49] ,
    \ces_7_0_io_ins_left[48] ,
    \ces_7_0_io_ins_left[47] ,
    \ces_7_0_io_ins_left[46] ,
    \ces_7_0_io_ins_left[45] ,
    \ces_7_0_io_ins_left[44] ,
    \ces_7_0_io_ins_left[43] ,
    \ces_7_0_io_ins_left[42] ,
    \ces_7_0_io_ins_left[41] ,
    \ces_7_0_io_ins_left[40] ,
    \ces_7_0_io_ins_left[39] ,
    \ces_7_0_io_ins_left[38] ,
    \ces_7_0_io_ins_left[37] ,
    \ces_7_0_io_ins_left[36] ,
    \ces_7_0_io_ins_left[35] ,
    \ces_7_0_io_ins_left[34] ,
    \ces_7_0_io_ins_left[33] ,
    \ces_7_0_io_ins_left[32] ,
    \ces_7_0_io_ins_left[31] ,
    \ces_7_0_io_ins_left[30] ,
    \ces_7_0_io_ins_left[29] ,
    \ces_7_0_io_ins_left[28] ,
    \ces_7_0_io_ins_left[27] ,
    \ces_7_0_io_ins_left[26] ,
    \ces_7_0_io_ins_left[25] ,
    \ces_7_0_io_ins_left[24] ,
    \ces_7_0_io_ins_left[23] ,
    \ces_7_0_io_ins_left[22] ,
    \ces_7_0_io_ins_left[21] ,
    \ces_7_0_io_ins_left[20] ,
    \ces_7_0_io_ins_left[19] ,
    \ces_7_0_io_ins_left[18] ,
    \ces_7_0_io_ins_left[17] ,
    \ces_7_0_io_ins_left[16] ,
    \ces_7_0_io_ins_left[15] ,
    \ces_7_0_io_ins_left[14] ,
    \ces_7_0_io_ins_left[13] ,
    \ces_7_0_io_ins_left[12] ,
    \ces_7_0_io_ins_left[11] ,
    \ces_7_0_io_ins_left[10] ,
    \ces_7_0_io_ins_left[9] ,
    \ces_7_0_io_ins_left[8] ,
    \ces_7_0_io_ins_left[7] ,
    \ces_7_0_io_ins_left[6] ,
    \ces_7_0_io_ins_left[5] ,
    \ces_7_0_io_ins_left[4] ,
    \ces_7_0_io_ins_left[3] ,
    \ces_7_0_io_ins_left[2] ,
    \ces_7_0_io_ins_left[1] ,
    \ces_7_0_io_ins_left[0] }),
    .io_outs_right({\ces_7_1_io_outs_right[63] ,
    \ces_7_1_io_outs_right[62] ,
    \ces_7_1_io_outs_right[61] ,
    \ces_7_1_io_outs_right[60] ,
    \ces_7_1_io_outs_right[59] ,
    \ces_7_1_io_outs_right[58] ,
    \ces_7_1_io_outs_right[57] ,
    \ces_7_1_io_outs_right[56] ,
    \ces_7_1_io_outs_right[55] ,
    \ces_7_1_io_outs_right[54] ,
    \ces_7_1_io_outs_right[53] ,
    \ces_7_1_io_outs_right[52] ,
    \ces_7_1_io_outs_right[51] ,
    \ces_7_1_io_outs_right[50] ,
    \ces_7_1_io_outs_right[49] ,
    \ces_7_1_io_outs_right[48] ,
    \ces_7_1_io_outs_right[47] ,
    \ces_7_1_io_outs_right[46] ,
    \ces_7_1_io_outs_right[45] ,
    \ces_7_1_io_outs_right[44] ,
    \ces_7_1_io_outs_right[43] ,
    \ces_7_1_io_outs_right[42] ,
    \ces_7_1_io_outs_right[41] ,
    \ces_7_1_io_outs_right[40] ,
    \ces_7_1_io_outs_right[39] ,
    \ces_7_1_io_outs_right[38] ,
    \ces_7_1_io_outs_right[37] ,
    \ces_7_1_io_outs_right[36] ,
    \ces_7_1_io_outs_right[35] ,
    \ces_7_1_io_outs_right[34] ,
    \ces_7_1_io_outs_right[33] ,
    \ces_7_1_io_outs_right[32] ,
    \ces_7_1_io_outs_right[31] ,
    \ces_7_1_io_outs_right[30] ,
    \ces_7_1_io_outs_right[29] ,
    \ces_7_1_io_outs_right[28] ,
    \ces_7_1_io_outs_right[27] ,
    \ces_7_1_io_outs_right[26] ,
    \ces_7_1_io_outs_right[25] ,
    \ces_7_1_io_outs_right[24] ,
    \ces_7_1_io_outs_right[23] ,
    \ces_7_1_io_outs_right[22] ,
    \ces_7_1_io_outs_right[21] ,
    \ces_7_1_io_outs_right[20] ,
    \ces_7_1_io_outs_right[19] ,
    \ces_7_1_io_outs_right[18] ,
    \ces_7_1_io_outs_right[17] ,
    \ces_7_1_io_outs_right[16] ,
    \ces_7_1_io_outs_right[15] ,
    \ces_7_1_io_outs_right[14] ,
    \ces_7_1_io_outs_right[13] ,
    \ces_7_1_io_outs_right[12] ,
    \ces_7_1_io_outs_right[11] ,
    \ces_7_1_io_outs_right[10] ,
    \ces_7_1_io_outs_right[9] ,
    \ces_7_1_io_outs_right[8] ,
    \ces_7_1_io_outs_right[7] ,
    \ces_7_1_io_outs_right[6] ,
    \ces_7_1_io_outs_right[5] ,
    \ces_7_1_io_outs_right[4] ,
    \ces_7_1_io_outs_right[3] ,
    \ces_7_1_io_outs_right[2] ,
    \ces_7_1_io_outs_right[1] ,
    \ces_7_1_io_outs_right[0] }),
    .io_outs_up({net3772,
    net3771,
    net3770,
    net3769,
    net3767,
    net3766,
    net3765,
    net3764,
    net3763,
    net3762,
    net3761,
    net3760,
    net3759,
    net3758,
    net3756,
    net3755,
    net3754,
    net3753,
    net3752,
    net3751,
    net3750,
    net3749,
    net3748,
    net3747,
    net3745,
    net3744,
    net3743,
    net3742,
    net3741,
    net3740,
    net3739,
    net3738,
    net3737,
    net3736,
    net3734,
    net3733,
    net3732,
    net3731,
    net3730,
    net3729,
    net3728,
    net3727,
    net3726,
    net3725,
    net3723,
    net3722,
    net3721,
    net3720,
    net3719,
    net3718,
    net3717,
    net3716,
    net3715,
    net3714,
    net3776,
    net3775,
    net3774,
    net3773,
    net3768,
    net3757,
    net3746,
    net3735,
    net3724,
    net3713}));
 Element ces_7_2 (.clock(clknet_3_5_0_clock),
    .io_lsbIns_1(ces_7_1_io_lsbOuts_1),
    .io_lsbIns_2(ces_7_1_io_lsbOuts_2),
    .io_lsbIns_3(ces_7_1_io_lsbOuts_3),
    .io_lsbIns_4(ces_7_1_io_lsbOuts_4),
    .io_lsbIns_5(ces_7_1_io_lsbOuts_5),
    .io_lsbIns_6(ces_7_1_io_lsbOuts_6),
    .io_lsbIns_7(ces_7_1_io_lsbOuts_7),
    .io_lsbOuts_0(ces_7_2_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_2_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_2_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_2_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_2_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_2_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_2_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_2_io_lsbOuts_7),
    .io_ins_down({net188,
    net187,
    net186,
    net185,
    net183,
    net182,
    net181,
    net180,
    net179,
    net178,
    net177,
    net176,
    net175,
    net174,
    net172,
    net171,
    net170,
    net169,
    net168,
    net167,
    net166,
    net165,
    net164,
    net163,
    net161,
    net160,
    net159,
    net158,
    net157,
    net156,
    net155,
    net154,
    net153,
    net152,
    net150,
    net149,
    net148,
    net147,
    net146,
    net145,
    net144,
    net143,
    net142,
    net141,
    net139,
    net138,
    net137,
    net136,
    net135,
    net134,
    net133,
    net132,
    net131,
    net130,
    net192,
    net191,
    net190,
    net189,
    net184,
    net173,
    net162,
    net151,
    net140,
    net129}),
    .io_ins_left({\ces_7_2_io_ins_left[63] ,
    \ces_7_2_io_ins_left[62] ,
    \ces_7_2_io_ins_left[61] ,
    \ces_7_2_io_ins_left[60] ,
    \ces_7_2_io_ins_left[59] ,
    \ces_7_2_io_ins_left[58] ,
    \ces_7_2_io_ins_left[57] ,
    \ces_7_2_io_ins_left[56] ,
    \ces_7_2_io_ins_left[55] ,
    \ces_7_2_io_ins_left[54] ,
    \ces_7_2_io_ins_left[53] ,
    \ces_7_2_io_ins_left[52] ,
    \ces_7_2_io_ins_left[51] ,
    \ces_7_2_io_ins_left[50] ,
    \ces_7_2_io_ins_left[49] ,
    \ces_7_2_io_ins_left[48] ,
    \ces_7_2_io_ins_left[47] ,
    \ces_7_2_io_ins_left[46] ,
    \ces_7_2_io_ins_left[45] ,
    \ces_7_2_io_ins_left[44] ,
    \ces_7_2_io_ins_left[43] ,
    \ces_7_2_io_ins_left[42] ,
    \ces_7_2_io_ins_left[41] ,
    \ces_7_2_io_ins_left[40] ,
    \ces_7_2_io_ins_left[39] ,
    \ces_7_2_io_ins_left[38] ,
    \ces_7_2_io_ins_left[37] ,
    \ces_7_2_io_ins_left[36] ,
    \ces_7_2_io_ins_left[35] ,
    \ces_7_2_io_ins_left[34] ,
    \ces_7_2_io_ins_left[33] ,
    \ces_7_2_io_ins_left[32] ,
    \ces_7_2_io_ins_left[31] ,
    \ces_7_2_io_ins_left[30] ,
    \ces_7_2_io_ins_left[29] ,
    \ces_7_2_io_ins_left[28] ,
    \ces_7_2_io_ins_left[27] ,
    \ces_7_2_io_ins_left[26] ,
    \ces_7_2_io_ins_left[25] ,
    \ces_7_2_io_ins_left[24] ,
    \ces_7_2_io_ins_left[23] ,
    \ces_7_2_io_ins_left[22] ,
    \ces_7_2_io_ins_left[21] ,
    \ces_7_2_io_ins_left[20] ,
    \ces_7_2_io_ins_left[19] ,
    \ces_7_2_io_ins_left[18] ,
    \ces_7_2_io_ins_left[17] ,
    \ces_7_2_io_ins_left[16] ,
    \ces_7_2_io_ins_left[15] ,
    \ces_7_2_io_ins_left[14] ,
    \ces_7_2_io_ins_left[13] ,
    \ces_7_2_io_ins_left[12] ,
    \ces_7_2_io_ins_left[11] ,
    \ces_7_2_io_ins_left[10] ,
    \ces_7_2_io_ins_left[9] ,
    \ces_7_2_io_ins_left[8] ,
    \ces_7_2_io_ins_left[7] ,
    \ces_7_2_io_ins_left[6] ,
    \ces_7_2_io_ins_left[5] ,
    \ces_7_2_io_ins_left[4] ,
    \ces_7_2_io_ins_left[3] ,
    \ces_7_2_io_ins_left[2] ,
    \ces_7_2_io_ins_left[1] ,
    \ces_7_2_io_ins_left[0] }),
    .io_ins_right({\ces_7_1_io_outs_right[63] ,
    \ces_7_1_io_outs_right[62] ,
    \ces_7_1_io_outs_right[61] ,
    \ces_7_1_io_outs_right[60] ,
    \ces_7_1_io_outs_right[59] ,
    \ces_7_1_io_outs_right[58] ,
    \ces_7_1_io_outs_right[57] ,
    \ces_7_1_io_outs_right[56] ,
    \ces_7_1_io_outs_right[55] ,
    \ces_7_1_io_outs_right[54] ,
    \ces_7_1_io_outs_right[53] ,
    \ces_7_1_io_outs_right[52] ,
    \ces_7_1_io_outs_right[51] ,
    \ces_7_1_io_outs_right[50] ,
    \ces_7_1_io_outs_right[49] ,
    \ces_7_1_io_outs_right[48] ,
    \ces_7_1_io_outs_right[47] ,
    \ces_7_1_io_outs_right[46] ,
    \ces_7_1_io_outs_right[45] ,
    \ces_7_1_io_outs_right[44] ,
    \ces_7_1_io_outs_right[43] ,
    \ces_7_1_io_outs_right[42] ,
    \ces_7_1_io_outs_right[41] ,
    \ces_7_1_io_outs_right[40] ,
    \ces_7_1_io_outs_right[39] ,
    \ces_7_1_io_outs_right[38] ,
    \ces_7_1_io_outs_right[37] ,
    \ces_7_1_io_outs_right[36] ,
    \ces_7_1_io_outs_right[35] ,
    \ces_7_1_io_outs_right[34] ,
    \ces_7_1_io_outs_right[33] ,
    \ces_7_1_io_outs_right[32] ,
    \ces_7_1_io_outs_right[31] ,
    \ces_7_1_io_outs_right[30] ,
    \ces_7_1_io_outs_right[29] ,
    \ces_7_1_io_outs_right[28] ,
    \ces_7_1_io_outs_right[27] ,
    \ces_7_1_io_outs_right[26] ,
    \ces_7_1_io_outs_right[25] ,
    \ces_7_1_io_outs_right[24] ,
    \ces_7_1_io_outs_right[23] ,
    \ces_7_1_io_outs_right[22] ,
    \ces_7_1_io_outs_right[21] ,
    \ces_7_1_io_outs_right[20] ,
    \ces_7_1_io_outs_right[19] ,
    \ces_7_1_io_outs_right[18] ,
    \ces_7_1_io_outs_right[17] ,
    \ces_7_1_io_outs_right[16] ,
    \ces_7_1_io_outs_right[15] ,
    \ces_7_1_io_outs_right[14] ,
    \ces_7_1_io_outs_right[13] ,
    \ces_7_1_io_outs_right[12] ,
    \ces_7_1_io_outs_right[11] ,
    \ces_7_1_io_outs_right[10] ,
    \ces_7_1_io_outs_right[9] ,
    \ces_7_1_io_outs_right[8] ,
    \ces_7_1_io_outs_right[7] ,
    \ces_7_1_io_outs_right[6] ,
    \ces_7_1_io_outs_right[5] ,
    \ces_7_1_io_outs_right[4] ,
    \ces_7_1_io_outs_right[3] ,
    \ces_7_1_io_outs_right[2] ,
    \ces_7_1_io_outs_right[1] ,
    \ces_7_1_io_outs_right[0] }),
    .io_ins_up({\ces_6_2_io_outs_up[63] ,
    \ces_6_2_io_outs_up[62] ,
    \ces_6_2_io_outs_up[61] ,
    \ces_6_2_io_outs_up[60] ,
    \ces_6_2_io_outs_up[59] ,
    \ces_6_2_io_outs_up[58] ,
    \ces_6_2_io_outs_up[57] ,
    \ces_6_2_io_outs_up[56] ,
    \ces_6_2_io_outs_up[55] ,
    \ces_6_2_io_outs_up[54] ,
    \ces_6_2_io_outs_up[53] ,
    \ces_6_2_io_outs_up[52] ,
    \ces_6_2_io_outs_up[51] ,
    \ces_6_2_io_outs_up[50] ,
    \ces_6_2_io_outs_up[49] ,
    \ces_6_2_io_outs_up[48] ,
    \ces_6_2_io_outs_up[47] ,
    \ces_6_2_io_outs_up[46] ,
    \ces_6_2_io_outs_up[45] ,
    \ces_6_2_io_outs_up[44] ,
    \ces_6_2_io_outs_up[43] ,
    \ces_6_2_io_outs_up[42] ,
    \ces_6_2_io_outs_up[41] ,
    \ces_6_2_io_outs_up[40] ,
    \ces_6_2_io_outs_up[39] ,
    \ces_6_2_io_outs_up[38] ,
    \ces_6_2_io_outs_up[37] ,
    \ces_6_2_io_outs_up[36] ,
    \ces_6_2_io_outs_up[35] ,
    \ces_6_2_io_outs_up[34] ,
    \ces_6_2_io_outs_up[33] ,
    \ces_6_2_io_outs_up[32] ,
    \ces_6_2_io_outs_up[31] ,
    \ces_6_2_io_outs_up[30] ,
    \ces_6_2_io_outs_up[29] ,
    \ces_6_2_io_outs_up[28] ,
    \ces_6_2_io_outs_up[27] ,
    \ces_6_2_io_outs_up[26] ,
    \ces_6_2_io_outs_up[25] ,
    \ces_6_2_io_outs_up[24] ,
    \ces_6_2_io_outs_up[23] ,
    \ces_6_2_io_outs_up[22] ,
    \ces_6_2_io_outs_up[21] ,
    \ces_6_2_io_outs_up[20] ,
    \ces_6_2_io_outs_up[19] ,
    \ces_6_2_io_outs_up[18] ,
    \ces_6_2_io_outs_up[17] ,
    \ces_6_2_io_outs_up[16] ,
    \ces_6_2_io_outs_up[15] ,
    \ces_6_2_io_outs_up[14] ,
    \ces_6_2_io_outs_up[13] ,
    \ces_6_2_io_outs_up[12] ,
    \ces_6_2_io_outs_up[11] ,
    \ces_6_2_io_outs_up[10] ,
    \ces_6_2_io_outs_up[9] ,
    \ces_6_2_io_outs_up[8] ,
    \ces_6_2_io_outs_up[7] ,
    \ces_6_2_io_outs_up[6] ,
    \ces_6_2_io_outs_up[5] ,
    \ces_6_2_io_outs_up[4] ,
    \ces_6_2_io_outs_up[3] ,
    \ces_6_2_io_outs_up[2] ,
    \ces_6_2_io_outs_up[1] ,
    \ces_6_2_io_outs_up[0] }),
    .io_outs_down({\ces_6_2_io_ins_down[63] ,
    \ces_6_2_io_ins_down[62] ,
    \ces_6_2_io_ins_down[61] ,
    \ces_6_2_io_ins_down[60] ,
    \ces_6_2_io_ins_down[59] ,
    \ces_6_2_io_ins_down[58] ,
    \ces_6_2_io_ins_down[57] ,
    \ces_6_2_io_ins_down[56] ,
    \ces_6_2_io_ins_down[55] ,
    \ces_6_2_io_ins_down[54] ,
    \ces_6_2_io_ins_down[53] ,
    \ces_6_2_io_ins_down[52] ,
    \ces_6_2_io_ins_down[51] ,
    \ces_6_2_io_ins_down[50] ,
    \ces_6_2_io_ins_down[49] ,
    \ces_6_2_io_ins_down[48] ,
    \ces_6_2_io_ins_down[47] ,
    \ces_6_2_io_ins_down[46] ,
    \ces_6_2_io_ins_down[45] ,
    \ces_6_2_io_ins_down[44] ,
    \ces_6_2_io_ins_down[43] ,
    \ces_6_2_io_ins_down[42] ,
    \ces_6_2_io_ins_down[41] ,
    \ces_6_2_io_ins_down[40] ,
    \ces_6_2_io_ins_down[39] ,
    \ces_6_2_io_ins_down[38] ,
    \ces_6_2_io_ins_down[37] ,
    \ces_6_2_io_ins_down[36] ,
    \ces_6_2_io_ins_down[35] ,
    \ces_6_2_io_ins_down[34] ,
    \ces_6_2_io_ins_down[33] ,
    \ces_6_2_io_ins_down[32] ,
    \ces_6_2_io_ins_down[31] ,
    \ces_6_2_io_ins_down[30] ,
    \ces_6_2_io_ins_down[29] ,
    \ces_6_2_io_ins_down[28] ,
    \ces_6_2_io_ins_down[27] ,
    \ces_6_2_io_ins_down[26] ,
    \ces_6_2_io_ins_down[25] ,
    \ces_6_2_io_ins_down[24] ,
    \ces_6_2_io_ins_down[23] ,
    \ces_6_2_io_ins_down[22] ,
    \ces_6_2_io_ins_down[21] ,
    \ces_6_2_io_ins_down[20] ,
    \ces_6_2_io_ins_down[19] ,
    \ces_6_2_io_ins_down[18] ,
    \ces_6_2_io_ins_down[17] ,
    \ces_6_2_io_ins_down[16] ,
    \ces_6_2_io_ins_down[15] ,
    \ces_6_2_io_ins_down[14] ,
    \ces_6_2_io_ins_down[13] ,
    \ces_6_2_io_ins_down[12] ,
    \ces_6_2_io_ins_down[11] ,
    \ces_6_2_io_ins_down[10] ,
    \ces_6_2_io_ins_down[9] ,
    \ces_6_2_io_ins_down[8] ,
    \ces_6_2_io_ins_down[7] ,
    \ces_6_2_io_ins_down[6] ,
    \ces_6_2_io_ins_down[5] ,
    \ces_6_2_io_ins_down[4] ,
    \ces_6_2_io_ins_down[3] ,
    \ces_6_2_io_ins_down[2] ,
    \ces_6_2_io_ins_down[1] ,
    \ces_6_2_io_ins_down[0] }),
    .io_outs_left({\ces_7_1_io_ins_left[63] ,
    \ces_7_1_io_ins_left[62] ,
    \ces_7_1_io_ins_left[61] ,
    \ces_7_1_io_ins_left[60] ,
    \ces_7_1_io_ins_left[59] ,
    \ces_7_1_io_ins_left[58] ,
    \ces_7_1_io_ins_left[57] ,
    \ces_7_1_io_ins_left[56] ,
    \ces_7_1_io_ins_left[55] ,
    \ces_7_1_io_ins_left[54] ,
    \ces_7_1_io_ins_left[53] ,
    \ces_7_1_io_ins_left[52] ,
    \ces_7_1_io_ins_left[51] ,
    \ces_7_1_io_ins_left[50] ,
    \ces_7_1_io_ins_left[49] ,
    \ces_7_1_io_ins_left[48] ,
    \ces_7_1_io_ins_left[47] ,
    \ces_7_1_io_ins_left[46] ,
    \ces_7_1_io_ins_left[45] ,
    \ces_7_1_io_ins_left[44] ,
    \ces_7_1_io_ins_left[43] ,
    \ces_7_1_io_ins_left[42] ,
    \ces_7_1_io_ins_left[41] ,
    \ces_7_1_io_ins_left[40] ,
    \ces_7_1_io_ins_left[39] ,
    \ces_7_1_io_ins_left[38] ,
    \ces_7_1_io_ins_left[37] ,
    \ces_7_1_io_ins_left[36] ,
    \ces_7_1_io_ins_left[35] ,
    \ces_7_1_io_ins_left[34] ,
    \ces_7_1_io_ins_left[33] ,
    \ces_7_1_io_ins_left[32] ,
    \ces_7_1_io_ins_left[31] ,
    \ces_7_1_io_ins_left[30] ,
    \ces_7_1_io_ins_left[29] ,
    \ces_7_1_io_ins_left[28] ,
    \ces_7_1_io_ins_left[27] ,
    \ces_7_1_io_ins_left[26] ,
    \ces_7_1_io_ins_left[25] ,
    \ces_7_1_io_ins_left[24] ,
    \ces_7_1_io_ins_left[23] ,
    \ces_7_1_io_ins_left[22] ,
    \ces_7_1_io_ins_left[21] ,
    \ces_7_1_io_ins_left[20] ,
    \ces_7_1_io_ins_left[19] ,
    \ces_7_1_io_ins_left[18] ,
    \ces_7_1_io_ins_left[17] ,
    \ces_7_1_io_ins_left[16] ,
    \ces_7_1_io_ins_left[15] ,
    \ces_7_1_io_ins_left[14] ,
    \ces_7_1_io_ins_left[13] ,
    \ces_7_1_io_ins_left[12] ,
    \ces_7_1_io_ins_left[11] ,
    \ces_7_1_io_ins_left[10] ,
    \ces_7_1_io_ins_left[9] ,
    \ces_7_1_io_ins_left[8] ,
    \ces_7_1_io_ins_left[7] ,
    \ces_7_1_io_ins_left[6] ,
    \ces_7_1_io_ins_left[5] ,
    \ces_7_1_io_ins_left[4] ,
    \ces_7_1_io_ins_left[3] ,
    \ces_7_1_io_ins_left[2] ,
    \ces_7_1_io_ins_left[1] ,
    \ces_7_1_io_ins_left[0] }),
    .io_outs_right({\ces_7_2_io_outs_right[63] ,
    \ces_7_2_io_outs_right[62] ,
    \ces_7_2_io_outs_right[61] ,
    \ces_7_2_io_outs_right[60] ,
    \ces_7_2_io_outs_right[59] ,
    \ces_7_2_io_outs_right[58] ,
    \ces_7_2_io_outs_right[57] ,
    \ces_7_2_io_outs_right[56] ,
    \ces_7_2_io_outs_right[55] ,
    \ces_7_2_io_outs_right[54] ,
    \ces_7_2_io_outs_right[53] ,
    \ces_7_2_io_outs_right[52] ,
    \ces_7_2_io_outs_right[51] ,
    \ces_7_2_io_outs_right[50] ,
    \ces_7_2_io_outs_right[49] ,
    \ces_7_2_io_outs_right[48] ,
    \ces_7_2_io_outs_right[47] ,
    \ces_7_2_io_outs_right[46] ,
    \ces_7_2_io_outs_right[45] ,
    \ces_7_2_io_outs_right[44] ,
    \ces_7_2_io_outs_right[43] ,
    \ces_7_2_io_outs_right[42] ,
    \ces_7_2_io_outs_right[41] ,
    \ces_7_2_io_outs_right[40] ,
    \ces_7_2_io_outs_right[39] ,
    \ces_7_2_io_outs_right[38] ,
    \ces_7_2_io_outs_right[37] ,
    \ces_7_2_io_outs_right[36] ,
    \ces_7_2_io_outs_right[35] ,
    \ces_7_2_io_outs_right[34] ,
    \ces_7_2_io_outs_right[33] ,
    \ces_7_2_io_outs_right[32] ,
    \ces_7_2_io_outs_right[31] ,
    \ces_7_2_io_outs_right[30] ,
    \ces_7_2_io_outs_right[29] ,
    \ces_7_2_io_outs_right[28] ,
    \ces_7_2_io_outs_right[27] ,
    \ces_7_2_io_outs_right[26] ,
    \ces_7_2_io_outs_right[25] ,
    \ces_7_2_io_outs_right[24] ,
    \ces_7_2_io_outs_right[23] ,
    \ces_7_2_io_outs_right[22] ,
    \ces_7_2_io_outs_right[21] ,
    \ces_7_2_io_outs_right[20] ,
    \ces_7_2_io_outs_right[19] ,
    \ces_7_2_io_outs_right[18] ,
    \ces_7_2_io_outs_right[17] ,
    \ces_7_2_io_outs_right[16] ,
    \ces_7_2_io_outs_right[15] ,
    \ces_7_2_io_outs_right[14] ,
    \ces_7_2_io_outs_right[13] ,
    \ces_7_2_io_outs_right[12] ,
    \ces_7_2_io_outs_right[11] ,
    \ces_7_2_io_outs_right[10] ,
    \ces_7_2_io_outs_right[9] ,
    \ces_7_2_io_outs_right[8] ,
    \ces_7_2_io_outs_right[7] ,
    \ces_7_2_io_outs_right[6] ,
    \ces_7_2_io_outs_right[5] ,
    \ces_7_2_io_outs_right[4] ,
    \ces_7_2_io_outs_right[3] ,
    \ces_7_2_io_outs_right[2] ,
    \ces_7_2_io_outs_right[1] ,
    \ces_7_2_io_outs_right[0] }),
    .io_outs_up({net3836,
    net3835,
    net3834,
    net3833,
    net3831,
    net3830,
    net3829,
    net3828,
    net3827,
    net3826,
    net3825,
    net3824,
    net3823,
    net3822,
    net3820,
    net3819,
    net3818,
    net3817,
    net3816,
    net3815,
    net3814,
    net3813,
    net3812,
    net3811,
    net3809,
    net3808,
    net3807,
    net3806,
    net3805,
    net3804,
    net3803,
    net3802,
    net3801,
    net3800,
    net3798,
    net3797,
    net3796,
    net3795,
    net3794,
    net3793,
    net3792,
    net3791,
    net3790,
    net3789,
    net3787,
    net3786,
    net3785,
    net3784,
    net3783,
    net3782,
    net3781,
    net3780,
    net3779,
    net3778,
    net3840,
    net3839,
    net3838,
    net3837,
    net3832,
    net3821,
    net3810,
    net3799,
    net3788,
    net3777}));
 Element ces_7_3 (.clock(clknet_3_5_0_clock),
    .io_lsbIns_1(ces_7_2_io_lsbOuts_1),
    .io_lsbIns_2(ces_7_2_io_lsbOuts_2),
    .io_lsbIns_3(ces_7_2_io_lsbOuts_3),
    .io_lsbIns_4(ces_7_2_io_lsbOuts_4),
    .io_lsbIns_5(ces_7_2_io_lsbOuts_5),
    .io_lsbIns_6(ces_7_2_io_lsbOuts_6),
    .io_lsbIns_7(ces_7_2_io_lsbOuts_7),
    .io_lsbOuts_0(ces_7_3_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_3_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_3_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_3_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_3_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_3_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_3_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_3_io_lsbOuts_7),
    .io_ins_down({net252,
    net251,
    net250,
    net249,
    net247,
    net246,
    net245,
    net244,
    net243,
    net242,
    net241,
    net240,
    net239,
    net238,
    net236,
    net235,
    net234,
    net233,
    net232,
    net231,
    net230,
    net229,
    net228,
    net227,
    net225,
    net224,
    net223,
    net222,
    net221,
    net220,
    net219,
    net218,
    net217,
    net216,
    net214,
    net213,
    net212,
    net211,
    net210,
    net209,
    net208,
    net207,
    net206,
    net205,
    net203,
    net202,
    net201,
    net200,
    net199,
    net198,
    net197,
    net196,
    net195,
    net194,
    net256,
    net255,
    net254,
    net253,
    net248,
    net237,
    net226,
    net215,
    net204,
    net193}),
    .io_ins_left({\ces_7_3_io_ins_left[63] ,
    \ces_7_3_io_ins_left[62] ,
    \ces_7_3_io_ins_left[61] ,
    \ces_7_3_io_ins_left[60] ,
    \ces_7_3_io_ins_left[59] ,
    \ces_7_3_io_ins_left[58] ,
    \ces_7_3_io_ins_left[57] ,
    \ces_7_3_io_ins_left[56] ,
    \ces_7_3_io_ins_left[55] ,
    \ces_7_3_io_ins_left[54] ,
    \ces_7_3_io_ins_left[53] ,
    \ces_7_3_io_ins_left[52] ,
    \ces_7_3_io_ins_left[51] ,
    \ces_7_3_io_ins_left[50] ,
    \ces_7_3_io_ins_left[49] ,
    \ces_7_3_io_ins_left[48] ,
    \ces_7_3_io_ins_left[47] ,
    \ces_7_3_io_ins_left[46] ,
    \ces_7_3_io_ins_left[45] ,
    \ces_7_3_io_ins_left[44] ,
    \ces_7_3_io_ins_left[43] ,
    \ces_7_3_io_ins_left[42] ,
    \ces_7_3_io_ins_left[41] ,
    \ces_7_3_io_ins_left[40] ,
    \ces_7_3_io_ins_left[39] ,
    \ces_7_3_io_ins_left[38] ,
    \ces_7_3_io_ins_left[37] ,
    \ces_7_3_io_ins_left[36] ,
    \ces_7_3_io_ins_left[35] ,
    \ces_7_3_io_ins_left[34] ,
    \ces_7_3_io_ins_left[33] ,
    \ces_7_3_io_ins_left[32] ,
    \ces_7_3_io_ins_left[31] ,
    \ces_7_3_io_ins_left[30] ,
    \ces_7_3_io_ins_left[29] ,
    \ces_7_3_io_ins_left[28] ,
    \ces_7_3_io_ins_left[27] ,
    \ces_7_3_io_ins_left[26] ,
    \ces_7_3_io_ins_left[25] ,
    \ces_7_3_io_ins_left[24] ,
    \ces_7_3_io_ins_left[23] ,
    \ces_7_3_io_ins_left[22] ,
    \ces_7_3_io_ins_left[21] ,
    \ces_7_3_io_ins_left[20] ,
    \ces_7_3_io_ins_left[19] ,
    \ces_7_3_io_ins_left[18] ,
    \ces_7_3_io_ins_left[17] ,
    \ces_7_3_io_ins_left[16] ,
    \ces_7_3_io_ins_left[15] ,
    \ces_7_3_io_ins_left[14] ,
    \ces_7_3_io_ins_left[13] ,
    \ces_7_3_io_ins_left[12] ,
    \ces_7_3_io_ins_left[11] ,
    \ces_7_3_io_ins_left[10] ,
    \ces_7_3_io_ins_left[9] ,
    \ces_7_3_io_ins_left[8] ,
    \ces_7_3_io_ins_left[7] ,
    \ces_7_3_io_ins_left[6] ,
    \ces_7_3_io_ins_left[5] ,
    \ces_7_3_io_ins_left[4] ,
    \ces_7_3_io_ins_left[3] ,
    \ces_7_3_io_ins_left[2] ,
    \ces_7_3_io_ins_left[1] ,
    \ces_7_3_io_ins_left[0] }),
    .io_ins_right({\ces_7_2_io_outs_right[63] ,
    \ces_7_2_io_outs_right[62] ,
    \ces_7_2_io_outs_right[61] ,
    \ces_7_2_io_outs_right[60] ,
    \ces_7_2_io_outs_right[59] ,
    \ces_7_2_io_outs_right[58] ,
    \ces_7_2_io_outs_right[57] ,
    \ces_7_2_io_outs_right[56] ,
    \ces_7_2_io_outs_right[55] ,
    \ces_7_2_io_outs_right[54] ,
    \ces_7_2_io_outs_right[53] ,
    \ces_7_2_io_outs_right[52] ,
    \ces_7_2_io_outs_right[51] ,
    \ces_7_2_io_outs_right[50] ,
    \ces_7_2_io_outs_right[49] ,
    \ces_7_2_io_outs_right[48] ,
    \ces_7_2_io_outs_right[47] ,
    \ces_7_2_io_outs_right[46] ,
    \ces_7_2_io_outs_right[45] ,
    \ces_7_2_io_outs_right[44] ,
    \ces_7_2_io_outs_right[43] ,
    \ces_7_2_io_outs_right[42] ,
    \ces_7_2_io_outs_right[41] ,
    \ces_7_2_io_outs_right[40] ,
    \ces_7_2_io_outs_right[39] ,
    \ces_7_2_io_outs_right[38] ,
    \ces_7_2_io_outs_right[37] ,
    \ces_7_2_io_outs_right[36] ,
    \ces_7_2_io_outs_right[35] ,
    \ces_7_2_io_outs_right[34] ,
    \ces_7_2_io_outs_right[33] ,
    \ces_7_2_io_outs_right[32] ,
    \ces_7_2_io_outs_right[31] ,
    \ces_7_2_io_outs_right[30] ,
    \ces_7_2_io_outs_right[29] ,
    \ces_7_2_io_outs_right[28] ,
    \ces_7_2_io_outs_right[27] ,
    \ces_7_2_io_outs_right[26] ,
    \ces_7_2_io_outs_right[25] ,
    \ces_7_2_io_outs_right[24] ,
    \ces_7_2_io_outs_right[23] ,
    \ces_7_2_io_outs_right[22] ,
    \ces_7_2_io_outs_right[21] ,
    \ces_7_2_io_outs_right[20] ,
    \ces_7_2_io_outs_right[19] ,
    \ces_7_2_io_outs_right[18] ,
    \ces_7_2_io_outs_right[17] ,
    \ces_7_2_io_outs_right[16] ,
    \ces_7_2_io_outs_right[15] ,
    \ces_7_2_io_outs_right[14] ,
    \ces_7_2_io_outs_right[13] ,
    \ces_7_2_io_outs_right[12] ,
    \ces_7_2_io_outs_right[11] ,
    \ces_7_2_io_outs_right[10] ,
    \ces_7_2_io_outs_right[9] ,
    \ces_7_2_io_outs_right[8] ,
    \ces_7_2_io_outs_right[7] ,
    \ces_7_2_io_outs_right[6] ,
    \ces_7_2_io_outs_right[5] ,
    \ces_7_2_io_outs_right[4] ,
    \ces_7_2_io_outs_right[3] ,
    \ces_7_2_io_outs_right[2] ,
    \ces_7_2_io_outs_right[1] ,
    \ces_7_2_io_outs_right[0] }),
    .io_ins_up({\ces_6_3_io_outs_up[63] ,
    \ces_6_3_io_outs_up[62] ,
    \ces_6_3_io_outs_up[61] ,
    \ces_6_3_io_outs_up[60] ,
    \ces_6_3_io_outs_up[59] ,
    \ces_6_3_io_outs_up[58] ,
    \ces_6_3_io_outs_up[57] ,
    \ces_6_3_io_outs_up[56] ,
    \ces_6_3_io_outs_up[55] ,
    \ces_6_3_io_outs_up[54] ,
    \ces_6_3_io_outs_up[53] ,
    \ces_6_3_io_outs_up[52] ,
    \ces_6_3_io_outs_up[51] ,
    \ces_6_3_io_outs_up[50] ,
    \ces_6_3_io_outs_up[49] ,
    \ces_6_3_io_outs_up[48] ,
    \ces_6_3_io_outs_up[47] ,
    \ces_6_3_io_outs_up[46] ,
    \ces_6_3_io_outs_up[45] ,
    \ces_6_3_io_outs_up[44] ,
    \ces_6_3_io_outs_up[43] ,
    \ces_6_3_io_outs_up[42] ,
    \ces_6_3_io_outs_up[41] ,
    \ces_6_3_io_outs_up[40] ,
    \ces_6_3_io_outs_up[39] ,
    \ces_6_3_io_outs_up[38] ,
    \ces_6_3_io_outs_up[37] ,
    \ces_6_3_io_outs_up[36] ,
    \ces_6_3_io_outs_up[35] ,
    \ces_6_3_io_outs_up[34] ,
    \ces_6_3_io_outs_up[33] ,
    \ces_6_3_io_outs_up[32] ,
    \ces_6_3_io_outs_up[31] ,
    \ces_6_3_io_outs_up[30] ,
    \ces_6_3_io_outs_up[29] ,
    \ces_6_3_io_outs_up[28] ,
    \ces_6_3_io_outs_up[27] ,
    \ces_6_3_io_outs_up[26] ,
    \ces_6_3_io_outs_up[25] ,
    \ces_6_3_io_outs_up[24] ,
    \ces_6_3_io_outs_up[23] ,
    \ces_6_3_io_outs_up[22] ,
    \ces_6_3_io_outs_up[21] ,
    \ces_6_3_io_outs_up[20] ,
    \ces_6_3_io_outs_up[19] ,
    \ces_6_3_io_outs_up[18] ,
    \ces_6_3_io_outs_up[17] ,
    \ces_6_3_io_outs_up[16] ,
    \ces_6_3_io_outs_up[15] ,
    \ces_6_3_io_outs_up[14] ,
    \ces_6_3_io_outs_up[13] ,
    \ces_6_3_io_outs_up[12] ,
    \ces_6_3_io_outs_up[11] ,
    \ces_6_3_io_outs_up[10] ,
    \ces_6_3_io_outs_up[9] ,
    \ces_6_3_io_outs_up[8] ,
    \ces_6_3_io_outs_up[7] ,
    \ces_6_3_io_outs_up[6] ,
    \ces_6_3_io_outs_up[5] ,
    \ces_6_3_io_outs_up[4] ,
    \ces_6_3_io_outs_up[3] ,
    \ces_6_3_io_outs_up[2] ,
    \ces_6_3_io_outs_up[1] ,
    \ces_6_3_io_outs_up[0] }),
    .io_outs_down({\ces_6_3_io_ins_down[63] ,
    \ces_6_3_io_ins_down[62] ,
    \ces_6_3_io_ins_down[61] ,
    \ces_6_3_io_ins_down[60] ,
    \ces_6_3_io_ins_down[59] ,
    \ces_6_3_io_ins_down[58] ,
    \ces_6_3_io_ins_down[57] ,
    \ces_6_3_io_ins_down[56] ,
    \ces_6_3_io_ins_down[55] ,
    \ces_6_3_io_ins_down[54] ,
    \ces_6_3_io_ins_down[53] ,
    \ces_6_3_io_ins_down[52] ,
    \ces_6_3_io_ins_down[51] ,
    \ces_6_3_io_ins_down[50] ,
    \ces_6_3_io_ins_down[49] ,
    \ces_6_3_io_ins_down[48] ,
    \ces_6_3_io_ins_down[47] ,
    \ces_6_3_io_ins_down[46] ,
    \ces_6_3_io_ins_down[45] ,
    \ces_6_3_io_ins_down[44] ,
    \ces_6_3_io_ins_down[43] ,
    \ces_6_3_io_ins_down[42] ,
    \ces_6_3_io_ins_down[41] ,
    \ces_6_3_io_ins_down[40] ,
    \ces_6_3_io_ins_down[39] ,
    \ces_6_3_io_ins_down[38] ,
    \ces_6_3_io_ins_down[37] ,
    \ces_6_3_io_ins_down[36] ,
    \ces_6_3_io_ins_down[35] ,
    \ces_6_3_io_ins_down[34] ,
    \ces_6_3_io_ins_down[33] ,
    \ces_6_3_io_ins_down[32] ,
    \ces_6_3_io_ins_down[31] ,
    \ces_6_3_io_ins_down[30] ,
    \ces_6_3_io_ins_down[29] ,
    \ces_6_3_io_ins_down[28] ,
    \ces_6_3_io_ins_down[27] ,
    \ces_6_3_io_ins_down[26] ,
    \ces_6_3_io_ins_down[25] ,
    \ces_6_3_io_ins_down[24] ,
    \ces_6_3_io_ins_down[23] ,
    \ces_6_3_io_ins_down[22] ,
    \ces_6_3_io_ins_down[21] ,
    \ces_6_3_io_ins_down[20] ,
    \ces_6_3_io_ins_down[19] ,
    \ces_6_3_io_ins_down[18] ,
    \ces_6_3_io_ins_down[17] ,
    \ces_6_3_io_ins_down[16] ,
    \ces_6_3_io_ins_down[15] ,
    \ces_6_3_io_ins_down[14] ,
    \ces_6_3_io_ins_down[13] ,
    \ces_6_3_io_ins_down[12] ,
    \ces_6_3_io_ins_down[11] ,
    \ces_6_3_io_ins_down[10] ,
    \ces_6_3_io_ins_down[9] ,
    \ces_6_3_io_ins_down[8] ,
    \ces_6_3_io_ins_down[7] ,
    \ces_6_3_io_ins_down[6] ,
    \ces_6_3_io_ins_down[5] ,
    \ces_6_3_io_ins_down[4] ,
    \ces_6_3_io_ins_down[3] ,
    \ces_6_3_io_ins_down[2] ,
    \ces_6_3_io_ins_down[1] ,
    \ces_6_3_io_ins_down[0] }),
    .io_outs_left({\ces_7_2_io_ins_left[63] ,
    \ces_7_2_io_ins_left[62] ,
    \ces_7_2_io_ins_left[61] ,
    \ces_7_2_io_ins_left[60] ,
    \ces_7_2_io_ins_left[59] ,
    \ces_7_2_io_ins_left[58] ,
    \ces_7_2_io_ins_left[57] ,
    \ces_7_2_io_ins_left[56] ,
    \ces_7_2_io_ins_left[55] ,
    \ces_7_2_io_ins_left[54] ,
    \ces_7_2_io_ins_left[53] ,
    \ces_7_2_io_ins_left[52] ,
    \ces_7_2_io_ins_left[51] ,
    \ces_7_2_io_ins_left[50] ,
    \ces_7_2_io_ins_left[49] ,
    \ces_7_2_io_ins_left[48] ,
    \ces_7_2_io_ins_left[47] ,
    \ces_7_2_io_ins_left[46] ,
    \ces_7_2_io_ins_left[45] ,
    \ces_7_2_io_ins_left[44] ,
    \ces_7_2_io_ins_left[43] ,
    \ces_7_2_io_ins_left[42] ,
    \ces_7_2_io_ins_left[41] ,
    \ces_7_2_io_ins_left[40] ,
    \ces_7_2_io_ins_left[39] ,
    \ces_7_2_io_ins_left[38] ,
    \ces_7_2_io_ins_left[37] ,
    \ces_7_2_io_ins_left[36] ,
    \ces_7_2_io_ins_left[35] ,
    \ces_7_2_io_ins_left[34] ,
    \ces_7_2_io_ins_left[33] ,
    \ces_7_2_io_ins_left[32] ,
    \ces_7_2_io_ins_left[31] ,
    \ces_7_2_io_ins_left[30] ,
    \ces_7_2_io_ins_left[29] ,
    \ces_7_2_io_ins_left[28] ,
    \ces_7_2_io_ins_left[27] ,
    \ces_7_2_io_ins_left[26] ,
    \ces_7_2_io_ins_left[25] ,
    \ces_7_2_io_ins_left[24] ,
    \ces_7_2_io_ins_left[23] ,
    \ces_7_2_io_ins_left[22] ,
    \ces_7_2_io_ins_left[21] ,
    \ces_7_2_io_ins_left[20] ,
    \ces_7_2_io_ins_left[19] ,
    \ces_7_2_io_ins_left[18] ,
    \ces_7_2_io_ins_left[17] ,
    \ces_7_2_io_ins_left[16] ,
    \ces_7_2_io_ins_left[15] ,
    \ces_7_2_io_ins_left[14] ,
    \ces_7_2_io_ins_left[13] ,
    \ces_7_2_io_ins_left[12] ,
    \ces_7_2_io_ins_left[11] ,
    \ces_7_2_io_ins_left[10] ,
    \ces_7_2_io_ins_left[9] ,
    \ces_7_2_io_ins_left[8] ,
    \ces_7_2_io_ins_left[7] ,
    \ces_7_2_io_ins_left[6] ,
    \ces_7_2_io_ins_left[5] ,
    \ces_7_2_io_ins_left[4] ,
    \ces_7_2_io_ins_left[3] ,
    \ces_7_2_io_ins_left[2] ,
    \ces_7_2_io_ins_left[1] ,
    \ces_7_2_io_ins_left[0] }),
    .io_outs_right({\ces_7_3_io_outs_right[63] ,
    \ces_7_3_io_outs_right[62] ,
    \ces_7_3_io_outs_right[61] ,
    \ces_7_3_io_outs_right[60] ,
    \ces_7_3_io_outs_right[59] ,
    \ces_7_3_io_outs_right[58] ,
    \ces_7_3_io_outs_right[57] ,
    \ces_7_3_io_outs_right[56] ,
    \ces_7_3_io_outs_right[55] ,
    \ces_7_3_io_outs_right[54] ,
    \ces_7_3_io_outs_right[53] ,
    \ces_7_3_io_outs_right[52] ,
    \ces_7_3_io_outs_right[51] ,
    \ces_7_3_io_outs_right[50] ,
    \ces_7_3_io_outs_right[49] ,
    \ces_7_3_io_outs_right[48] ,
    \ces_7_3_io_outs_right[47] ,
    \ces_7_3_io_outs_right[46] ,
    \ces_7_3_io_outs_right[45] ,
    \ces_7_3_io_outs_right[44] ,
    \ces_7_3_io_outs_right[43] ,
    \ces_7_3_io_outs_right[42] ,
    \ces_7_3_io_outs_right[41] ,
    \ces_7_3_io_outs_right[40] ,
    \ces_7_3_io_outs_right[39] ,
    \ces_7_3_io_outs_right[38] ,
    \ces_7_3_io_outs_right[37] ,
    \ces_7_3_io_outs_right[36] ,
    \ces_7_3_io_outs_right[35] ,
    \ces_7_3_io_outs_right[34] ,
    \ces_7_3_io_outs_right[33] ,
    \ces_7_3_io_outs_right[32] ,
    \ces_7_3_io_outs_right[31] ,
    \ces_7_3_io_outs_right[30] ,
    \ces_7_3_io_outs_right[29] ,
    \ces_7_3_io_outs_right[28] ,
    \ces_7_3_io_outs_right[27] ,
    \ces_7_3_io_outs_right[26] ,
    \ces_7_3_io_outs_right[25] ,
    \ces_7_3_io_outs_right[24] ,
    \ces_7_3_io_outs_right[23] ,
    \ces_7_3_io_outs_right[22] ,
    \ces_7_3_io_outs_right[21] ,
    \ces_7_3_io_outs_right[20] ,
    \ces_7_3_io_outs_right[19] ,
    \ces_7_3_io_outs_right[18] ,
    \ces_7_3_io_outs_right[17] ,
    \ces_7_3_io_outs_right[16] ,
    \ces_7_3_io_outs_right[15] ,
    \ces_7_3_io_outs_right[14] ,
    \ces_7_3_io_outs_right[13] ,
    \ces_7_3_io_outs_right[12] ,
    \ces_7_3_io_outs_right[11] ,
    \ces_7_3_io_outs_right[10] ,
    \ces_7_3_io_outs_right[9] ,
    \ces_7_3_io_outs_right[8] ,
    \ces_7_3_io_outs_right[7] ,
    \ces_7_3_io_outs_right[6] ,
    \ces_7_3_io_outs_right[5] ,
    \ces_7_3_io_outs_right[4] ,
    \ces_7_3_io_outs_right[3] ,
    \ces_7_3_io_outs_right[2] ,
    \ces_7_3_io_outs_right[1] ,
    \ces_7_3_io_outs_right[0] }),
    .io_outs_up({net3900,
    net3899,
    net3898,
    net3897,
    net3895,
    net3894,
    net3893,
    net3892,
    net3891,
    net3890,
    net3889,
    net3888,
    net3887,
    net3886,
    net3884,
    net3883,
    net3882,
    net3881,
    net3880,
    net3879,
    net3878,
    net3877,
    net3876,
    net3875,
    net3873,
    net3872,
    net3871,
    net3870,
    net3869,
    net3868,
    net3867,
    net3866,
    net3865,
    net3864,
    net3862,
    net3861,
    net3860,
    net3859,
    net3858,
    net3857,
    net3856,
    net3855,
    net3854,
    net3853,
    net3851,
    net3850,
    net3849,
    net3848,
    net3847,
    net3846,
    net3845,
    net3844,
    net3843,
    net3842,
    net3904,
    net3903,
    net3902,
    net3901,
    net3896,
    net3885,
    net3874,
    net3863,
    net3852,
    net3841}));
 Element ces_7_4 (.clock(clknet_3_7_0_clock),
    .io_lsbIns_1(ces_7_3_io_lsbOuts_1),
    .io_lsbIns_2(ces_7_3_io_lsbOuts_2),
    .io_lsbIns_3(ces_7_3_io_lsbOuts_3),
    .io_lsbIns_4(ces_7_3_io_lsbOuts_4),
    .io_lsbIns_5(ces_7_3_io_lsbOuts_5),
    .io_lsbIns_6(ces_7_3_io_lsbOuts_6),
    .io_lsbIns_7(ces_7_3_io_lsbOuts_7),
    .io_lsbOuts_0(ces_7_4_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_4_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_4_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_4_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_4_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_4_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_4_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_4_io_lsbOuts_7),
    .io_ins_down({net316,
    net315,
    net314,
    net313,
    net311,
    net310,
    net309,
    net308,
    net307,
    net306,
    net305,
    net304,
    net303,
    net302,
    net300,
    net299,
    net298,
    net297,
    net296,
    net295,
    net294,
    net293,
    net292,
    net291,
    net289,
    net288,
    net287,
    net286,
    net285,
    net284,
    net283,
    net282,
    net281,
    net280,
    net278,
    net277,
    net276,
    net275,
    net274,
    net273,
    net272,
    net271,
    net270,
    net269,
    net267,
    net266,
    net265,
    net264,
    net263,
    net262,
    net261,
    net260,
    net259,
    net258,
    net320,
    net319,
    net318,
    net317,
    net312,
    net301,
    net290,
    net279,
    net268,
    net257}),
    .io_ins_left({\ces_7_4_io_ins_left[63] ,
    \ces_7_4_io_ins_left[62] ,
    \ces_7_4_io_ins_left[61] ,
    \ces_7_4_io_ins_left[60] ,
    \ces_7_4_io_ins_left[59] ,
    \ces_7_4_io_ins_left[58] ,
    \ces_7_4_io_ins_left[57] ,
    \ces_7_4_io_ins_left[56] ,
    \ces_7_4_io_ins_left[55] ,
    \ces_7_4_io_ins_left[54] ,
    \ces_7_4_io_ins_left[53] ,
    \ces_7_4_io_ins_left[52] ,
    \ces_7_4_io_ins_left[51] ,
    \ces_7_4_io_ins_left[50] ,
    \ces_7_4_io_ins_left[49] ,
    \ces_7_4_io_ins_left[48] ,
    \ces_7_4_io_ins_left[47] ,
    \ces_7_4_io_ins_left[46] ,
    \ces_7_4_io_ins_left[45] ,
    \ces_7_4_io_ins_left[44] ,
    \ces_7_4_io_ins_left[43] ,
    \ces_7_4_io_ins_left[42] ,
    \ces_7_4_io_ins_left[41] ,
    \ces_7_4_io_ins_left[40] ,
    \ces_7_4_io_ins_left[39] ,
    \ces_7_4_io_ins_left[38] ,
    \ces_7_4_io_ins_left[37] ,
    \ces_7_4_io_ins_left[36] ,
    \ces_7_4_io_ins_left[35] ,
    \ces_7_4_io_ins_left[34] ,
    \ces_7_4_io_ins_left[33] ,
    \ces_7_4_io_ins_left[32] ,
    \ces_7_4_io_ins_left[31] ,
    \ces_7_4_io_ins_left[30] ,
    \ces_7_4_io_ins_left[29] ,
    \ces_7_4_io_ins_left[28] ,
    \ces_7_4_io_ins_left[27] ,
    \ces_7_4_io_ins_left[26] ,
    \ces_7_4_io_ins_left[25] ,
    \ces_7_4_io_ins_left[24] ,
    \ces_7_4_io_ins_left[23] ,
    \ces_7_4_io_ins_left[22] ,
    \ces_7_4_io_ins_left[21] ,
    \ces_7_4_io_ins_left[20] ,
    \ces_7_4_io_ins_left[19] ,
    \ces_7_4_io_ins_left[18] ,
    \ces_7_4_io_ins_left[17] ,
    \ces_7_4_io_ins_left[16] ,
    \ces_7_4_io_ins_left[15] ,
    \ces_7_4_io_ins_left[14] ,
    \ces_7_4_io_ins_left[13] ,
    \ces_7_4_io_ins_left[12] ,
    \ces_7_4_io_ins_left[11] ,
    \ces_7_4_io_ins_left[10] ,
    \ces_7_4_io_ins_left[9] ,
    \ces_7_4_io_ins_left[8] ,
    \ces_7_4_io_ins_left[7] ,
    \ces_7_4_io_ins_left[6] ,
    \ces_7_4_io_ins_left[5] ,
    \ces_7_4_io_ins_left[4] ,
    \ces_7_4_io_ins_left[3] ,
    \ces_7_4_io_ins_left[2] ,
    \ces_7_4_io_ins_left[1] ,
    \ces_7_4_io_ins_left[0] }),
    .io_ins_right({\ces_7_3_io_outs_right[63] ,
    \ces_7_3_io_outs_right[62] ,
    \ces_7_3_io_outs_right[61] ,
    \ces_7_3_io_outs_right[60] ,
    \ces_7_3_io_outs_right[59] ,
    \ces_7_3_io_outs_right[58] ,
    \ces_7_3_io_outs_right[57] ,
    \ces_7_3_io_outs_right[56] ,
    \ces_7_3_io_outs_right[55] ,
    \ces_7_3_io_outs_right[54] ,
    \ces_7_3_io_outs_right[53] ,
    \ces_7_3_io_outs_right[52] ,
    \ces_7_3_io_outs_right[51] ,
    \ces_7_3_io_outs_right[50] ,
    \ces_7_3_io_outs_right[49] ,
    \ces_7_3_io_outs_right[48] ,
    \ces_7_3_io_outs_right[47] ,
    \ces_7_3_io_outs_right[46] ,
    \ces_7_3_io_outs_right[45] ,
    \ces_7_3_io_outs_right[44] ,
    \ces_7_3_io_outs_right[43] ,
    \ces_7_3_io_outs_right[42] ,
    \ces_7_3_io_outs_right[41] ,
    \ces_7_3_io_outs_right[40] ,
    \ces_7_3_io_outs_right[39] ,
    \ces_7_3_io_outs_right[38] ,
    \ces_7_3_io_outs_right[37] ,
    \ces_7_3_io_outs_right[36] ,
    \ces_7_3_io_outs_right[35] ,
    \ces_7_3_io_outs_right[34] ,
    \ces_7_3_io_outs_right[33] ,
    \ces_7_3_io_outs_right[32] ,
    \ces_7_3_io_outs_right[31] ,
    \ces_7_3_io_outs_right[30] ,
    \ces_7_3_io_outs_right[29] ,
    \ces_7_3_io_outs_right[28] ,
    \ces_7_3_io_outs_right[27] ,
    \ces_7_3_io_outs_right[26] ,
    \ces_7_3_io_outs_right[25] ,
    \ces_7_3_io_outs_right[24] ,
    \ces_7_3_io_outs_right[23] ,
    \ces_7_3_io_outs_right[22] ,
    \ces_7_3_io_outs_right[21] ,
    \ces_7_3_io_outs_right[20] ,
    \ces_7_3_io_outs_right[19] ,
    \ces_7_3_io_outs_right[18] ,
    \ces_7_3_io_outs_right[17] ,
    \ces_7_3_io_outs_right[16] ,
    \ces_7_3_io_outs_right[15] ,
    \ces_7_3_io_outs_right[14] ,
    \ces_7_3_io_outs_right[13] ,
    \ces_7_3_io_outs_right[12] ,
    \ces_7_3_io_outs_right[11] ,
    \ces_7_3_io_outs_right[10] ,
    \ces_7_3_io_outs_right[9] ,
    \ces_7_3_io_outs_right[8] ,
    \ces_7_3_io_outs_right[7] ,
    \ces_7_3_io_outs_right[6] ,
    \ces_7_3_io_outs_right[5] ,
    \ces_7_3_io_outs_right[4] ,
    \ces_7_3_io_outs_right[3] ,
    \ces_7_3_io_outs_right[2] ,
    \ces_7_3_io_outs_right[1] ,
    \ces_7_3_io_outs_right[0] }),
    .io_ins_up({\ces_6_4_io_outs_up[63] ,
    \ces_6_4_io_outs_up[62] ,
    \ces_6_4_io_outs_up[61] ,
    \ces_6_4_io_outs_up[60] ,
    \ces_6_4_io_outs_up[59] ,
    \ces_6_4_io_outs_up[58] ,
    \ces_6_4_io_outs_up[57] ,
    \ces_6_4_io_outs_up[56] ,
    \ces_6_4_io_outs_up[55] ,
    \ces_6_4_io_outs_up[54] ,
    \ces_6_4_io_outs_up[53] ,
    \ces_6_4_io_outs_up[52] ,
    \ces_6_4_io_outs_up[51] ,
    \ces_6_4_io_outs_up[50] ,
    \ces_6_4_io_outs_up[49] ,
    \ces_6_4_io_outs_up[48] ,
    \ces_6_4_io_outs_up[47] ,
    \ces_6_4_io_outs_up[46] ,
    \ces_6_4_io_outs_up[45] ,
    \ces_6_4_io_outs_up[44] ,
    \ces_6_4_io_outs_up[43] ,
    \ces_6_4_io_outs_up[42] ,
    \ces_6_4_io_outs_up[41] ,
    \ces_6_4_io_outs_up[40] ,
    \ces_6_4_io_outs_up[39] ,
    \ces_6_4_io_outs_up[38] ,
    \ces_6_4_io_outs_up[37] ,
    \ces_6_4_io_outs_up[36] ,
    \ces_6_4_io_outs_up[35] ,
    \ces_6_4_io_outs_up[34] ,
    \ces_6_4_io_outs_up[33] ,
    \ces_6_4_io_outs_up[32] ,
    \ces_6_4_io_outs_up[31] ,
    \ces_6_4_io_outs_up[30] ,
    \ces_6_4_io_outs_up[29] ,
    \ces_6_4_io_outs_up[28] ,
    \ces_6_4_io_outs_up[27] ,
    \ces_6_4_io_outs_up[26] ,
    \ces_6_4_io_outs_up[25] ,
    \ces_6_4_io_outs_up[24] ,
    \ces_6_4_io_outs_up[23] ,
    \ces_6_4_io_outs_up[22] ,
    \ces_6_4_io_outs_up[21] ,
    \ces_6_4_io_outs_up[20] ,
    \ces_6_4_io_outs_up[19] ,
    \ces_6_4_io_outs_up[18] ,
    \ces_6_4_io_outs_up[17] ,
    \ces_6_4_io_outs_up[16] ,
    \ces_6_4_io_outs_up[15] ,
    \ces_6_4_io_outs_up[14] ,
    \ces_6_4_io_outs_up[13] ,
    \ces_6_4_io_outs_up[12] ,
    \ces_6_4_io_outs_up[11] ,
    \ces_6_4_io_outs_up[10] ,
    \ces_6_4_io_outs_up[9] ,
    \ces_6_4_io_outs_up[8] ,
    \ces_6_4_io_outs_up[7] ,
    \ces_6_4_io_outs_up[6] ,
    \ces_6_4_io_outs_up[5] ,
    \ces_6_4_io_outs_up[4] ,
    \ces_6_4_io_outs_up[3] ,
    \ces_6_4_io_outs_up[2] ,
    \ces_6_4_io_outs_up[1] ,
    \ces_6_4_io_outs_up[0] }),
    .io_outs_down({\ces_6_4_io_ins_down[63] ,
    \ces_6_4_io_ins_down[62] ,
    \ces_6_4_io_ins_down[61] ,
    \ces_6_4_io_ins_down[60] ,
    \ces_6_4_io_ins_down[59] ,
    \ces_6_4_io_ins_down[58] ,
    \ces_6_4_io_ins_down[57] ,
    \ces_6_4_io_ins_down[56] ,
    \ces_6_4_io_ins_down[55] ,
    \ces_6_4_io_ins_down[54] ,
    \ces_6_4_io_ins_down[53] ,
    \ces_6_4_io_ins_down[52] ,
    \ces_6_4_io_ins_down[51] ,
    \ces_6_4_io_ins_down[50] ,
    \ces_6_4_io_ins_down[49] ,
    \ces_6_4_io_ins_down[48] ,
    \ces_6_4_io_ins_down[47] ,
    \ces_6_4_io_ins_down[46] ,
    \ces_6_4_io_ins_down[45] ,
    \ces_6_4_io_ins_down[44] ,
    \ces_6_4_io_ins_down[43] ,
    \ces_6_4_io_ins_down[42] ,
    \ces_6_4_io_ins_down[41] ,
    \ces_6_4_io_ins_down[40] ,
    \ces_6_4_io_ins_down[39] ,
    \ces_6_4_io_ins_down[38] ,
    \ces_6_4_io_ins_down[37] ,
    \ces_6_4_io_ins_down[36] ,
    \ces_6_4_io_ins_down[35] ,
    \ces_6_4_io_ins_down[34] ,
    \ces_6_4_io_ins_down[33] ,
    \ces_6_4_io_ins_down[32] ,
    \ces_6_4_io_ins_down[31] ,
    \ces_6_4_io_ins_down[30] ,
    \ces_6_4_io_ins_down[29] ,
    \ces_6_4_io_ins_down[28] ,
    \ces_6_4_io_ins_down[27] ,
    \ces_6_4_io_ins_down[26] ,
    \ces_6_4_io_ins_down[25] ,
    \ces_6_4_io_ins_down[24] ,
    \ces_6_4_io_ins_down[23] ,
    \ces_6_4_io_ins_down[22] ,
    \ces_6_4_io_ins_down[21] ,
    \ces_6_4_io_ins_down[20] ,
    \ces_6_4_io_ins_down[19] ,
    \ces_6_4_io_ins_down[18] ,
    \ces_6_4_io_ins_down[17] ,
    \ces_6_4_io_ins_down[16] ,
    \ces_6_4_io_ins_down[15] ,
    \ces_6_4_io_ins_down[14] ,
    \ces_6_4_io_ins_down[13] ,
    \ces_6_4_io_ins_down[12] ,
    \ces_6_4_io_ins_down[11] ,
    \ces_6_4_io_ins_down[10] ,
    \ces_6_4_io_ins_down[9] ,
    \ces_6_4_io_ins_down[8] ,
    \ces_6_4_io_ins_down[7] ,
    \ces_6_4_io_ins_down[6] ,
    \ces_6_4_io_ins_down[5] ,
    \ces_6_4_io_ins_down[4] ,
    \ces_6_4_io_ins_down[3] ,
    \ces_6_4_io_ins_down[2] ,
    \ces_6_4_io_ins_down[1] ,
    \ces_6_4_io_ins_down[0] }),
    .io_outs_left({\ces_7_3_io_ins_left[63] ,
    \ces_7_3_io_ins_left[62] ,
    \ces_7_3_io_ins_left[61] ,
    \ces_7_3_io_ins_left[60] ,
    \ces_7_3_io_ins_left[59] ,
    \ces_7_3_io_ins_left[58] ,
    \ces_7_3_io_ins_left[57] ,
    \ces_7_3_io_ins_left[56] ,
    \ces_7_3_io_ins_left[55] ,
    \ces_7_3_io_ins_left[54] ,
    \ces_7_3_io_ins_left[53] ,
    \ces_7_3_io_ins_left[52] ,
    \ces_7_3_io_ins_left[51] ,
    \ces_7_3_io_ins_left[50] ,
    \ces_7_3_io_ins_left[49] ,
    \ces_7_3_io_ins_left[48] ,
    \ces_7_3_io_ins_left[47] ,
    \ces_7_3_io_ins_left[46] ,
    \ces_7_3_io_ins_left[45] ,
    \ces_7_3_io_ins_left[44] ,
    \ces_7_3_io_ins_left[43] ,
    \ces_7_3_io_ins_left[42] ,
    \ces_7_3_io_ins_left[41] ,
    \ces_7_3_io_ins_left[40] ,
    \ces_7_3_io_ins_left[39] ,
    \ces_7_3_io_ins_left[38] ,
    \ces_7_3_io_ins_left[37] ,
    \ces_7_3_io_ins_left[36] ,
    \ces_7_3_io_ins_left[35] ,
    \ces_7_3_io_ins_left[34] ,
    \ces_7_3_io_ins_left[33] ,
    \ces_7_3_io_ins_left[32] ,
    \ces_7_3_io_ins_left[31] ,
    \ces_7_3_io_ins_left[30] ,
    \ces_7_3_io_ins_left[29] ,
    \ces_7_3_io_ins_left[28] ,
    \ces_7_3_io_ins_left[27] ,
    \ces_7_3_io_ins_left[26] ,
    \ces_7_3_io_ins_left[25] ,
    \ces_7_3_io_ins_left[24] ,
    \ces_7_3_io_ins_left[23] ,
    \ces_7_3_io_ins_left[22] ,
    \ces_7_3_io_ins_left[21] ,
    \ces_7_3_io_ins_left[20] ,
    \ces_7_3_io_ins_left[19] ,
    \ces_7_3_io_ins_left[18] ,
    \ces_7_3_io_ins_left[17] ,
    \ces_7_3_io_ins_left[16] ,
    \ces_7_3_io_ins_left[15] ,
    \ces_7_3_io_ins_left[14] ,
    \ces_7_3_io_ins_left[13] ,
    \ces_7_3_io_ins_left[12] ,
    \ces_7_3_io_ins_left[11] ,
    \ces_7_3_io_ins_left[10] ,
    \ces_7_3_io_ins_left[9] ,
    \ces_7_3_io_ins_left[8] ,
    \ces_7_3_io_ins_left[7] ,
    \ces_7_3_io_ins_left[6] ,
    \ces_7_3_io_ins_left[5] ,
    \ces_7_3_io_ins_left[4] ,
    \ces_7_3_io_ins_left[3] ,
    \ces_7_3_io_ins_left[2] ,
    \ces_7_3_io_ins_left[1] ,
    \ces_7_3_io_ins_left[0] }),
    .io_outs_right({\ces_7_4_io_outs_right[63] ,
    \ces_7_4_io_outs_right[62] ,
    \ces_7_4_io_outs_right[61] ,
    \ces_7_4_io_outs_right[60] ,
    \ces_7_4_io_outs_right[59] ,
    \ces_7_4_io_outs_right[58] ,
    \ces_7_4_io_outs_right[57] ,
    \ces_7_4_io_outs_right[56] ,
    \ces_7_4_io_outs_right[55] ,
    \ces_7_4_io_outs_right[54] ,
    \ces_7_4_io_outs_right[53] ,
    \ces_7_4_io_outs_right[52] ,
    \ces_7_4_io_outs_right[51] ,
    \ces_7_4_io_outs_right[50] ,
    \ces_7_4_io_outs_right[49] ,
    \ces_7_4_io_outs_right[48] ,
    \ces_7_4_io_outs_right[47] ,
    \ces_7_4_io_outs_right[46] ,
    \ces_7_4_io_outs_right[45] ,
    \ces_7_4_io_outs_right[44] ,
    \ces_7_4_io_outs_right[43] ,
    \ces_7_4_io_outs_right[42] ,
    \ces_7_4_io_outs_right[41] ,
    \ces_7_4_io_outs_right[40] ,
    \ces_7_4_io_outs_right[39] ,
    \ces_7_4_io_outs_right[38] ,
    \ces_7_4_io_outs_right[37] ,
    \ces_7_4_io_outs_right[36] ,
    \ces_7_4_io_outs_right[35] ,
    \ces_7_4_io_outs_right[34] ,
    \ces_7_4_io_outs_right[33] ,
    \ces_7_4_io_outs_right[32] ,
    \ces_7_4_io_outs_right[31] ,
    \ces_7_4_io_outs_right[30] ,
    \ces_7_4_io_outs_right[29] ,
    \ces_7_4_io_outs_right[28] ,
    \ces_7_4_io_outs_right[27] ,
    \ces_7_4_io_outs_right[26] ,
    \ces_7_4_io_outs_right[25] ,
    \ces_7_4_io_outs_right[24] ,
    \ces_7_4_io_outs_right[23] ,
    \ces_7_4_io_outs_right[22] ,
    \ces_7_4_io_outs_right[21] ,
    \ces_7_4_io_outs_right[20] ,
    \ces_7_4_io_outs_right[19] ,
    \ces_7_4_io_outs_right[18] ,
    \ces_7_4_io_outs_right[17] ,
    \ces_7_4_io_outs_right[16] ,
    \ces_7_4_io_outs_right[15] ,
    \ces_7_4_io_outs_right[14] ,
    \ces_7_4_io_outs_right[13] ,
    \ces_7_4_io_outs_right[12] ,
    \ces_7_4_io_outs_right[11] ,
    \ces_7_4_io_outs_right[10] ,
    \ces_7_4_io_outs_right[9] ,
    \ces_7_4_io_outs_right[8] ,
    \ces_7_4_io_outs_right[7] ,
    \ces_7_4_io_outs_right[6] ,
    \ces_7_4_io_outs_right[5] ,
    \ces_7_4_io_outs_right[4] ,
    \ces_7_4_io_outs_right[3] ,
    \ces_7_4_io_outs_right[2] ,
    \ces_7_4_io_outs_right[1] ,
    \ces_7_4_io_outs_right[0] }),
    .io_outs_up({net3964,
    net3963,
    net3962,
    net3961,
    net3959,
    net3958,
    net3957,
    net3956,
    net3955,
    net3954,
    net3953,
    net3952,
    net3951,
    net3950,
    net3948,
    net3947,
    net3946,
    net3945,
    net3944,
    net3943,
    net3942,
    net3941,
    net3940,
    net3939,
    net3937,
    net3936,
    net3935,
    net3934,
    net3933,
    net3932,
    net3931,
    net3930,
    net3929,
    net3928,
    net3926,
    net3925,
    net3924,
    net3923,
    net3922,
    net3921,
    net3920,
    net3919,
    net3918,
    net3917,
    net3915,
    net3914,
    net3913,
    net3912,
    net3911,
    net3910,
    net3909,
    net3908,
    net3907,
    net3906,
    net3968,
    net3967,
    net3966,
    net3965,
    net3960,
    net3949,
    net3938,
    net3927,
    net3916,
    net3905}));
 Element ces_7_5 (.clock(clknet_3_7_0_clock),
    .io_lsbIns_1(ces_7_4_io_lsbOuts_1),
    .io_lsbIns_2(ces_7_4_io_lsbOuts_2),
    .io_lsbIns_3(ces_7_4_io_lsbOuts_3),
    .io_lsbIns_4(ces_7_4_io_lsbOuts_4),
    .io_lsbIns_5(ces_7_4_io_lsbOuts_5),
    .io_lsbIns_6(ces_7_4_io_lsbOuts_6),
    .io_lsbIns_7(ces_7_4_io_lsbOuts_7),
    .io_lsbOuts_0(ces_7_5_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_5_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_5_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_5_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_5_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_5_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_5_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_5_io_lsbOuts_7),
    .io_ins_down({net380,
    net379,
    net378,
    net377,
    net375,
    net374,
    net373,
    net372,
    net371,
    net370,
    net369,
    net368,
    net367,
    net366,
    net364,
    net363,
    net362,
    net361,
    net360,
    net359,
    net358,
    net357,
    net356,
    net355,
    net353,
    net352,
    net351,
    net350,
    net349,
    net348,
    net347,
    net346,
    net345,
    net344,
    net342,
    net341,
    net340,
    net339,
    net338,
    net337,
    net336,
    net335,
    net334,
    net333,
    net331,
    net330,
    net329,
    net328,
    net327,
    net326,
    net325,
    net324,
    net323,
    net322,
    net384,
    net383,
    net382,
    net381,
    net376,
    net365,
    net354,
    net343,
    net332,
    net321}),
    .io_ins_left({\ces_7_5_io_ins_left[63] ,
    \ces_7_5_io_ins_left[62] ,
    \ces_7_5_io_ins_left[61] ,
    \ces_7_5_io_ins_left[60] ,
    \ces_7_5_io_ins_left[59] ,
    \ces_7_5_io_ins_left[58] ,
    \ces_7_5_io_ins_left[57] ,
    \ces_7_5_io_ins_left[56] ,
    \ces_7_5_io_ins_left[55] ,
    \ces_7_5_io_ins_left[54] ,
    \ces_7_5_io_ins_left[53] ,
    \ces_7_5_io_ins_left[52] ,
    \ces_7_5_io_ins_left[51] ,
    \ces_7_5_io_ins_left[50] ,
    \ces_7_5_io_ins_left[49] ,
    \ces_7_5_io_ins_left[48] ,
    \ces_7_5_io_ins_left[47] ,
    \ces_7_5_io_ins_left[46] ,
    \ces_7_5_io_ins_left[45] ,
    \ces_7_5_io_ins_left[44] ,
    \ces_7_5_io_ins_left[43] ,
    \ces_7_5_io_ins_left[42] ,
    \ces_7_5_io_ins_left[41] ,
    \ces_7_5_io_ins_left[40] ,
    \ces_7_5_io_ins_left[39] ,
    \ces_7_5_io_ins_left[38] ,
    \ces_7_5_io_ins_left[37] ,
    \ces_7_5_io_ins_left[36] ,
    \ces_7_5_io_ins_left[35] ,
    \ces_7_5_io_ins_left[34] ,
    \ces_7_5_io_ins_left[33] ,
    \ces_7_5_io_ins_left[32] ,
    \ces_7_5_io_ins_left[31] ,
    \ces_7_5_io_ins_left[30] ,
    \ces_7_5_io_ins_left[29] ,
    \ces_7_5_io_ins_left[28] ,
    \ces_7_5_io_ins_left[27] ,
    \ces_7_5_io_ins_left[26] ,
    \ces_7_5_io_ins_left[25] ,
    \ces_7_5_io_ins_left[24] ,
    \ces_7_5_io_ins_left[23] ,
    \ces_7_5_io_ins_left[22] ,
    \ces_7_5_io_ins_left[21] ,
    \ces_7_5_io_ins_left[20] ,
    \ces_7_5_io_ins_left[19] ,
    \ces_7_5_io_ins_left[18] ,
    \ces_7_5_io_ins_left[17] ,
    \ces_7_5_io_ins_left[16] ,
    \ces_7_5_io_ins_left[15] ,
    \ces_7_5_io_ins_left[14] ,
    \ces_7_5_io_ins_left[13] ,
    \ces_7_5_io_ins_left[12] ,
    \ces_7_5_io_ins_left[11] ,
    \ces_7_5_io_ins_left[10] ,
    \ces_7_5_io_ins_left[9] ,
    \ces_7_5_io_ins_left[8] ,
    \ces_7_5_io_ins_left[7] ,
    \ces_7_5_io_ins_left[6] ,
    \ces_7_5_io_ins_left[5] ,
    \ces_7_5_io_ins_left[4] ,
    \ces_7_5_io_ins_left[3] ,
    \ces_7_5_io_ins_left[2] ,
    \ces_7_5_io_ins_left[1] ,
    \ces_7_5_io_ins_left[0] }),
    .io_ins_right({\ces_7_4_io_outs_right[63] ,
    \ces_7_4_io_outs_right[62] ,
    \ces_7_4_io_outs_right[61] ,
    \ces_7_4_io_outs_right[60] ,
    \ces_7_4_io_outs_right[59] ,
    \ces_7_4_io_outs_right[58] ,
    \ces_7_4_io_outs_right[57] ,
    \ces_7_4_io_outs_right[56] ,
    \ces_7_4_io_outs_right[55] ,
    \ces_7_4_io_outs_right[54] ,
    \ces_7_4_io_outs_right[53] ,
    \ces_7_4_io_outs_right[52] ,
    \ces_7_4_io_outs_right[51] ,
    \ces_7_4_io_outs_right[50] ,
    \ces_7_4_io_outs_right[49] ,
    \ces_7_4_io_outs_right[48] ,
    \ces_7_4_io_outs_right[47] ,
    \ces_7_4_io_outs_right[46] ,
    \ces_7_4_io_outs_right[45] ,
    \ces_7_4_io_outs_right[44] ,
    \ces_7_4_io_outs_right[43] ,
    \ces_7_4_io_outs_right[42] ,
    \ces_7_4_io_outs_right[41] ,
    \ces_7_4_io_outs_right[40] ,
    \ces_7_4_io_outs_right[39] ,
    \ces_7_4_io_outs_right[38] ,
    \ces_7_4_io_outs_right[37] ,
    \ces_7_4_io_outs_right[36] ,
    \ces_7_4_io_outs_right[35] ,
    \ces_7_4_io_outs_right[34] ,
    \ces_7_4_io_outs_right[33] ,
    \ces_7_4_io_outs_right[32] ,
    \ces_7_4_io_outs_right[31] ,
    \ces_7_4_io_outs_right[30] ,
    \ces_7_4_io_outs_right[29] ,
    \ces_7_4_io_outs_right[28] ,
    \ces_7_4_io_outs_right[27] ,
    \ces_7_4_io_outs_right[26] ,
    \ces_7_4_io_outs_right[25] ,
    \ces_7_4_io_outs_right[24] ,
    \ces_7_4_io_outs_right[23] ,
    \ces_7_4_io_outs_right[22] ,
    \ces_7_4_io_outs_right[21] ,
    \ces_7_4_io_outs_right[20] ,
    \ces_7_4_io_outs_right[19] ,
    \ces_7_4_io_outs_right[18] ,
    \ces_7_4_io_outs_right[17] ,
    \ces_7_4_io_outs_right[16] ,
    \ces_7_4_io_outs_right[15] ,
    \ces_7_4_io_outs_right[14] ,
    \ces_7_4_io_outs_right[13] ,
    \ces_7_4_io_outs_right[12] ,
    \ces_7_4_io_outs_right[11] ,
    \ces_7_4_io_outs_right[10] ,
    \ces_7_4_io_outs_right[9] ,
    \ces_7_4_io_outs_right[8] ,
    \ces_7_4_io_outs_right[7] ,
    \ces_7_4_io_outs_right[6] ,
    \ces_7_4_io_outs_right[5] ,
    \ces_7_4_io_outs_right[4] ,
    \ces_7_4_io_outs_right[3] ,
    \ces_7_4_io_outs_right[2] ,
    \ces_7_4_io_outs_right[1] ,
    \ces_7_4_io_outs_right[0] }),
    .io_ins_up({\ces_6_5_io_outs_up[63] ,
    \ces_6_5_io_outs_up[62] ,
    \ces_6_5_io_outs_up[61] ,
    \ces_6_5_io_outs_up[60] ,
    \ces_6_5_io_outs_up[59] ,
    \ces_6_5_io_outs_up[58] ,
    \ces_6_5_io_outs_up[57] ,
    \ces_6_5_io_outs_up[56] ,
    \ces_6_5_io_outs_up[55] ,
    \ces_6_5_io_outs_up[54] ,
    \ces_6_5_io_outs_up[53] ,
    \ces_6_5_io_outs_up[52] ,
    \ces_6_5_io_outs_up[51] ,
    \ces_6_5_io_outs_up[50] ,
    \ces_6_5_io_outs_up[49] ,
    \ces_6_5_io_outs_up[48] ,
    \ces_6_5_io_outs_up[47] ,
    \ces_6_5_io_outs_up[46] ,
    \ces_6_5_io_outs_up[45] ,
    \ces_6_5_io_outs_up[44] ,
    \ces_6_5_io_outs_up[43] ,
    \ces_6_5_io_outs_up[42] ,
    \ces_6_5_io_outs_up[41] ,
    \ces_6_5_io_outs_up[40] ,
    \ces_6_5_io_outs_up[39] ,
    \ces_6_5_io_outs_up[38] ,
    \ces_6_5_io_outs_up[37] ,
    \ces_6_5_io_outs_up[36] ,
    \ces_6_5_io_outs_up[35] ,
    \ces_6_5_io_outs_up[34] ,
    \ces_6_5_io_outs_up[33] ,
    \ces_6_5_io_outs_up[32] ,
    \ces_6_5_io_outs_up[31] ,
    \ces_6_5_io_outs_up[30] ,
    \ces_6_5_io_outs_up[29] ,
    \ces_6_5_io_outs_up[28] ,
    \ces_6_5_io_outs_up[27] ,
    \ces_6_5_io_outs_up[26] ,
    \ces_6_5_io_outs_up[25] ,
    \ces_6_5_io_outs_up[24] ,
    \ces_6_5_io_outs_up[23] ,
    \ces_6_5_io_outs_up[22] ,
    \ces_6_5_io_outs_up[21] ,
    \ces_6_5_io_outs_up[20] ,
    \ces_6_5_io_outs_up[19] ,
    \ces_6_5_io_outs_up[18] ,
    \ces_6_5_io_outs_up[17] ,
    \ces_6_5_io_outs_up[16] ,
    \ces_6_5_io_outs_up[15] ,
    \ces_6_5_io_outs_up[14] ,
    \ces_6_5_io_outs_up[13] ,
    \ces_6_5_io_outs_up[12] ,
    \ces_6_5_io_outs_up[11] ,
    \ces_6_5_io_outs_up[10] ,
    \ces_6_5_io_outs_up[9] ,
    \ces_6_5_io_outs_up[8] ,
    \ces_6_5_io_outs_up[7] ,
    \ces_6_5_io_outs_up[6] ,
    \ces_6_5_io_outs_up[5] ,
    \ces_6_5_io_outs_up[4] ,
    \ces_6_5_io_outs_up[3] ,
    \ces_6_5_io_outs_up[2] ,
    \ces_6_5_io_outs_up[1] ,
    \ces_6_5_io_outs_up[0] }),
    .io_outs_down({\ces_6_5_io_ins_down[63] ,
    \ces_6_5_io_ins_down[62] ,
    \ces_6_5_io_ins_down[61] ,
    \ces_6_5_io_ins_down[60] ,
    \ces_6_5_io_ins_down[59] ,
    \ces_6_5_io_ins_down[58] ,
    \ces_6_5_io_ins_down[57] ,
    \ces_6_5_io_ins_down[56] ,
    \ces_6_5_io_ins_down[55] ,
    \ces_6_5_io_ins_down[54] ,
    \ces_6_5_io_ins_down[53] ,
    \ces_6_5_io_ins_down[52] ,
    \ces_6_5_io_ins_down[51] ,
    \ces_6_5_io_ins_down[50] ,
    \ces_6_5_io_ins_down[49] ,
    \ces_6_5_io_ins_down[48] ,
    \ces_6_5_io_ins_down[47] ,
    \ces_6_5_io_ins_down[46] ,
    \ces_6_5_io_ins_down[45] ,
    \ces_6_5_io_ins_down[44] ,
    \ces_6_5_io_ins_down[43] ,
    \ces_6_5_io_ins_down[42] ,
    \ces_6_5_io_ins_down[41] ,
    \ces_6_5_io_ins_down[40] ,
    \ces_6_5_io_ins_down[39] ,
    \ces_6_5_io_ins_down[38] ,
    \ces_6_5_io_ins_down[37] ,
    \ces_6_5_io_ins_down[36] ,
    \ces_6_5_io_ins_down[35] ,
    \ces_6_5_io_ins_down[34] ,
    \ces_6_5_io_ins_down[33] ,
    \ces_6_5_io_ins_down[32] ,
    \ces_6_5_io_ins_down[31] ,
    \ces_6_5_io_ins_down[30] ,
    \ces_6_5_io_ins_down[29] ,
    \ces_6_5_io_ins_down[28] ,
    \ces_6_5_io_ins_down[27] ,
    \ces_6_5_io_ins_down[26] ,
    \ces_6_5_io_ins_down[25] ,
    \ces_6_5_io_ins_down[24] ,
    \ces_6_5_io_ins_down[23] ,
    \ces_6_5_io_ins_down[22] ,
    \ces_6_5_io_ins_down[21] ,
    \ces_6_5_io_ins_down[20] ,
    \ces_6_5_io_ins_down[19] ,
    \ces_6_5_io_ins_down[18] ,
    \ces_6_5_io_ins_down[17] ,
    \ces_6_5_io_ins_down[16] ,
    \ces_6_5_io_ins_down[15] ,
    \ces_6_5_io_ins_down[14] ,
    \ces_6_5_io_ins_down[13] ,
    \ces_6_5_io_ins_down[12] ,
    \ces_6_5_io_ins_down[11] ,
    \ces_6_5_io_ins_down[10] ,
    \ces_6_5_io_ins_down[9] ,
    \ces_6_5_io_ins_down[8] ,
    \ces_6_5_io_ins_down[7] ,
    \ces_6_5_io_ins_down[6] ,
    \ces_6_5_io_ins_down[5] ,
    \ces_6_5_io_ins_down[4] ,
    \ces_6_5_io_ins_down[3] ,
    \ces_6_5_io_ins_down[2] ,
    \ces_6_5_io_ins_down[1] ,
    \ces_6_5_io_ins_down[0] }),
    .io_outs_left({\ces_7_4_io_ins_left[63] ,
    \ces_7_4_io_ins_left[62] ,
    \ces_7_4_io_ins_left[61] ,
    \ces_7_4_io_ins_left[60] ,
    \ces_7_4_io_ins_left[59] ,
    \ces_7_4_io_ins_left[58] ,
    \ces_7_4_io_ins_left[57] ,
    \ces_7_4_io_ins_left[56] ,
    \ces_7_4_io_ins_left[55] ,
    \ces_7_4_io_ins_left[54] ,
    \ces_7_4_io_ins_left[53] ,
    \ces_7_4_io_ins_left[52] ,
    \ces_7_4_io_ins_left[51] ,
    \ces_7_4_io_ins_left[50] ,
    \ces_7_4_io_ins_left[49] ,
    \ces_7_4_io_ins_left[48] ,
    \ces_7_4_io_ins_left[47] ,
    \ces_7_4_io_ins_left[46] ,
    \ces_7_4_io_ins_left[45] ,
    \ces_7_4_io_ins_left[44] ,
    \ces_7_4_io_ins_left[43] ,
    \ces_7_4_io_ins_left[42] ,
    \ces_7_4_io_ins_left[41] ,
    \ces_7_4_io_ins_left[40] ,
    \ces_7_4_io_ins_left[39] ,
    \ces_7_4_io_ins_left[38] ,
    \ces_7_4_io_ins_left[37] ,
    \ces_7_4_io_ins_left[36] ,
    \ces_7_4_io_ins_left[35] ,
    \ces_7_4_io_ins_left[34] ,
    \ces_7_4_io_ins_left[33] ,
    \ces_7_4_io_ins_left[32] ,
    \ces_7_4_io_ins_left[31] ,
    \ces_7_4_io_ins_left[30] ,
    \ces_7_4_io_ins_left[29] ,
    \ces_7_4_io_ins_left[28] ,
    \ces_7_4_io_ins_left[27] ,
    \ces_7_4_io_ins_left[26] ,
    \ces_7_4_io_ins_left[25] ,
    \ces_7_4_io_ins_left[24] ,
    \ces_7_4_io_ins_left[23] ,
    \ces_7_4_io_ins_left[22] ,
    \ces_7_4_io_ins_left[21] ,
    \ces_7_4_io_ins_left[20] ,
    \ces_7_4_io_ins_left[19] ,
    \ces_7_4_io_ins_left[18] ,
    \ces_7_4_io_ins_left[17] ,
    \ces_7_4_io_ins_left[16] ,
    \ces_7_4_io_ins_left[15] ,
    \ces_7_4_io_ins_left[14] ,
    \ces_7_4_io_ins_left[13] ,
    \ces_7_4_io_ins_left[12] ,
    \ces_7_4_io_ins_left[11] ,
    \ces_7_4_io_ins_left[10] ,
    \ces_7_4_io_ins_left[9] ,
    \ces_7_4_io_ins_left[8] ,
    \ces_7_4_io_ins_left[7] ,
    \ces_7_4_io_ins_left[6] ,
    \ces_7_4_io_ins_left[5] ,
    \ces_7_4_io_ins_left[4] ,
    \ces_7_4_io_ins_left[3] ,
    \ces_7_4_io_ins_left[2] ,
    \ces_7_4_io_ins_left[1] ,
    \ces_7_4_io_ins_left[0] }),
    .io_outs_right({\ces_7_5_io_outs_right[63] ,
    \ces_7_5_io_outs_right[62] ,
    \ces_7_5_io_outs_right[61] ,
    \ces_7_5_io_outs_right[60] ,
    \ces_7_5_io_outs_right[59] ,
    \ces_7_5_io_outs_right[58] ,
    \ces_7_5_io_outs_right[57] ,
    \ces_7_5_io_outs_right[56] ,
    \ces_7_5_io_outs_right[55] ,
    \ces_7_5_io_outs_right[54] ,
    \ces_7_5_io_outs_right[53] ,
    \ces_7_5_io_outs_right[52] ,
    \ces_7_5_io_outs_right[51] ,
    \ces_7_5_io_outs_right[50] ,
    \ces_7_5_io_outs_right[49] ,
    \ces_7_5_io_outs_right[48] ,
    \ces_7_5_io_outs_right[47] ,
    \ces_7_5_io_outs_right[46] ,
    \ces_7_5_io_outs_right[45] ,
    \ces_7_5_io_outs_right[44] ,
    \ces_7_5_io_outs_right[43] ,
    \ces_7_5_io_outs_right[42] ,
    \ces_7_5_io_outs_right[41] ,
    \ces_7_5_io_outs_right[40] ,
    \ces_7_5_io_outs_right[39] ,
    \ces_7_5_io_outs_right[38] ,
    \ces_7_5_io_outs_right[37] ,
    \ces_7_5_io_outs_right[36] ,
    \ces_7_5_io_outs_right[35] ,
    \ces_7_5_io_outs_right[34] ,
    \ces_7_5_io_outs_right[33] ,
    \ces_7_5_io_outs_right[32] ,
    \ces_7_5_io_outs_right[31] ,
    \ces_7_5_io_outs_right[30] ,
    \ces_7_5_io_outs_right[29] ,
    \ces_7_5_io_outs_right[28] ,
    \ces_7_5_io_outs_right[27] ,
    \ces_7_5_io_outs_right[26] ,
    \ces_7_5_io_outs_right[25] ,
    \ces_7_5_io_outs_right[24] ,
    \ces_7_5_io_outs_right[23] ,
    \ces_7_5_io_outs_right[22] ,
    \ces_7_5_io_outs_right[21] ,
    \ces_7_5_io_outs_right[20] ,
    \ces_7_5_io_outs_right[19] ,
    \ces_7_5_io_outs_right[18] ,
    \ces_7_5_io_outs_right[17] ,
    \ces_7_5_io_outs_right[16] ,
    \ces_7_5_io_outs_right[15] ,
    \ces_7_5_io_outs_right[14] ,
    \ces_7_5_io_outs_right[13] ,
    \ces_7_5_io_outs_right[12] ,
    \ces_7_5_io_outs_right[11] ,
    \ces_7_5_io_outs_right[10] ,
    \ces_7_5_io_outs_right[9] ,
    \ces_7_5_io_outs_right[8] ,
    \ces_7_5_io_outs_right[7] ,
    \ces_7_5_io_outs_right[6] ,
    \ces_7_5_io_outs_right[5] ,
    \ces_7_5_io_outs_right[4] ,
    \ces_7_5_io_outs_right[3] ,
    \ces_7_5_io_outs_right[2] ,
    \ces_7_5_io_outs_right[1] ,
    \ces_7_5_io_outs_right[0] }),
    .io_outs_up({net4028,
    net4027,
    net4026,
    net4025,
    net4023,
    net4022,
    net4021,
    net4020,
    net4019,
    net4018,
    net4017,
    net4016,
    net4015,
    net4014,
    net4012,
    net4011,
    net4010,
    net4009,
    net4008,
    net4007,
    net4006,
    net4005,
    net4004,
    net4003,
    net4001,
    net4000,
    net3999,
    net3998,
    net3997,
    net3996,
    net3995,
    net3994,
    net3993,
    net3992,
    net3990,
    net3989,
    net3988,
    net3987,
    net3986,
    net3985,
    net3984,
    net3983,
    net3982,
    net3981,
    net3979,
    net3978,
    net3977,
    net3976,
    net3975,
    net3974,
    net3973,
    net3972,
    net3971,
    net3970,
    net4032,
    net4031,
    net4030,
    net4029,
    net4024,
    net4013,
    net4002,
    net3991,
    net3980,
    net3969}));
 Element ces_7_6 (.clock(clknet_3_7_0_clock),
    .io_lsbIns_1(ces_7_5_io_lsbOuts_1),
    .io_lsbIns_2(ces_7_5_io_lsbOuts_2),
    .io_lsbIns_3(ces_7_5_io_lsbOuts_3),
    .io_lsbIns_4(ces_7_5_io_lsbOuts_4),
    .io_lsbIns_5(ces_7_5_io_lsbOuts_5),
    .io_lsbIns_6(ces_7_5_io_lsbOuts_6),
    .io_lsbIns_7(ces_7_5_io_lsbOuts_7),
    .io_lsbOuts_0(ces_7_6_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_6_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_6_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_6_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_6_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_6_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_6_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_6_io_lsbOuts_7),
    .io_ins_down({net444,
    net443,
    net442,
    net441,
    net439,
    net438,
    net437,
    net436,
    net435,
    net434,
    net433,
    net432,
    net431,
    net430,
    net428,
    net427,
    net426,
    net425,
    net424,
    net423,
    net422,
    net421,
    net420,
    net419,
    net417,
    net416,
    net415,
    net414,
    net413,
    net412,
    net411,
    net410,
    net409,
    net408,
    net406,
    net405,
    net404,
    net403,
    net402,
    net401,
    net400,
    net399,
    net398,
    net397,
    net395,
    net394,
    net393,
    net392,
    net391,
    net390,
    net389,
    net388,
    net387,
    net386,
    net448,
    net447,
    net446,
    net445,
    net440,
    net429,
    net418,
    net407,
    net396,
    net385}),
    .io_ins_left({\ces_7_6_io_ins_left[63] ,
    \ces_7_6_io_ins_left[62] ,
    \ces_7_6_io_ins_left[61] ,
    \ces_7_6_io_ins_left[60] ,
    \ces_7_6_io_ins_left[59] ,
    \ces_7_6_io_ins_left[58] ,
    \ces_7_6_io_ins_left[57] ,
    \ces_7_6_io_ins_left[56] ,
    \ces_7_6_io_ins_left[55] ,
    \ces_7_6_io_ins_left[54] ,
    \ces_7_6_io_ins_left[53] ,
    \ces_7_6_io_ins_left[52] ,
    \ces_7_6_io_ins_left[51] ,
    \ces_7_6_io_ins_left[50] ,
    \ces_7_6_io_ins_left[49] ,
    \ces_7_6_io_ins_left[48] ,
    \ces_7_6_io_ins_left[47] ,
    \ces_7_6_io_ins_left[46] ,
    \ces_7_6_io_ins_left[45] ,
    \ces_7_6_io_ins_left[44] ,
    \ces_7_6_io_ins_left[43] ,
    \ces_7_6_io_ins_left[42] ,
    \ces_7_6_io_ins_left[41] ,
    \ces_7_6_io_ins_left[40] ,
    \ces_7_6_io_ins_left[39] ,
    \ces_7_6_io_ins_left[38] ,
    \ces_7_6_io_ins_left[37] ,
    \ces_7_6_io_ins_left[36] ,
    \ces_7_6_io_ins_left[35] ,
    \ces_7_6_io_ins_left[34] ,
    \ces_7_6_io_ins_left[33] ,
    \ces_7_6_io_ins_left[32] ,
    \ces_7_6_io_ins_left[31] ,
    \ces_7_6_io_ins_left[30] ,
    \ces_7_6_io_ins_left[29] ,
    \ces_7_6_io_ins_left[28] ,
    \ces_7_6_io_ins_left[27] ,
    \ces_7_6_io_ins_left[26] ,
    \ces_7_6_io_ins_left[25] ,
    \ces_7_6_io_ins_left[24] ,
    \ces_7_6_io_ins_left[23] ,
    \ces_7_6_io_ins_left[22] ,
    \ces_7_6_io_ins_left[21] ,
    \ces_7_6_io_ins_left[20] ,
    \ces_7_6_io_ins_left[19] ,
    \ces_7_6_io_ins_left[18] ,
    \ces_7_6_io_ins_left[17] ,
    \ces_7_6_io_ins_left[16] ,
    \ces_7_6_io_ins_left[15] ,
    \ces_7_6_io_ins_left[14] ,
    \ces_7_6_io_ins_left[13] ,
    \ces_7_6_io_ins_left[12] ,
    \ces_7_6_io_ins_left[11] ,
    \ces_7_6_io_ins_left[10] ,
    \ces_7_6_io_ins_left[9] ,
    \ces_7_6_io_ins_left[8] ,
    \ces_7_6_io_ins_left[7] ,
    \ces_7_6_io_ins_left[6] ,
    \ces_7_6_io_ins_left[5] ,
    \ces_7_6_io_ins_left[4] ,
    \ces_7_6_io_ins_left[3] ,
    \ces_7_6_io_ins_left[2] ,
    \ces_7_6_io_ins_left[1] ,
    \ces_7_6_io_ins_left[0] }),
    .io_ins_right({\ces_7_5_io_outs_right[63] ,
    \ces_7_5_io_outs_right[62] ,
    \ces_7_5_io_outs_right[61] ,
    \ces_7_5_io_outs_right[60] ,
    \ces_7_5_io_outs_right[59] ,
    \ces_7_5_io_outs_right[58] ,
    \ces_7_5_io_outs_right[57] ,
    \ces_7_5_io_outs_right[56] ,
    \ces_7_5_io_outs_right[55] ,
    \ces_7_5_io_outs_right[54] ,
    \ces_7_5_io_outs_right[53] ,
    \ces_7_5_io_outs_right[52] ,
    \ces_7_5_io_outs_right[51] ,
    \ces_7_5_io_outs_right[50] ,
    \ces_7_5_io_outs_right[49] ,
    \ces_7_5_io_outs_right[48] ,
    \ces_7_5_io_outs_right[47] ,
    \ces_7_5_io_outs_right[46] ,
    \ces_7_5_io_outs_right[45] ,
    \ces_7_5_io_outs_right[44] ,
    \ces_7_5_io_outs_right[43] ,
    \ces_7_5_io_outs_right[42] ,
    \ces_7_5_io_outs_right[41] ,
    \ces_7_5_io_outs_right[40] ,
    \ces_7_5_io_outs_right[39] ,
    \ces_7_5_io_outs_right[38] ,
    \ces_7_5_io_outs_right[37] ,
    \ces_7_5_io_outs_right[36] ,
    \ces_7_5_io_outs_right[35] ,
    \ces_7_5_io_outs_right[34] ,
    \ces_7_5_io_outs_right[33] ,
    \ces_7_5_io_outs_right[32] ,
    \ces_7_5_io_outs_right[31] ,
    \ces_7_5_io_outs_right[30] ,
    \ces_7_5_io_outs_right[29] ,
    \ces_7_5_io_outs_right[28] ,
    \ces_7_5_io_outs_right[27] ,
    \ces_7_5_io_outs_right[26] ,
    \ces_7_5_io_outs_right[25] ,
    \ces_7_5_io_outs_right[24] ,
    \ces_7_5_io_outs_right[23] ,
    \ces_7_5_io_outs_right[22] ,
    \ces_7_5_io_outs_right[21] ,
    \ces_7_5_io_outs_right[20] ,
    \ces_7_5_io_outs_right[19] ,
    \ces_7_5_io_outs_right[18] ,
    \ces_7_5_io_outs_right[17] ,
    \ces_7_5_io_outs_right[16] ,
    \ces_7_5_io_outs_right[15] ,
    \ces_7_5_io_outs_right[14] ,
    \ces_7_5_io_outs_right[13] ,
    \ces_7_5_io_outs_right[12] ,
    \ces_7_5_io_outs_right[11] ,
    \ces_7_5_io_outs_right[10] ,
    \ces_7_5_io_outs_right[9] ,
    \ces_7_5_io_outs_right[8] ,
    \ces_7_5_io_outs_right[7] ,
    \ces_7_5_io_outs_right[6] ,
    \ces_7_5_io_outs_right[5] ,
    \ces_7_5_io_outs_right[4] ,
    \ces_7_5_io_outs_right[3] ,
    \ces_7_5_io_outs_right[2] ,
    \ces_7_5_io_outs_right[1] ,
    \ces_7_5_io_outs_right[0] }),
    .io_ins_up({\ces_6_6_io_outs_up[63] ,
    \ces_6_6_io_outs_up[62] ,
    \ces_6_6_io_outs_up[61] ,
    \ces_6_6_io_outs_up[60] ,
    \ces_6_6_io_outs_up[59] ,
    \ces_6_6_io_outs_up[58] ,
    \ces_6_6_io_outs_up[57] ,
    \ces_6_6_io_outs_up[56] ,
    \ces_6_6_io_outs_up[55] ,
    \ces_6_6_io_outs_up[54] ,
    \ces_6_6_io_outs_up[53] ,
    \ces_6_6_io_outs_up[52] ,
    \ces_6_6_io_outs_up[51] ,
    \ces_6_6_io_outs_up[50] ,
    \ces_6_6_io_outs_up[49] ,
    \ces_6_6_io_outs_up[48] ,
    \ces_6_6_io_outs_up[47] ,
    \ces_6_6_io_outs_up[46] ,
    \ces_6_6_io_outs_up[45] ,
    \ces_6_6_io_outs_up[44] ,
    \ces_6_6_io_outs_up[43] ,
    \ces_6_6_io_outs_up[42] ,
    \ces_6_6_io_outs_up[41] ,
    \ces_6_6_io_outs_up[40] ,
    \ces_6_6_io_outs_up[39] ,
    \ces_6_6_io_outs_up[38] ,
    \ces_6_6_io_outs_up[37] ,
    \ces_6_6_io_outs_up[36] ,
    \ces_6_6_io_outs_up[35] ,
    \ces_6_6_io_outs_up[34] ,
    \ces_6_6_io_outs_up[33] ,
    \ces_6_6_io_outs_up[32] ,
    \ces_6_6_io_outs_up[31] ,
    \ces_6_6_io_outs_up[30] ,
    \ces_6_6_io_outs_up[29] ,
    \ces_6_6_io_outs_up[28] ,
    \ces_6_6_io_outs_up[27] ,
    \ces_6_6_io_outs_up[26] ,
    \ces_6_6_io_outs_up[25] ,
    \ces_6_6_io_outs_up[24] ,
    \ces_6_6_io_outs_up[23] ,
    \ces_6_6_io_outs_up[22] ,
    \ces_6_6_io_outs_up[21] ,
    \ces_6_6_io_outs_up[20] ,
    \ces_6_6_io_outs_up[19] ,
    \ces_6_6_io_outs_up[18] ,
    \ces_6_6_io_outs_up[17] ,
    \ces_6_6_io_outs_up[16] ,
    \ces_6_6_io_outs_up[15] ,
    \ces_6_6_io_outs_up[14] ,
    \ces_6_6_io_outs_up[13] ,
    \ces_6_6_io_outs_up[12] ,
    \ces_6_6_io_outs_up[11] ,
    \ces_6_6_io_outs_up[10] ,
    \ces_6_6_io_outs_up[9] ,
    \ces_6_6_io_outs_up[8] ,
    \ces_6_6_io_outs_up[7] ,
    \ces_6_6_io_outs_up[6] ,
    \ces_6_6_io_outs_up[5] ,
    \ces_6_6_io_outs_up[4] ,
    \ces_6_6_io_outs_up[3] ,
    \ces_6_6_io_outs_up[2] ,
    \ces_6_6_io_outs_up[1] ,
    \ces_6_6_io_outs_up[0] }),
    .io_outs_down({\ces_6_6_io_ins_down[63] ,
    \ces_6_6_io_ins_down[62] ,
    \ces_6_6_io_ins_down[61] ,
    \ces_6_6_io_ins_down[60] ,
    \ces_6_6_io_ins_down[59] ,
    \ces_6_6_io_ins_down[58] ,
    \ces_6_6_io_ins_down[57] ,
    \ces_6_6_io_ins_down[56] ,
    \ces_6_6_io_ins_down[55] ,
    \ces_6_6_io_ins_down[54] ,
    \ces_6_6_io_ins_down[53] ,
    \ces_6_6_io_ins_down[52] ,
    \ces_6_6_io_ins_down[51] ,
    \ces_6_6_io_ins_down[50] ,
    \ces_6_6_io_ins_down[49] ,
    \ces_6_6_io_ins_down[48] ,
    \ces_6_6_io_ins_down[47] ,
    \ces_6_6_io_ins_down[46] ,
    \ces_6_6_io_ins_down[45] ,
    \ces_6_6_io_ins_down[44] ,
    \ces_6_6_io_ins_down[43] ,
    \ces_6_6_io_ins_down[42] ,
    \ces_6_6_io_ins_down[41] ,
    \ces_6_6_io_ins_down[40] ,
    \ces_6_6_io_ins_down[39] ,
    \ces_6_6_io_ins_down[38] ,
    \ces_6_6_io_ins_down[37] ,
    \ces_6_6_io_ins_down[36] ,
    \ces_6_6_io_ins_down[35] ,
    \ces_6_6_io_ins_down[34] ,
    \ces_6_6_io_ins_down[33] ,
    \ces_6_6_io_ins_down[32] ,
    \ces_6_6_io_ins_down[31] ,
    \ces_6_6_io_ins_down[30] ,
    \ces_6_6_io_ins_down[29] ,
    \ces_6_6_io_ins_down[28] ,
    \ces_6_6_io_ins_down[27] ,
    \ces_6_6_io_ins_down[26] ,
    \ces_6_6_io_ins_down[25] ,
    \ces_6_6_io_ins_down[24] ,
    \ces_6_6_io_ins_down[23] ,
    \ces_6_6_io_ins_down[22] ,
    \ces_6_6_io_ins_down[21] ,
    \ces_6_6_io_ins_down[20] ,
    \ces_6_6_io_ins_down[19] ,
    \ces_6_6_io_ins_down[18] ,
    \ces_6_6_io_ins_down[17] ,
    \ces_6_6_io_ins_down[16] ,
    \ces_6_6_io_ins_down[15] ,
    \ces_6_6_io_ins_down[14] ,
    \ces_6_6_io_ins_down[13] ,
    \ces_6_6_io_ins_down[12] ,
    \ces_6_6_io_ins_down[11] ,
    \ces_6_6_io_ins_down[10] ,
    \ces_6_6_io_ins_down[9] ,
    \ces_6_6_io_ins_down[8] ,
    \ces_6_6_io_ins_down[7] ,
    \ces_6_6_io_ins_down[6] ,
    \ces_6_6_io_ins_down[5] ,
    \ces_6_6_io_ins_down[4] ,
    \ces_6_6_io_ins_down[3] ,
    \ces_6_6_io_ins_down[2] ,
    \ces_6_6_io_ins_down[1] ,
    \ces_6_6_io_ins_down[0] }),
    .io_outs_left({\ces_7_5_io_ins_left[63] ,
    \ces_7_5_io_ins_left[62] ,
    \ces_7_5_io_ins_left[61] ,
    \ces_7_5_io_ins_left[60] ,
    \ces_7_5_io_ins_left[59] ,
    \ces_7_5_io_ins_left[58] ,
    \ces_7_5_io_ins_left[57] ,
    \ces_7_5_io_ins_left[56] ,
    \ces_7_5_io_ins_left[55] ,
    \ces_7_5_io_ins_left[54] ,
    \ces_7_5_io_ins_left[53] ,
    \ces_7_5_io_ins_left[52] ,
    \ces_7_5_io_ins_left[51] ,
    \ces_7_5_io_ins_left[50] ,
    \ces_7_5_io_ins_left[49] ,
    \ces_7_5_io_ins_left[48] ,
    \ces_7_5_io_ins_left[47] ,
    \ces_7_5_io_ins_left[46] ,
    \ces_7_5_io_ins_left[45] ,
    \ces_7_5_io_ins_left[44] ,
    \ces_7_5_io_ins_left[43] ,
    \ces_7_5_io_ins_left[42] ,
    \ces_7_5_io_ins_left[41] ,
    \ces_7_5_io_ins_left[40] ,
    \ces_7_5_io_ins_left[39] ,
    \ces_7_5_io_ins_left[38] ,
    \ces_7_5_io_ins_left[37] ,
    \ces_7_5_io_ins_left[36] ,
    \ces_7_5_io_ins_left[35] ,
    \ces_7_5_io_ins_left[34] ,
    \ces_7_5_io_ins_left[33] ,
    \ces_7_5_io_ins_left[32] ,
    \ces_7_5_io_ins_left[31] ,
    \ces_7_5_io_ins_left[30] ,
    \ces_7_5_io_ins_left[29] ,
    \ces_7_5_io_ins_left[28] ,
    \ces_7_5_io_ins_left[27] ,
    \ces_7_5_io_ins_left[26] ,
    \ces_7_5_io_ins_left[25] ,
    \ces_7_5_io_ins_left[24] ,
    \ces_7_5_io_ins_left[23] ,
    \ces_7_5_io_ins_left[22] ,
    \ces_7_5_io_ins_left[21] ,
    \ces_7_5_io_ins_left[20] ,
    \ces_7_5_io_ins_left[19] ,
    \ces_7_5_io_ins_left[18] ,
    \ces_7_5_io_ins_left[17] ,
    \ces_7_5_io_ins_left[16] ,
    \ces_7_5_io_ins_left[15] ,
    \ces_7_5_io_ins_left[14] ,
    \ces_7_5_io_ins_left[13] ,
    \ces_7_5_io_ins_left[12] ,
    \ces_7_5_io_ins_left[11] ,
    \ces_7_5_io_ins_left[10] ,
    \ces_7_5_io_ins_left[9] ,
    \ces_7_5_io_ins_left[8] ,
    \ces_7_5_io_ins_left[7] ,
    \ces_7_5_io_ins_left[6] ,
    \ces_7_5_io_ins_left[5] ,
    \ces_7_5_io_ins_left[4] ,
    \ces_7_5_io_ins_left[3] ,
    \ces_7_5_io_ins_left[2] ,
    \ces_7_5_io_ins_left[1] ,
    \ces_7_5_io_ins_left[0] }),
    .io_outs_right({\ces_7_6_io_outs_right[63] ,
    \ces_7_6_io_outs_right[62] ,
    \ces_7_6_io_outs_right[61] ,
    \ces_7_6_io_outs_right[60] ,
    \ces_7_6_io_outs_right[59] ,
    \ces_7_6_io_outs_right[58] ,
    \ces_7_6_io_outs_right[57] ,
    \ces_7_6_io_outs_right[56] ,
    \ces_7_6_io_outs_right[55] ,
    \ces_7_6_io_outs_right[54] ,
    \ces_7_6_io_outs_right[53] ,
    \ces_7_6_io_outs_right[52] ,
    \ces_7_6_io_outs_right[51] ,
    \ces_7_6_io_outs_right[50] ,
    \ces_7_6_io_outs_right[49] ,
    \ces_7_6_io_outs_right[48] ,
    \ces_7_6_io_outs_right[47] ,
    \ces_7_6_io_outs_right[46] ,
    \ces_7_6_io_outs_right[45] ,
    \ces_7_6_io_outs_right[44] ,
    \ces_7_6_io_outs_right[43] ,
    \ces_7_6_io_outs_right[42] ,
    \ces_7_6_io_outs_right[41] ,
    \ces_7_6_io_outs_right[40] ,
    \ces_7_6_io_outs_right[39] ,
    \ces_7_6_io_outs_right[38] ,
    \ces_7_6_io_outs_right[37] ,
    \ces_7_6_io_outs_right[36] ,
    \ces_7_6_io_outs_right[35] ,
    \ces_7_6_io_outs_right[34] ,
    \ces_7_6_io_outs_right[33] ,
    \ces_7_6_io_outs_right[32] ,
    \ces_7_6_io_outs_right[31] ,
    \ces_7_6_io_outs_right[30] ,
    \ces_7_6_io_outs_right[29] ,
    \ces_7_6_io_outs_right[28] ,
    \ces_7_6_io_outs_right[27] ,
    \ces_7_6_io_outs_right[26] ,
    \ces_7_6_io_outs_right[25] ,
    \ces_7_6_io_outs_right[24] ,
    \ces_7_6_io_outs_right[23] ,
    \ces_7_6_io_outs_right[22] ,
    \ces_7_6_io_outs_right[21] ,
    \ces_7_6_io_outs_right[20] ,
    \ces_7_6_io_outs_right[19] ,
    \ces_7_6_io_outs_right[18] ,
    \ces_7_6_io_outs_right[17] ,
    \ces_7_6_io_outs_right[16] ,
    \ces_7_6_io_outs_right[15] ,
    \ces_7_6_io_outs_right[14] ,
    \ces_7_6_io_outs_right[13] ,
    \ces_7_6_io_outs_right[12] ,
    \ces_7_6_io_outs_right[11] ,
    \ces_7_6_io_outs_right[10] ,
    \ces_7_6_io_outs_right[9] ,
    \ces_7_6_io_outs_right[8] ,
    \ces_7_6_io_outs_right[7] ,
    \ces_7_6_io_outs_right[6] ,
    \ces_7_6_io_outs_right[5] ,
    \ces_7_6_io_outs_right[4] ,
    \ces_7_6_io_outs_right[3] ,
    \ces_7_6_io_outs_right[2] ,
    \ces_7_6_io_outs_right[1] ,
    \ces_7_6_io_outs_right[0] }),
    .io_outs_up({net4092,
    net4091,
    net4090,
    net4089,
    net4087,
    net4086,
    net4085,
    net4084,
    net4083,
    net4082,
    net4081,
    net4080,
    net4079,
    net4078,
    net4076,
    net4075,
    net4074,
    net4073,
    net4072,
    net4071,
    net4070,
    net4069,
    net4068,
    net4067,
    net4065,
    net4064,
    net4063,
    net4062,
    net4061,
    net4060,
    net4059,
    net4058,
    net4057,
    net4056,
    net4054,
    net4053,
    net4052,
    net4051,
    net4050,
    net4049,
    net4048,
    net4047,
    net4046,
    net4045,
    net4043,
    net4042,
    net4041,
    net4040,
    net4039,
    net4038,
    net4037,
    net4036,
    net4035,
    net4034,
    net4096,
    net4095,
    net4094,
    net4093,
    net4088,
    net4077,
    net4066,
    net4055,
    net4044,
    net4033}));
 Element ces_7_7 (.clock(clknet_3_7_0_clock),
    .io_lsbIns_1(ces_7_6_io_lsbOuts_1),
    .io_lsbIns_2(ces_7_6_io_lsbOuts_2),
    .io_lsbIns_3(ces_7_6_io_lsbOuts_3),
    .io_lsbIns_4(ces_7_6_io_lsbOuts_4),
    .io_lsbIns_5(ces_7_6_io_lsbOuts_5),
    .io_lsbIns_6(ces_7_6_io_lsbOuts_6),
    .io_lsbIns_7(ces_7_6_io_lsbOuts_7),
    .io_lsbOuts_0(ces_7_7_io_lsbOuts_0),
    .io_lsbOuts_1(ces_7_7_io_lsbOuts_1),
    .io_lsbOuts_2(ces_7_7_io_lsbOuts_2),
    .io_lsbOuts_3(ces_7_7_io_lsbOuts_3),
    .io_lsbOuts_4(ces_7_7_io_lsbOuts_4),
    .io_lsbOuts_5(ces_7_7_io_lsbOuts_5),
    .io_lsbOuts_6(ces_7_7_io_lsbOuts_6),
    .io_lsbOuts_7(ces_7_7_io_lsbOuts_7),
    .io_ins_down({net508,
    net507,
    net506,
    net505,
    net503,
    net502,
    net501,
    net500,
    net499,
    net498,
    net497,
    net496,
    net495,
    net494,
    net492,
    net491,
    net490,
    net489,
    net488,
    net487,
    net486,
    net485,
    net484,
    net483,
    net481,
    net480,
    net479,
    net478,
    net477,
    net476,
    net475,
    net474,
    net473,
    net472,
    net470,
    net469,
    net468,
    net467,
    net466,
    net465,
    net464,
    net463,
    net462,
    net461,
    net459,
    net458,
    net457,
    net456,
    net455,
    net454,
    net453,
    net452,
    net451,
    net450,
    net512,
    net511,
    net510,
    net509,
    net504,
    net493,
    net482,
    net471,
    net460,
    net449}),
    .io_ins_left({net1020,
    net1019,
    net1018,
    net1017,
    net1015,
    net1014,
    net1013,
    net1012,
    net1011,
    net1010,
    net1009,
    net1008,
    net1007,
    net1006,
    net1004,
    net1003,
    net1002,
    net1001,
    net1000,
    net999,
    net998,
    net997,
    net996,
    net995,
    net993,
    net992,
    net991,
    net990,
    net989,
    net988,
    net987,
    net986,
    net985,
    net984,
    net982,
    net981,
    net980,
    net979,
    net978,
    net977,
    net976,
    net975,
    net974,
    net973,
    net971,
    net970,
    net969,
    net968,
    net967,
    net966,
    net965,
    net964,
    net963,
    net962,
    net1024,
    net1023,
    net1022,
    net1021,
    net1016,
    net1005,
    net994,
    net983,
    net972,
    net961}),
    .io_ins_right({\ces_7_6_io_outs_right[63] ,
    \ces_7_6_io_outs_right[62] ,
    \ces_7_6_io_outs_right[61] ,
    \ces_7_6_io_outs_right[60] ,
    \ces_7_6_io_outs_right[59] ,
    \ces_7_6_io_outs_right[58] ,
    \ces_7_6_io_outs_right[57] ,
    \ces_7_6_io_outs_right[56] ,
    \ces_7_6_io_outs_right[55] ,
    \ces_7_6_io_outs_right[54] ,
    \ces_7_6_io_outs_right[53] ,
    \ces_7_6_io_outs_right[52] ,
    \ces_7_6_io_outs_right[51] ,
    \ces_7_6_io_outs_right[50] ,
    \ces_7_6_io_outs_right[49] ,
    \ces_7_6_io_outs_right[48] ,
    \ces_7_6_io_outs_right[47] ,
    \ces_7_6_io_outs_right[46] ,
    \ces_7_6_io_outs_right[45] ,
    \ces_7_6_io_outs_right[44] ,
    \ces_7_6_io_outs_right[43] ,
    \ces_7_6_io_outs_right[42] ,
    \ces_7_6_io_outs_right[41] ,
    \ces_7_6_io_outs_right[40] ,
    \ces_7_6_io_outs_right[39] ,
    \ces_7_6_io_outs_right[38] ,
    \ces_7_6_io_outs_right[37] ,
    \ces_7_6_io_outs_right[36] ,
    \ces_7_6_io_outs_right[35] ,
    \ces_7_6_io_outs_right[34] ,
    \ces_7_6_io_outs_right[33] ,
    \ces_7_6_io_outs_right[32] ,
    \ces_7_6_io_outs_right[31] ,
    \ces_7_6_io_outs_right[30] ,
    \ces_7_6_io_outs_right[29] ,
    \ces_7_6_io_outs_right[28] ,
    \ces_7_6_io_outs_right[27] ,
    \ces_7_6_io_outs_right[26] ,
    \ces_7_6_io_outs_right[25] ,
    \ces_7_6_io_outs_right[24] ,
    \ces_7_6_io_outs_right[23] ,
    \ces_7_6_io_outs_right[22] ,
    \ces_7_6_io_outs_right[21] ,
    \ces_7_6_io_outs_right[20] ,
    \ces_7_6_io_outs_right[19] ,
    \ces_7_6_io_outs_right[18] ,
    \ces_7_6_io_outs_right[17] ,
    \ces_7_6_io_outs_right[16] ,
    \ces_7_6_io_outs_right[15] ,
    \ces_7_6_io_outs_right[14] ,
    \ces_7_6_io_outs_right[13] ,
    \ces_7_6_io_outs_right[12] ,
    \ces_7_6_io_outs_right[11] ,
    \ces_7_6_io_outs_right[10] ,
    \ces_7_6_io_outs_right[9] ,
    \ces_7_6_io_outs_right[8] ,
    \ces_7_6_io_outs_right[7] ,
    \ces_7_6_io_outs_right[6] ,
    \ces_7_6_io_outs_right[5] ,
    \ces_7_6_io_outs_right[4] ,
    \ces_7_6_io_outs_right[3] ,
    \ces_7_6_io_outs_right[2] ,
    \ces_7_6_io_outs_right[1] ,
    \ces_7_6_io_outs_right[0] }),
    .io_ins_up({\ces_6_7_io_outs_up[63] ,
    \ces_6_7_io_outs_up[62] ,
    \ces_6_7_io_outs_up[61] ,
    \ces_6_7_io_outs_up[60] ,
    \ces_6_7_io_outs_up[59] ,
    \ces_6_7_io_outs_up[58] ,
    \ces_6_7_io_outs_up[57] ,
    \ces_6_7_io_outs_up[56] ,
    \ces_6_7_io_outs_up[55] ,
    \ces_6_7_io_outs_up[54] ,
    \ces_6_7_io_outs_up[53] ,
    \ces_6_7_io_outs_up[52] ,
    \ces_6_7_io_outs_up[51] ,
    \ces_6_7_io_outs_up[50] ,
    \ces_6_7_io_outs_up[49] ,
    \ces_6_7_io_outs_up[48] ,
    \ces_6_7_io_outs_up[47] ,
    \ces_6_7_io_outs_up[46] ,
    \ces_6_7_io_outs_up[45] ,
    \ces_6_7_io_outs_up[44] ,
    \ces_6_7_io_outs_up[43] ,
    \ces_6_7_io_outs_up[42] ,
    \ces_6_7_io_outs_up[41] ,
    \ces_6_7_io_outs_up[40] ,
    \ces_6_7_io_outs_up[39] ,
    \ces_6_7_io_outs_up[38] ,
    \ces_6_7_io_outs_up[37] ,
    \ces_6_7_io_outs_up[36] ,
    \ces_6_7_io_outs_up[35] ,
    \ces_6_7_io_outs_up[34] ,
    \ces_6_7_io_outs_up[33] ,
    \ces_6_7_io_outs_up[32] ,
    \ces_6_7_io_outs_up[31] ,
    \ces_6_7_io_outs_up[30] ,
    \ces_6_7_io_outs_up[29] ,
    \ces_6_7_io_outs_up[28] ,
    \ces_6_7_io_outs_up[27] ,
    \ces_6_7_io_outs_up[26] ,
    \ces_6_7_io_outs_up[25] ,
    \ces_6_7_io_outs_up[24] ,
    \ces_6_7_io_outs_up[23] ,
    \ces_6_7_io_outs_up[22] ,
    \ces_6_7_io_outs_up[21] ,
    \ces_6_7_io_outs_up[20] ,
    \ces_6_7_io_outs_up[19] ,
    \ces_6_7_io_outs_up[18] ,
    \ces_6_7_io_outs_up[17] ,
    \ces_6_7_io_outs_up[16] ,
    \ces_6_7_io_outs_up[15] ,
    \ces_6_7_io_outs_up[14] ,
    \ces_6_7_io_outs_up[13] ,
    \ces_6_7_io_outs_up[12] ,
    \ces_6_7_io_outs_up[11] ,
    \ces_6_7_io_outs_up[10] ,
    \ces_6_7_io_outs_up[9] ,
    \ces_6_7_io_outs_up[8] ,
    \ces_6_7_io_outs_up[7] ,
    \ces_6_7_io_outs_up[6] ,
    \ces_6_7_io_outs_up[5] ,
    \ces_6_7_io_outs_up[4] ,
    \ces_6_7_io_outs_up[3] ,
    \ces_6_7_io_outs_up[2] ,
    \ces_6_7_io_outs_up[1] ,
    \ces_6_7_io_outs_up[0] }),
    .io_outs_down({\ces_6_7_io_ins_down[63] ,
    \ces_6_7_io_ins_down[62] ,
    \ces_6_7_io_ins_down[61] ,
    \ces_6_7_io_ins_down[60] ,
    \ces_6_7_io_ins_down[59] ,
    \ces_6_7_io_ins_down[58] ,
    \ces_6_7_io_ins_down[57] ,
    \ces_6_7_io_ins_down[56] ,
    \ces_6_7_io_ins_down[55] ,
    \ces_6_7_io_ins_down[54] ,
    \ces_6_7_io_ins_down[53] ,
    \ces_6_7_io_ins_down[52] ,
    \ces_6_7_io_ins_down[51] ,
    \ces_6_7_io_ins_down[50] ,
    \ces_6_7_io_ins_down[49] ,
    \ces_6_7_io_ins_down[48] ,
    \ces_6_7_io_ins_down[47] ,
    \ces_6_7_io_ins_down[46] ,
    \ces_6_7_io_ins_down[45] ,
    \ces_6_7_io_ins_down[44] ,
    \ces_6_7_io_ins_down[43] ,
    \ces_6_7_io_ins_down[42] ,
    \ces_6_7_io_ins_down[41] ,
    \ces_6_7_io_ins_down[40] ,
    \ces_6_7_io_ins_down[39] ,
    \ces_6_7_io_ins_down[38] ,
    \ces_6_7_io_ins_down[37] ,
    \ces_6_7_io_ins_down[36] ,
    \ces_6_7_io_ins_down[35] ,
    \ces_6_7_io_ins_down[34] ,
    \ces_6_7_io_ins_down[33] ,
    \ces_6_7_io_ins_down[32] ,
    \ces_6_7_io_ins_down[31] ,
    \ces_6_7_io_ins_down[30] ,
    \ces_6_7_io_ins_down[29] ,
    \ces_6_7_io_ins_down[28] ,
    \ces_6_7_io_ins_down[27] ,
    \ces_6_7_io_ins_down[26] ,
    \ces_6_7_io_ins_down[25] ,
    \ces_6_7_io_ins_down[24] ,
    \ces_6_7_io_ins_down[23] ,
    \ces_6_7_io_ins_down[22] ,
    \ces_6_7_io_ins_down[21] ,
    \ces_6_7_io_ins_down[20] ,
    \ces_6_7_io_ins_down[19] ,
    \ces_6_7_io_ins_down[18] ,
    \ces_6_7_io_ins_down[17] ,
    \ces_6_7_io_ins_down[16] ,
    \ces_6_7_io_ins_down[15] ,
    \ces_6_7_io_ins_down[14] ,
    \ces_6_7_io_ins_down[13] ,
    \ces_6_7_io_ins_down[12] ,
    \ces_6_7_io_ins_down[11] ,
    \ces_6_7_io_ins_down[10] ,
    \ces_6_7_io_ins_down[9] ,
    \ces_6_7_io_ins_down[8] ,
    \ces_6_7_io_ins_down[7] ,
    \ces_6_7_io_ins_down[6] ,
    \ces_6_7_io_ins_down[5] ,
    \ces_6_7_io_ins_down[4] ,
    \ces_6_7_io_ins_down[3] ,
    \ces_6_7_io_ins_down[2] ,
    \ces_6_7_io_ins_down[1] ,
    \ces_6_7_io_ins_down[0] }),
    .io_outs_left({\ces_7_6_io_ins_left[63] ,
    \ces_7_6_io_ins_left[62] ,
    \ces_7_6_io_ins_left[61] ,
    \ces_7_6_io_ins_left[60] ,
    \ces_7_6_io_ins_left[59] ,
    \ces_7_6_io_ins_left[58] ,
    \ces_7_6_io_ins_left[57] ,
    \ces_7_6_io_ins_left[56] ,
    \ces_7_6_io_ins_left[55] ,
    \ces_7_6_io_ins_left[54] ,
    \ces_7_6_io_ins_left[53] ,
    \ces_7_6_io_ins_left[52] ,
    \ces_7_6_io_ins_left[51] ,
    \ces_7_6_io_ins_left[50] ,
    \ces_7_6_io_ins_left[49] ,
    \ces_7_6_io_ins_left[48] ,
    \ces_7_6_io_ins_left[47] ,
    \ces_7_6_io_ins_left[46] ,
    \ces_7_6_io_ins_left[45] ,
    \ces_7_6_io_ins_left[44] ,
    \ces_7_6_io_ins_left[43] ,
    \ces_7_6_io_ins_left[42] ,
    \ces_7_6_io_ins_left[41] ,
    \ces_7_6_io_ins_left[40] ,
    \ces_7_6_io_ins_left[39] ,
    \ces_7_6_io_ins_left[38] ,
    \ces_7_6_io_ins_left[37] ,
    \ces_7_6_io_ins_left[36] ,
    \ces_7_6_io_ins_left[35] ,
    \ces_7_6_io_ins_left[34] ,
    \ces_7_6_io_ins_left[33] ,
    \ces_7_6_io_ins_left[32] ,
    \ces_7_6_io_ins_left[31] ,
    \ces_7_6_io_ins_left[30] ,
    \ces_7_6_io_ins_left[29] ,
    \ces_7_6_io_ins_left[28] ,
    \ces_7_6_io_ins_left[27] ,
    \ces_7_6_io_ins_left[26] ,
    \ces_7_6_io_ins_left[25] ,
    \ces_7_6_io_ins_left[24] ,
    \ces_7_6_io_ins_left[23] ,
    \ces_7_6_io_ins_left[22] ,
    \ces_7_6_io_ins_left[21] ,
    \ces_7_6_io_ins_left[20] ,
    \ces_7_6_io_ins_left[19] ,
    \ces_7_6_io_ins_left[18] ,
    \ces_7_6_io_ins_left[17] ,
    \ces_7_6_io_ins_left[16] ,
    \ces_7_6_io_ins_left[15] ,
    \ces_7_6_io_ins_left[14] ,
    \ces_7_6_io_ins_left[13] ,
    \ces_7_6_io_ins_left[12] ,
    \ces_7_6_io_ins_left[11] ,
    \ces_7_6_io_ins_left[10] ,
    \ces_7_6_io_ins_left[9] ,
    \ces_7_6_io_ins_left[8] ,
    \ces_7_6_io_ins_left[7] ,
    \ces_7_6_io_ins_left[6] ,
    \ces_7_6_io_ins_left[5] ,
    \ces_7_6_io_ins_left[4] ,
    \ces_7_6_io_ins_left[3] ,
    \ces_7_6_io_ins_left[2] ,
    \ces_7_6_io_ins_left[1] ,
    \ces_7_6_io_ins_left[0] }),
    .io_outs_right({net3644,
    net3643,
    net3642,
    net3641,
    net3639,
    net3638,
    net3637,
    net3636,
    net3635,
    net3634,
    net3633,
    net3632,
    net3631,
    net3630,
    net3628,
    net3627,
    net3626,
    net3625,
    net3624,
    net3623,
    net3622,
    net3621,
    net3620,
    net3619,
    net3617,
    net3616,
    net3615,
    net3614,
    net3613,
    net3612,
    net3611,
    net3610,
    net3609,
    net3608,
    net3606,
    net3605,
    net3604,
    net3603,
    net3602,
    net3601,
    net3600,
    net3599,
    net3598,
    net3597,
    net3595,
    net3594,
    net3593,
    net3592,
    net3591,
    net3590,
    net3589,
    net3588,
    net3587,
    net3586,
    net3648,
    net3647,
    net3646,
    net3645,
    net3640,
    net3629,
    net3618,
    net3607,
    net3596,
    net3585}),
    .io_outs_up({net4156,
    net4155,
    net4154,
    net4153,
    net4151,
    net4150,
    net4149,
    net4148,
    net4147,
    net4146,
    net4145,
    net4144,
    net4143,
    net4142,
    net4140,
    net4139,
    net4138,
    net4137,
    net4136,
    net4135,
    net4134,
    net4133,
    net4132,
    net4131,
    net4129,
    net4128,
    net4127,
    net4126,
    net4125,
    net4124,
    net4123,
    net4122,
    net4121,
    net4120,
    net4118,
    net4117,
    net4116,
    net4115,
    net4114,
    net4113,
    net4112,
    net4111,
    net4110,
    net4109,
    net4107,
    net4106,
    net4105,
    net4104,
    net4103,
    net4102,
    net4101,
    net4100,
    net4099,
    net4098,
    net4160,
    net4159,
    net4158,
    net4157,
    net4152,
    net4141,
    net4130,
    net4119,
    net4108,
    net4097}));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_0$_DFF_P_  (.CLK(clknet_3_0_0_clock_regs),
    .D(ces_0_7_io_lsbOuts_0),
    .QN(_001_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_1$_DFF_P_  (.CLK(clknet_3_2_0_clock_regs),
    .D(ces_0_7_io_lsbOuts_1),
    .QN(_000_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_10$_DFF_P_  (.CLK(clknet_3_2_0_clock_regs),
    .D(ces_1_7_io_lsbOuts_2),
    .QN(_010_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_11$_DFF_P_  (.CLK(clknet_3_2_0_clock_regs),
    .D(ces_1_7_io_lsbOuts_3),
    .QN(_011_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_12$_DFF_P_  (.CLK(clknet_3_0_0_clock_regs),
    .D(ces_1_7_io_lsbOuts_4),
    .QN(_012_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_13$_DFF_P_  (.CLK(clknet_3_2_0_clock_regs),
    .D(ces_1_7_io_lsbOuts_5),
    .QN(_013_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_14$_DFF_P_  (.CLK(clknet_3_0_0_clock_regs),
    .D(ces_1_7_io_lsbOuts_6),
    .QN(_014_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_15$_DFF_P_  (.CLK(clknet_3_0_0_clock_regs),
    .D(ces_1_7_io_lsbOuts_7),
    .QN(_015_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_16$_DFF_P_  (.CLK(clknet_3_1_0_clock_regs),
    .D(ces_2_7_io_lsbOuts_0),
    .QN(_016_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_17$_DFF_P_  (.CLK(clknet_3_3_0_clock_regs),
    .D(ces_2_7_io_lsbOuts_1),
    .QN(_017_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_18$_DFF_P_  (.CLK(clknet_3_3_0_clock_regs),
    .D(ces_2_7_io_lsbOuts_2),
    .QN(_018_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_19$_DFF_P_  (.CLK(clknet_3_1_0_clock_regs),
    .D(ces_2_7_io_lsbOuts_3),
    .QN(_019_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_2$_DFF_P_  (.CLK(clknet_3_0_0_clock_regs),
    .D(ces_0_7_io_lsbOuts_2),
    .QN(_002_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_20$_DFF_P_  (.CLK(clknet_3_1_0_clock_regs),
    .D(ces_2_7_io_lsbOuts_4),
    .QN(_020_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_21$_DFF_P_  (.CLK(clknet_3_3_0_clock_regs),
    .D(ces_2_7_io_lsbOuts_5),
    .QN(_021_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_22$_DFF_P_  (.CLK(clknet_3_3_0_clock_regs),
    .D(ces_2_7_io_lsbOuts_6),
    .QN(_022_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_23$_DFF_P_  (.CLK(clknet_3_3_0_clock_regs),
    .D(ces_2_7_io_lsbOuts_7),
    .QN(_023_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_24$_DFF_P_  (.CLK(clknet_3_1_0_clock_regs),
    .D(ces_3_7_io_lsbOuts_0),
    .QN(_024_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_25$_DFF_P_  (.CLK(clknet_3_1_0_clock_regs),
    .D(ces_3_7_io_lsbOuts_1),
    .QN(_025_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_26$_DFF_P_  (.CLK(clknet_3_3_0_clock_regs),
    .D(ces_3_7_io_lsbOuts_2),
    .QN(_026_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_27$_DFF_P_  (.CLK(clknet_3_1_0_clock_regs),
    .D(ces_3_7_io_lsbOuts_3),
    .QN(_027_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_28$_DFF_P_  (.CLK(clknet_3_3_0_clock_regs),
    .D(ces_3_7_io_lsbOuts_4),
    .QN(_028_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_29$_DFF_P_  (.CLK(clknet_3_1_0_clock_regs),
    .D(ces_3_7_io_lsbOuts_5),
    .QN(_029_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_3$_DFF_P_  (.CLK(clknet_3_2_0_clock_regs),
    .D(ces_0_7_io_lsbOuts_3),
    .QN(_003_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_30$_DFF_P_  (.CLK(clknet_3_1_0_clock_regs),
    .D(ces_3_7_io_lsbOuts_6),
    .QN(_030_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_31$_DFF_P_  (.CLK(clknet_3_3_0_clock_regs),
    .D(ces_3_7_io_lsbOuts_7),
    .QN(_031_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_32$_DFF_P_  (.CLK(clknet_3_7_0_clock_regs),
    .D(ces_4_7_io_lsbOuts_0),
    .QN(_032_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_33$_DFF_P_  (.CLK(clknet_3_6_0_clock_regs),
    .D(ces_4_7_io_lsbOuts_1),
    .QN(_033_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_34$_DFF_P_  (.CLK(clknet_3_6_0_clock_regs),
    .D(ces_4_7_io_lsbOuts_2),
    .QN(_034_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_35$_DFF_P_  (.CLK(clknet_3_6_0_clock_regs),
    .D(ces_4_7_io_lsbOuts_3),
    .QN(_035_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_36$_DFF_P_  (.CLK(clknet_3_6_0_clock_regs),
    .D(ces_4_7_io_lsbOuts_4),
    .QN(_036_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_37$_DFF_P_  (.CLK(clknet_3_7_0_clock_regs),
    .D(ces_4_7_io_lsbOuts_5),
    .QN(_037_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_38$_DFF_P_  (.CLK(clknet_3_6_0_clock_regs),
    .D(ces_4_7_io_lsbOuts_6),
    .QN(_038_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_39$_DFF_P_  (.CLK(clknet_3_6_0_clock_regs),
    .D(ces_4_7_io_lsbOuts_7),
    .QN(_039_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_4$_DFF_P_  (.CLK(clknet_3_0_0_clock_regs),
    .D(ces_0_7_io_lsbOuts_4),
    .QN(_004_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_40$_DFF_P_  (.CLK(clknet_3_7_0_clock_regs),
    .D(ces_5_7_io_lsbOuts_0),
    .QN(_040_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_41$_DFF_P_  (.CLK(clknet_3_6_0_clock_regs),
    .D(ces_5_7_io_lsbOuts_1),
    .QN(_041_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_42$_DFF_P_  (.CLK(clknet_3_7_0_clock_regs),
    .D(ces_5_7_io_lsbOuts_2),
    .QN(_042_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_43$_DFF_P_  (.CLK(clknet_3_6_0_clock_regs),
    .D(ces_5_7_io_lsbOuts_3),
    .QN(_043_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_44$_DFF_P_  (.CLK(clknet_3_6_0_clock_regs),
    .D(ces_5_7_io_lsbOuts_4),
    .QN(_044_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_45$_DFF_P_  (.CLK(clknet_3_7_0_clock_regs),
    .D(ces_5_7_io_lsbOuts_5),
    .QN(_045_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_46$_DFF_P_  (.CLK(clknet_3_7_0_clock_regs),
    .D(ces_5_7_io_lsbOuts_6),
    .QN(_046_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_47$_DFF_P_  (.CLK(clknet_3_7_0_clock_regs),
    .D(ces_5_7_io_lsbOuts_7),
    .QN(_047_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_48$_DFF_P_  (.CLK(clknet_3_4_0_clock_regs),
    .D(ces_6_7_io_lsbOuts_0),
    .QN(_048_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_49$_DFF_P_  (.CLK(clknet_3_4_0_clock_regs),
    .D(ces_6_7_io_lsbOuts_1),
    .QN(_049_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_5$_DFF_P_  (.CLK(clknet_3_2_0_clock_regs),
    .D(ces_0_7_io_lsbOuts_5),
    .QN(_005_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_50$_DFF_P_  (.CLK(clknet_3_5_0_clock_regs),
    .D(ces_6_7_io_lsbOuts_2),
    .QN(_050_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_51$_DFF_P_  (.CLK(clknet_3_4_0_clock_regs),
    .D(ces_6_7_io_lsbOuts_3),
    .QN(_051_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_52$_DFF_P_  (.CLK(clknet_3_4_0_clock_regs),
    .D(ces_6_7_io_lsbOuts_4),
    .QN(_052_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_53$_DFF_P_  (.CLK(clknet_3_5_0_clock_regs),
    .D(ces_6_7_io_lsbOuts_5),
    .QN(_053_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_54$_DFF_P_  (.CLK(clknet_3_5_0_clock_regs),
    .D(ces_6_7_io_lsbOuts_6),
    .QN(_054_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_55$_DFF_P_  (.CLK(clknet_3_4_0_clock_regs),
    .D(ces_6_7_io_lsbOuts_7),
    .QN(_055_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_56$_DFF_P_  (.CLK(clknet_3_5_0_clock_regs),
    .D(ces_7_7_io_lsbOuts_0),
    .QN(_056_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_57$_DFF_P_  (.CLK(clknet_3_4_0_clock_regs),
    .D(ces_7_7_io_lsbOuts_1),
    .QN(_057_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_58$_DFF_P_  (.CLK(clknet_3_5_0_clock_regs),
    .D(ces_7_7_io_lsbOuts_2),
    .QN(_058_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_59$_DFF_P_  (.CLK(clknet_3_5_0_clock_regs),
    .D(ces_7_7_io_lsbOuts_3),
    .QN(_059_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_6$_DFF_P_  (.CLK(clknet_3_0_0_clock_regs),
    .D(ces_0_7_io_lsbOuts_6),
    .QN(_006_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_60$_DFF_P_  (.CLK(clknet_3_5_0_clock_regs),
    .D(ces_7_7_io_lsbOuts_4),
    .QN(_060_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_61$_DFF_P_  (.CLK(clknet_3_5_0_clock_regs),
    .D(ces_7_7_io_lsbOuts_5),
    .QN(_061_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_62$_DFF_P_  (.CLK(clknet_3_4_0_clock_regs),
    .D(ces_7_7_io_lsbOuts_6),
    .QN(_062_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_63$_DFF_P_  (.CLK(clknet_3_5_0_clock_regs),
    .D(ces_7_7_io_lsbOuts_7),
    .QN(_063_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_7$_DFF_P_  (.CLK(clknet_3_0_0_clock_regs),
    .D(ces_0_7_io_lsbOuts_7),
    .QN(_007_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_8$_DFF_P_  (.CLK(clknet_3_2_0_clock_regs),
    .D(ces_1_7_io_lsbOuts_0),
    .QN(_008_));
 DFFHQNx2_ASAP7_75t_R \io_lsbs_9$_DFF_P_  (.CLK(clknet_3_0_0_clock_regs),
    .D(ces_1_7_io_lsbOuts_1),
    .QN(_009_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_354_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_355_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_356_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_357_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_358_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_359_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_360_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_361_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_362_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_363_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_364_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_365_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_530_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_531_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_532_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_533_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_534_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_535_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_536_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_537_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_538_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_539_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_540_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_541_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_706_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_707_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_708_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_709_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_710_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_711_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_712_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_713_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_714_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_715_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_716_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_717_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_882_Right_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_883_Right_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_884_Right_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_885_Right_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_886_Right_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_887_Right_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_888_Right_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_889_Right_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_890_Right_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_891_Right_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_892_Right_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_893_Right_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1058_Right_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1059_Right_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1060_Right_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1061_Right_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1062_Right_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1063_Right_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1064_Right_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1065_Right_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1066_Right_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1067_Right_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1068_Right_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1069_Right_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1234_Right_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1235_Right_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1236_Right_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1237_Right_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1238_Right_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1239_Right_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1240_Right_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1241_Right_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1242_Right_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1243_Right_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1244_Right_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1245_Right_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1410_Right_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1411_Right_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1412_Right_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1413_Right_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1414_Right_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1415_Right_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1416_Right_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1417_Right_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1418_Right_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1419_Right_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1420_Right_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1421_Right_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1422_Right_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1423_Right_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_9_Right_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_9_Right_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_9_Right_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_9_Right_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_9_Right_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_9_Right_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_9_Right_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_9_Right_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_9_Right_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_9_Right_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_9_Right_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_9_Right_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_9_Right_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_9_Right_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_9_Right_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_9_Right_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_9_Right_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_9_Right_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_9_Right_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_9_Right_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_9_Right_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_9_Right_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_9_Right_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_9_Right_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_9_Right_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_9_Right_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_9_Right_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_9_Right_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_9_Right_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_9_Right_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_9_Right_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_9_Right_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_9_Right_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_9_Right_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_9_Right_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_9_Right_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_9_Right_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_9_Right_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_9_Right_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_9_Right_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_9_Right_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_9_Right_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_9_Right_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_9_Right_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_9_Right_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_9_Right_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_9_Right_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_9_Right_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_9_Right_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_9_Right_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_9_Right_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_9_Right_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_9_Right_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_9_Right_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_9_Right_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_9_Right_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_9_Right_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_9_Right_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_9_Right_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_9_Right_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_9_Right_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_9_Right_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_9_Right_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_9_Right_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_9_Right_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_9_Right_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_9_Right_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_9_Right_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_9_Right_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_9_Right_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_9_Right_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_9_Right_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_9_Right_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_9_Right_185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_9_Right_186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_9_Right_187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_9_Right_188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_9_Right_189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_9_Right_190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_9_Right_191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_9_Right_192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_9_Right_193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_9_Right_194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_9_Right_195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_9_Right_196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_9_Right_197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_9_Right_198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_9_Right_199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_9_Right_200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_9_Right_201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_9_Right_202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_9_Right_203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_9_Right_204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_9_Right_205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_9_Right_206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_9_Right_207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_9_Right_208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_9_Right_209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_9_Right_210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_9_Right_211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_9_Right_212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_9_Right_213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_9_Right_214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_9_Right_215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_9_Right_216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_9_Right_217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_9_Right_218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_9_Right_219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_9_Right_220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_9_Right_221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_9_Right_222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_9_Right_223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_9_Right_224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_9_Right_225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_9_Right_226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_9_Right_227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_9_Right_228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_9_Right_229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_9_Right_230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_9_Right_231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_9_Right_232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_9_Right_233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_9_Right_234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_9_Right_235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_9_Right_236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_9_Right_237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_9_Right_238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_9_Right_239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_9_Right_240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_9_Right_241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_9_Right_242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_9_Right_243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_9_Right_244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_9_Right_245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_9_Right_246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_9_Right_247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_9_Right_248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_9_Right_249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_9_Right_250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_9_Right_251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_9_Right_252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_9_Right_253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_9_Right_254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_9_Right_255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_9_Right_256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_9_Right_257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_9_Right_258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_9_Right_259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_9_Right_260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_9_Right_261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_9_Right_262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_9_Right_263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_9_Right_264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_9_Right_265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_9_Right_266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_9_Right_267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_9_Right_268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_9_Right_269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_9_Right_270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_9_Right_271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_9_Right_272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_9_Right_273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_9_Right_274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_9_Right_275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_9_Right_276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_9_Right_277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_9_Right_278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_9_Right_279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_9_Right_280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_9_Right_281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_9_Right_282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_9_Right_283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_9_Right_284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_9_Right_285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_9_Right_286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_9_Right_287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_9_Right_288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_9_Right_289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_9_Right_290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_9_Right_291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_9_Right_292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_9_Right_293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_9_Right_294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_9_Right_295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_9_Right_296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_9_Right_297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_9_Right_298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_9_Right_299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_9_Right_300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_9_Right_301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_9_Right_302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_9_Right_303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_9_Right_304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_9_Right_305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_9_Right_306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_9_Right_307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_9_Right_308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_9_Right_309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_9_Right_310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_9_Right_311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_9_Right_312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_9_Right_313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_9_Right_314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_9_Right_315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_9_Right_316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_9_Right_317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_9_Right_318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_9_Right_319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_9_Right_320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_9_Right_321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_9_Right_322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_9_Right_323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_9_Right_324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_9_Right_325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_9_Right_326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_9_Right_327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_9_Right_328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_9_Right_329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_9_Right_330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_9_Right_331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_9_Right_332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_9_Right_333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_9_Right_334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_9_Right_335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_9_Right_336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_9_Right_337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_9_Right_338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_9_Right_339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_9_Right_340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_9_Right_341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_9_Right_342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_9_Right_343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_9_Right_344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_9_Right_345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_9_Right_346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_9_Right_347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_9_Right_348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_9_Right_349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_9_Right_350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_9_Right_351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_9_Right_352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_9_Right_353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_9_Right_354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_9_Right_355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_9_Right_356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_9_Right_357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_9_Right_358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_9_Right_359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_9_Right_360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_9_Right_361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_9_Right_362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_9_Right_363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_9_Right_364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_9_Right_365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_9_Right_366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_9_Right_367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_9_Right_368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_9_Right_369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_9_Right_370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_9_Right_371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_9_Right_372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_9_Right_373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_9_Right_374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_9_Right_375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_9_Right_376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_9_Right_377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_9_Right_378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_9_Right_379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_9_Right_380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_295_9_Right_381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_296_9_Right_382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_297_9_Right_383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_298_9_Right_384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_299_9_Right_385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_300_9_Right_386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_301_9_Right_387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_302_9_Right_388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_303_9_Right_389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_304_9_Right_390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_305_9_Right_391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_306_9_Right_392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_307_9_Right_393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_308_9_Right_394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_309_9_Right_395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_310_9_Right_396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_311_9_Right_397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_312_9_Right_398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_313_9_Right_399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_314_9_Right_400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_315_9_Right_401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_316_9_Right_402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_317_9_Right_403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_318_9_Right_404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_319_9_Right_405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_320_9_Right_406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_321_9_Right_407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_322_9_Right_408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_323_9_Right_409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_324_9_Right_410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_325_9_Right_411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_326_9_Right_412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_327_9_Right_413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_328_9_Right_414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_329_9_Right_415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_330_9_Right_416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_331_9_Right_417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_332_9_Right_418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_333_9_Right_419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_334_9_Right_420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_335_9_Right_421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_336_9_Right_422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_337_9_Right_423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_338_9_Right_424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_339_9_Right_425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_340_9_Right_426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_341_9_Right_427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_342_9_Right_428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_343_9_Right_429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_344_9_Right_430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_345_9_Right_431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_346_9_Right_432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_347_9_Right_433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_348_9_Right_434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_349_9_Right_435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_350_9_Right_436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_351_9_Right_437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_352_9_Right_438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_353_9_Right_439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_366_9_Right_440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_367_9_Right_441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_368_9_Right_442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_369_9_Right_443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_370_9_Right_444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_371_9_Right_445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_372_9_Right_446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_373_9_Right_447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_374_9_Right_448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_375_9_Right_449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_376_9_Right_450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_377_9_Right_451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_378_9_Right_452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_379_9_Right_453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_380_9_Right_454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_381_9_Right_455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_382_9_Right_456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_383_9_Right_457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_384_9_Right_458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_385_9_Right_459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_386_9_Right_460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_387_9_Right_461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_388_9_Right_462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_389_9_Right_463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_390_9_Right_464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_391_9_Right_465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_392_9_Right_466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_393_9_Right_467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_394_9_Right_468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_395_9_Right_469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_396_9_Right_470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_397_9_Right_471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_398_9_Right_472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_399_9_Right_473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_400_9_Right_474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_401_9_Right_475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_402_9_Right_476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_403_9_Right_477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_404_9_Right_478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_405_9_Right_479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_406_9_Right_480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_407_9_Right_481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_408_9_Right_482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_409_9_Right_483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_410_9_Right_484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_411_9_Right_485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_412_9_Right_486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_413_9_Right_487 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_414_9_Right_488 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_415_9_Right_489 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_416_9_Right_490 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_417_9_Right_491 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_418_9_Right_492 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_419_9_Right_493 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_420_9_Right_494 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_421_9_Right_495 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_422_9_Right_496 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_423_9_Right_497 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_424_9_Right_498 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_425_9_Right_499 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_426_9_Right_500 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_427_9_Right_501 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_428_9_Right_502 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_429_9_Right_503 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_430_9_Right_504 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_431_9_Right_505 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_432_9_Right_506 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_433_9_Right_507 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_434_9_Right_508 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_435_9_Right_509 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_436_9_Right_510 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_437_9_Right_511 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_438_9_Right_512 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_439_9_Right_513 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_440_9_Right_514 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_441_9_Right_515 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_442_9_Right_516 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_443_9_Right_517 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_444_9_Right_518 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_445_9_Right_519 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_446_9_Right_520 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_447_9_Right_521 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_448_9_Right_522 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_449_9_Right_523 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_450_9_Right_524 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_451_9_Right_525 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_452_9_Right_526 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_453_9_Right_527 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_454_9_Right_528 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_455_9_Right_529 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_456_9_Right_530 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_457_9_Right_531 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_458_9_Right_532 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_459_9_Right_533 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_460_9_Right_534 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_461_9_Right_535 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_462_9_Right_536 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_463_9_Right_537 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_464_9_Right_538 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_465_9_Right_539 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_466_9_Right_540 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_467_9_Right_541 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_468_9_Right_542 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_469_9_Right_543 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_470_9_Right_544 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_471_9_Right_545 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_472_9_Right_546 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_473_9_Right_547 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_474_9_Right_548 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_475_9_Right_549 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_476_9_Right_550 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_477_9_Right_551 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_478_9_Right_552 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_479_9_Right_553 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_480_9_Right_554 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_481_9_Right_555 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_482_9_Right_556 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_483_9_Right_557 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_484_9_Right_558 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_485_9_Right_559 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_486_9_Right_560 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_487_9_Right_561 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_488_9_Right_562 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_489_9_Right_563 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_490_9_Right_564 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_491_9_Right_565 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_492_9_Right_566 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_493_9_Right_567 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_494_9_Right_568 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_495_9_Right_569 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_496_9_Right_570 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_497_9_Right_571 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_498_9_Right_572 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_499_9_Right_573 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_500_9_Right_574 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_501_9_Right_575 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_502_9_Right_576 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_503_9_Right_577 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_504_9_Right_578 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_505_9_Right_579 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_506_9_Right_580 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_507_9_Right_581 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_508_9_Right_582 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_509_9_Right_583 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_510_9_Right_584 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_511_9_Right_585 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_512_9_Right_586 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_513_9_Right_587 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_514_9_Right_588 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_515_9_Right_589 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_516_9_Right_590 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_517_9_Right_591 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_518_9_Right_592 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_519_9_Right_593 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_520_9_Right_594 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_521_9_Right_595 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_522_9_Right_596 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_523_9_Right_597 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_524_9_Right_598 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_525_9_Right_599 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_526_9_Right_600 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_527_9_Right_601 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_528_9_Right_602 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_529_9_Right_603 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_542_9_Right_604 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_543_9_Right_605 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_544_9_Right_606 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_545_9_Right_607 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_546_9_Right_608 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_547_9_Right_609 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_548_9_Right_610 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_549_9_Right_611 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_550_9_Right_612 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_551_9_Right_613 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_552_9_Right_614 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_553_9_Right_615 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_554_9_Right_616 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_555_9_Right_617 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_556_9_Right_618 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_557_9_Right_619 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_558_9_Right_620 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_559_9_Right_621 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_560_9_Right_622 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_561_9_Right_623 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_562_9_Right_624 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_563_9_Right_625 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_564_9_Right_626 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_565_9_Right_627 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_566_9_Right_628 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_567_9_Right_629 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_568_9_Right_630 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_569_9_Right_631 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_570_9_Right_632 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_571_9_Right_633 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_572_9_Right_634 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_573_9_Right_635 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_574_9_Right_636 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_575_9_Right_637 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_576_9_Right_638 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_577_9_Right_639 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_578_9_Right_640 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_579_9_Right_641 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_580_9_Right_642 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_581_9_Right_643 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_582_9_Right_644 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_583_9_Right_645 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_584_9_Right_646 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_585_9_Right_647 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_586_9_Right_648 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_587_9_Right_649 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_588_9_Right_650 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_589_9_Right_651 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_590_9_Right_652 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_591_9_Right_653 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_592_9_Right_654 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_593_9_Right_655 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_594_9_Right_656 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_595_9_Right_657 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_596_9_Right_658 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_597_9_Right_659 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_598_9_Right_660 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_599_9_Right_661 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_600_9_Right_662 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_601_9_Right_663 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_602_9_Right_664 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_603_9_Right_665 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_604_9_Right_666 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_605_9_Right_667 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_606_9_Right_668 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_607_9_Right_669 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_608_9_Right_670 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_609_9_Right_671 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_610_9_Right_672 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_611_9_Right_673 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_612_9_Right_674 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_613_9_Right_675 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_614_9_Right_676 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_615_9_Right_677 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_616_9_Right_678 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_617_9_Right_679 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_618_9_Right_680 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_619_9_Right_681 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_620_9_Right_682 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_621_9_Right_683 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_622_9_Right_684 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_623_9_Right_685 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_624_9_Right_686 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_625_9_Right_687 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_626_9_Right_688 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_627_9_Right_689 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_628_9_Right_690 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_629_9_Right_691 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_630_9_Right_692 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_631_9_Right_693 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_632_9_Right_694 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_633_9_Right_695 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_634_9_Right_696 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_635_9_Right_697 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_636_9_Right_698 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_637_9_Right_699 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_638_9_Right_700 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_639_9_Right_701 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_640_9_Right_702 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_641_9_Right_703 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_642_9_Right_704 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_643_9_Right_705 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_644_9_Right_706 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_645_9_Right_707 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_646_9_Right_708 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_647_9_Right_709 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_648_9_Right_710 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_649_9_Right_711 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_650_9_Right_712 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_651_9_Right_713 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_652_9_Right_714 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_653_9_Right_715 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_654_9_Right_716 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_655_9_Right_717 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_656_9_Right_718 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_657_9_Right_719 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_658_9_Right_720 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_659_9_Right_721 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_660_9_Right_722 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_661_9_Right_723 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_662_9_Right_724 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_663_9_Right_725 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_664_9_Right_726 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_665_9_Right_727 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_666_9_Right_728 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_667_9_Right_729 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_668_9_Right_730 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_669_9_Right_731 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_670_9_Right_732 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_671_9_Right_733 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_672_9_Right_734 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_673_9_Right_735 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_674_9_Right_736 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_675_9_Right_737 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_676_9_Right_738 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_677_9_Right_739 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_678_9_Right_740 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_679_9_Right_741 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_680_9_Right_742 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_681_9_Right_743 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_682_9_Right_744 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_683_9_Right_745 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_684_9_Right_746 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_685_9_Right_747 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_686_9_Right_748 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_687_9_Right_749 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_688_9_Right_750 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_689_9_Right_751 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_690_9_Right_752 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_691_9_Right_753 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_692_9_Right_754 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_693_9_Right_755 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_694_9_Right_756 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_695_9_Right_757 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_696_9_Right_758 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_697_9_Right_759 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_698_9_Right_760 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_699_9_Right_761 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_700_9_Right_762 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_701_9_Right_763 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_702_9_Right_764 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_703_9_Right_765 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_704_9_Right_766 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_705_9_Right_767 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_718_9_Right_768 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_719_9_Right_769 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_720_9_Right_770 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_721_9_Right_771 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_722_9_Right_772 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_723_9_Right_773 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_724_9_Right_774 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_725_9_Right_775 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_726_9_Right_776 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_727_9_Right_777 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_728_9_Right_778 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_729_9_Right_779 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_730_9_Right_780 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_731_9_Right_781 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_732_9_Right_782 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_733_9_Right_783 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_734_9_Right_784 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_735_9_Right_785 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_736_9_Right_786 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_737_9_Right_787 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_738_9_Right_788 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_739_9_Right_789 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_740_9_Right_790 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_741_9_Right_791 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_742_9_Right_792 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_743_9_Right_793 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_744_9_Right_794 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_745_9_Right_795 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_746_9_Right_796 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_747_9_Right_797 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_748_9_Right_798 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_749_9_Right_799 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_750_9_Right_800 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_751_9_Right_801 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_752_9_Right_802 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_753_9_Right_803 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_754_9_Right_804 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_755_9_Right_805 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_756_9_Right_806 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_757_9_Right_807 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_758_9_Right_808 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_759_9_Right_809 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_760_9_Right_810 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_761_9_Right_811 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_762_9_Right_812 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_763_9_Right_813 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_764_9_Right_814 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_765_9_Right_815 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_766_9_Right_816 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_767_9_Right_817 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_768_9_Right_818 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_769_9_Right_819 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_770_9_Right_820 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_771_9_Right_821 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_772_9_Right_822 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_773_9_Right_823 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_774_9_Right_824 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_775_9_Right_825 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_776_9_Right_826 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_777_9_Right_827 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_778_9_Right_828 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_779_9_Right_829 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_780_9_Right_830 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_781_9_Right_831 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_782_9_Right_832 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_783_9_Right_833 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_784_9_Right_834 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_785_9_Right_835 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_786_9_Right_836 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_787_9_Right_837 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_788_9_Right_838 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_789_9_Right_839 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_790_9_Right_840 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_791_9_Right_841 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_792_9_Right_842 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_793_9_Right_843 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_794_9_Right_844 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_795_9_Right_845 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_796_9_Right_846 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_797_9_Right_847 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_798_9_Right_848 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_799_9_Right_849 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_800_9_Right_850 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_801_9_Right_851 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_802_9_Right_852 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_803_9_Right_853 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_804_9_Right_854 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_805_9_Right_855 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_806_9_Right_856 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_807_9_Right_857 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_808_9_Right_858 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_809_9_Right_859 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_810_9_Right_860 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_811_9_Right_861 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_812_9_Right_862 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_813_9_Right_863 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_814_9_Right_864 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_815_9_Right_865 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_816_9_Right_866 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_817_9_Right_867 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_818_9_Right_868 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_819_9_Right_869 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_820_9_Right_870 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_821_9_Right_871 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_822_9_Right_872 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_823_9_Right_873 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_824_9_Right_874 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_825_9_Right_875 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_826_9_Right_876 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_827_9_Right_877 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_828_9_Right_878 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_829_9_Right_879 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_830_9_Right_880 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_831_9_Right_881 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_832_9_Right_882 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_833_9_Right_883 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_834_9_Right_884 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_835_9_Right_885 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_836_9_Right_886 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_837_9_Right_887 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_838_9_Right_888 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_839_9_Right_889 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_840_9_Right_890 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_841_9_Right_891 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_842_9_Right_892 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_843_9_Right_893 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_844_9_Right_894 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_845_9_Right_895 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_846_9_Right_896 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_847_9_Right_897 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_848_9_Right_898 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_849_9_Right_899 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_850_9_Right_900 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_851_9_Right_901 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_852_9_Right_902 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_853_9_Right_903 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_854_9_Right_904 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_855_9_Right_905 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_856_9_Right_906 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_857_9_Right_907 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_858_9_Right_908 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_859_9_Right_909 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_860_9_Right_910 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_861_9_Right_911 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_862_9_Right_912 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_863_9_Right_913 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_864_9_Right_914 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_865_9_Right_915 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_866_9_Right_916 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_867_9_Right_917 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_868_9_Right_918 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_869_9_Right_919 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_870_9_Right_920 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_871_9_Right_921 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_872_9_Right_922 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_873_9_Right_923 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_874_9_Right_924 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_875_9_Right_925 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_876_9_Right_926 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_877_9_Right_927 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_878_9_Right_928 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_879_9_Right_929 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_880_9_Right_930 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_881_9_Right_931 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_894_9_Right_932 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_895_9_Right_933 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_896_9_Right_934 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_897_9_Right_935 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_898_9_Right_936 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_899_9_Right_937 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_900_9_Right_938 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_901_9_Right_939 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_902_9_Right_940 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_903_9_Right_941 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_904_9_Right_942 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_905_9_Right_943 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_906_9_Right_944 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_907_9_Right_945 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_908_9_Right_946 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_909_9_Right_947 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_910_9_Right_948 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_911_9_Right_949 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_912_9_Right_950 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_913_9_Right_951 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_914_9_Right_952 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_915_9_Right_953 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_916_9_Right_954 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_917_9_Right_955 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_918_9_Right_956 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_919_9_Right_957 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_920_9_Right_958 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_921_9_Right_959 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_922_9_Right_960 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_923_9_Right_961 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_924_9_Right_962 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_925_9_Right_963 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_926_9_Right_964 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_927_9_Right_965 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_928_9_Right_966 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_929_9_Right_967 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_930_9_Right_968 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_931_9_Right_969 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_932_9_Right_970 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_933_9_Right_971 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_934_9_Right_972 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_935_9_Right_973 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_936_9_Right_974 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_937_9_Right_975 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_938_9_Right_976 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_939_9_Right_977 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_940_9_Right_978 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_941_9_Right_979 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_942_9_Right_980 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_943_9_Right_981 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_944_9_Right_982 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_945_9_Right_983 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_946_9_Right_984 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_947_9_Right_985 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_948_9_Right_986 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_949_9_Right_987 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_950_9_Right_988 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_951_9_Right_989 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_952_9_Right_990 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_953_9_Right_991 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_954_9_Right_992 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_955_9_Right_993 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_956_9_Right_994 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_957_9_Right_995 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_958_9_Right_996 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_959_9_Right_997 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_960_9_Right_998 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_961_9_Right_999 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_962_9_Right_1000 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_963_9_Right_1001 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_964_9_Right_1002 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_965_9_Right_1003 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_966_9_Right_1004 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_967_9_Right_1005 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_968_9_Right_1006 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_969_9_Right_1007 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_970_9_Right_1008 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_971_9_Right_1009 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_972_9_Right_1010 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_973_9_Right_1011 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_974_9_Right_1012 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_975_9_Right_1013 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_976_9_Right_1014 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_977_9_Right_1015 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_978_9_Right_1016 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_979_9_Right_1017 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_980_9_Right_1018 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_981_9_Right_1019 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_982_9_Right_1020 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_983_9_Right_1021 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_984_9_Right_1022 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_985_9_Right_1023 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_986_9_Right_1024 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_987_9_Right_1025 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_988_9_Right_1026 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_989_9_Right_1027 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_990_9_Right_1028 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_991_9_Right_1029 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_992_9_Right_1030 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_993_9_Right_1031 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_994_9_Right_1032 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_995_9_Right_1033 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_996_9_Right_1034 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_997_9_Right_1035 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_998_9_Right_1036 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_999_9_Right_1037 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1000_9_Right_1038 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1001_9_Right_1039 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1002_9_Right_1040 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1003_9_Right_1041 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1004_9_Right_1042 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1005_9_Right_1043 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1006_9_Right_1044 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1007_9_Right_1045 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1008_9_Right_1046 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1009_9_Right_1047 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1010_9_Right_1048 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1011_9_Right_1049 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1012_9_Right_1050 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1013_9_Right_1051 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1014_9_Right_1052 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1015_9_Right_1053 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1016_9_Right_1054 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1017_9_Right_1055 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1018_9_Right_1056 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1019_9_Right_1057 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1020_9_Right_1058 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1021_9_Right_1059 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1022_9_Right_1060 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1023_9_Right_1061 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1024_9_Right_1062 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1025_9_Right_1063 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1026_9_Right_1064 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1027_9_Right_1065 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1028_9_Right_1066 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1029_9_Right_1067 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1030_9_Right_1068 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1031_9_Right_1069 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1032_9_Right_1070 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1033_9_Right_1071 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1034_9_Right_1072 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1035_9_Right_1073 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1036_9_Right_1074 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1037_9_Right_1075 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1038_9_Right_1076 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1039_9_Right_1077 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1040_9_Right_1078 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1041_9_Right_1079 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1042_9_Right_1080 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1043_9_Right_1081 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1044_9_Right_1082 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1045_9_Right_1083 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1046_9_Right_1084 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1047_9_Right_1085 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1048_9_Right_1086 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1049_9_Right_1087 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1050_9_Right_1088 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1051_9_Right_1089 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1052_9_Right_1090 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1053_9_Right_1091 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1054_9_Right_1092 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1055_9_Right_1093 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1056_9_Right_1094 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1057_9_Right_1095 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1070_9_Right_1096 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1071_9_Right_1097 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1072_9_Right_1098 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1073_9_Right_1099 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1074_9_Right_1100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1075_9_Right_1101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1076_9_Right_1102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1077_9_Right_1103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1078_9_Right_1104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1079_9_Right_1105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1080_9_Right_1106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1081_9_Right_1107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1082_9_Right_1108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1083_9_Right_1109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1084_9_Right_1110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1085_9_Right_1111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1086_9_Right_1112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1087_9_Right_1113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1088_9_Right_1114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1089_9_Right_1115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1090_9_Right_1116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1091_9_Right_1117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1092_9_Right_1118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1093_9_Right_1119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1094_9_Right_1120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1095_9_Right_1121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1096_9_Right_1122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1097_9_Right_1123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1098_9_Right_1124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1099_9_Right_1125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1100_9_Right_1126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1101_9_Right_1127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1102_9_Right_1128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1103_9_Right_1129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1104_9_Right_1130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1105_9_Right_1131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1106_9_Right_1132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1107_9_Right_1133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1108_9_Right_1134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1109_9_Right_1135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1110_9_Right_1136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1111_9_Right_1137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1112_9_Right_1138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1113_9_Right_1139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1114_9_Right_1140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1115_9_Right_1141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1116_9_Right_1142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1117_9_Right_1143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1118_9_Right_1144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1119_9_Right_1145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1120_9_Right_1146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1121_9_Right_1147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1122_9_Right_1148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1123_9_Right_1149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1124_9_Right_1150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1125_9_Right_1151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1126_9_Right_1152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1127_9_Right_1153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1128_9_Right_1154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1129_9_Right_1155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1130_9_Right_1156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1131_9_Right_1157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1132_9_Right_1158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1133_9_Right_1159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1134_9_Right_1160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1135_9_Right_1161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1136_9_Right_1162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1137_9_Right_1163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1138_9_Right_1164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1139_9_Right_1165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1140_9_Right_1166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1141_9_Right_1167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1142_9_Right_1168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1143_9_Right_1169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1144_9_Right_1170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1145_9_Right_1171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1146_9_Right_1172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1147_9_Right_1173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1148_9_Right_1174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1149_9_Right_1175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1150_9_Right_1176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1151_9_Right_1177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1152_9_Right_1178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1153_9_Right_1179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1154_9_Right_1180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1155_9_Right_1181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1156_9_Right_1182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1157_9_Right_1183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1158_9_Right_1184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1159_9_Right_1185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1160_9_Right_1186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1161_9_Right_1187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1162_9_Right_1188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1163_9_Right_1189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1164_9_Right_1190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1165_9_Right_1191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1166_9_Right_1192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1167_9_Right_1193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1168_9_Right_1194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1169_9_Right_1195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1170_9_Right_1196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1171_9_Right_1197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1172_9_Right_1198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1173_9_Right_1199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1174_9_Right_1200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1175_9_Right_1201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1176_9_Right_1202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1177_9_Right_1203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1178_9_Right_1204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1179_9_Right_1205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1180_9_Right_1206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1181_9_Right_1207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1182_9_Right_1208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1183_9_Right_1209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1184_9_Right_1210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1185_9_Right_1211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1186_9_Right_1212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1187_9_Right_1213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1188_9_Right_1214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1189_9_Right_1215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1190_9_Right_1216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1191_9_Right_1217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1192_9_Right_1218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1193_9_Right_1219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1194_9_Right_1220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1195_9_Right_1221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1196_9_Right_1222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1197_9_Right_1223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1198_9_Right_1224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1199_9_Right_1225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1200_9_Right_1226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1201_9_Right_1227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1202_9_Right_1228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1203_9_Right_1229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1204_9_Right_1230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1205_9_Right_1231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1206_9_Right_1232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1207_9_Right_1233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1208_9_Right_1234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1209_9_Right_1235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1210_9_Right_1236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1211_9_Right_1237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1212_9_Right_1238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1213_9_Right_1239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1214_9_Right_1240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1215_9_Right_1241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1216_9_Right_1242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1217_9_Right_1243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1218_9_Right_1244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1219_9_Right_1245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1220_9_Right_1246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1221_9_Right_1247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1222_9_Right_1248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1223_9_Right_1249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1224_9_Right_1250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1225_9_Right_1251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1226_9_Right_1252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1227_9_Right_1253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1228_9_Right_1254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1229_9_Right_1255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1230_9_Right_1256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1231_9_Right_1257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1232_9_Right_1258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1233_9_Right_1259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1246_9_Right_1260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1247_9_Right_1261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1248_9_Right_1262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1249_9_Right_1263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1250_9_Right_1264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1251_9_Right_1265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1252_9_Right_1266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1253_9_Right_1267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1254_9_Right_1268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1255_9_Right_1269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1256_9_Right_1270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1257_9_Right_1271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1258_9_Right_1272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1259_9_Right_1273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1260_9_Right_1274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1261_9_Right_1275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1262_9_Right_1276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1263_9_Right_1277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1264_9_Right_1278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1265_9_Right_1279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1266_9_Right_1280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1267_9_Right_1281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1268_9_Right_1282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1269_9_Right_1283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1270_9_Right_1284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1271_9_Right_1285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1272_9_Right_1286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1273_9_Right_1287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1274_9_Right_1288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1275_9_Right_1289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1276_9_Right_1290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1277_9_Right_1291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1278_9_Right_1292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1279_9_Right_1293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1280_9_Right_1294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1281_9_Right_1295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1282_9_Right_1296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1283_9_Right_1297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1284_9_Right_1298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1285_9_Right_1299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1286_9_Right_1300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1287_9_Right_1301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1288_9_Right_1302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1289_9_Right_1303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1290_9_Right_1304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1291_9_Right_1305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1292_9_Right_1306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1293_9_Right_1307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1294_9_Right_1308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1295_9_Right_1309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1296_9_Right_1310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1297_9_Right_1311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1298_9_Right_1312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1299_9_Right_1313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1300_9_Right_1314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1301_9_Right_1315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1302_9_Right_1316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1303_9_Right_1317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1304_9_Right_1318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1305_9_Right_1319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1306_9_Right_1320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1307_9_Right_1321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1308_9_Right_1322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1309_9_Right_1323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1310_9_Right_1324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1311_9_Right_1325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1312_9_Right_1326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1313_9_Right_1327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1314_9_Right_1328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1315_9_Right_1329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1316_9_Right_1330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1317_9_Right_1331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1318_9_Right_1332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1319_9_Right_1333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1320_9_Right_1334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1321_9_Right_1335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1322_9_Right_1336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1323_9_Right_1337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1324_9_Right_1338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1325_9_Right_1339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1326_9_Right_1340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1327_9_Right_1341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1328_9_Right_1342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1329_9_Right_1343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1330_9_Right_1344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1331_9_Right_1345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1332_9_Right_1346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1333_9_Right_1347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1334_9_Right_1348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1335_9_Right_1349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1336_9_Right_1350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1337_9_Right_1351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1338_9_Right_1352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1339_9_Right_1353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1340_9_Right_1354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1341_9_Right_1355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1342_9_Right_1356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1343_9_Right_1357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1344_9_Right_1358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1345_9_Right_1359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1346_9_Right_1360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1347_9_Right_1361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1348_9_Right_1362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1349_9_Right_1363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1350_9_Right_1364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1351_9_Right_1365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1352_9_Right_1366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1353_9_Right_1367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1354_9_Right_1368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1355_9_Right_1369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1356_9_Right_1370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1357_9_Right_1371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1358_9_Right_1372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1359_9_Right_1373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1360_9_Right_1374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1361_9_Right_1375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1362_9_Right_1376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1363_9_Right_1377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1364_9_Right_1378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1365_9_Right_1379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1366_9_Right_1380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1367_9_Right_1381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1368_9_Right_1382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1369_9_Right_1383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1370_9_Right_1384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1371_9_Right_1385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1372_9_Right_1386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1373_9_Right_1387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1374_9_Right_1388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1375_9_Right_1389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1376_9_Right_1390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1377_9_Right_1391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1378_9_Right_1392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1379_9_Right_1393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1380_9_Right_1394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1381_9_Right_1395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1382_9_Right_1396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1383_9_Right_1397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1384_9_Right_1398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1385_9_Right_1399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1386_9_Right_1400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1387_9_Right_1401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1388_9_Right_1402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1389_9_Right_1403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1390_9_Right_1404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1391_9_Right_1405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1392_9_Right_1406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1393_9_Right_1407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1394_9_Right_1408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1395_9_Right_1409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1396_9_Right_1410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1397_9_Right_1411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1398_9_Right_1412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1399_9_Right_1413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1400_9_Right_1414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1401_9_Right_1415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1402_9_Right_1416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1403_9_Right_1417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1404_9_Right_1418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1405_9_Right_1419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1406_9_Right_1420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1407_9_Right_1421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1408_9_Right_1422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1409_9_Right_1423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_1424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_1425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_1426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_1427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_1428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_1429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_1430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_1431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_1432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_1433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_1434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_1435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_1436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_1437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_1_Left_1438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_1_Left_1439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_1_Left_1440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_1_Left_1441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_1_Left_1442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_1_Left_1443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_1_Left_1444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_1_Left_1445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_1_Left_1446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_1_Left_1447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_1_Left_1448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_1_Left_1449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_1_Left_1450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_1_Left_1451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_1_Left_1452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_1_Left_1453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_1_Left_1454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_1_Left_1455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_1_Left_1456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_1_Left_1457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_1_Left_1458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_1_Left_1459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_1_Left_1460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_1_Left_1461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_1_Left_1462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_1_Left_1463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_1_Left_1464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_1_Left_1465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_1_Left_1466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_1_Left_1467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_1_Left_1468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_1_Left_1469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_1_Left_1470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_1_Left_1471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_1_Left_1472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_1_Left_1473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_1_Left_1474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_1_Left_1475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_1_Left_1476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_1_Left_1477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_1_Left_1478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_1_Left_1479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_1_Left_1480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_1_Left_1481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_1_Left_1482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_1_Left_1483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_1_Left_1484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_1_Left_1485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_1_Left_1486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_1_Left_1487 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_1_Left_1488 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_1_Left_1489 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_1_Left_1490 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_1_Left_1491 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_1_Left_1492 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_1_Left_1493 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_1_Left_1494 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_1_Left_1495 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_1_Left_1496 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_1_Left_1497 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_1_Left_1498 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_1_Left_1499 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_1_Left_1500 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_1_Left_1501 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_1_Left_1502 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_1_Left_1503 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_1_Left_1504 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_1_Left_1505 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_1_Left_1506 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_1_Left_1507 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_1_Left_1508 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_1_Left_1509 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_1_Left_1510 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_1_Left_1511 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_1_Left_1512 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_1_Left_1513 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_1_Left_1514 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_1_Left_1515 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_1_Left_1516 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_1_Left_1517 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_1_Left_1518 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_1_Left_1519 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_1_Left_1520 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_1_Left_1521 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_1_Left_1522 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_1_Left_1523 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_1_Left_1524 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_1_Left_1525 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_1_Left_1526 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_1_Left_1527 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_1_Left_1528 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_1_Left_1529 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_1_Left_1530 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_1_Left_1531 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_1_Left_1532 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_1_Left_1533 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_1_Left_1534 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_1_Left_1535 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_1_Left_1536 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_1_Left_1537 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_1_Left_1538 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_1_Left_1539 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_1_Left_1540 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_1_Left_1541 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_1_Left_1542 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_1_Left_1543 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_1_Left_1544 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_1_Left_1545 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_1_Left_1546 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_1_Left_1547 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_1_Left_1548 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_1_Left_1549 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_1_Left_1550 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_1_Left_1551 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_1_Left_1552 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_1_Left_1553 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_1_Left_1554 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_1_Left_1555 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_1_Left_1556 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_1_Left_1557 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_1_Left_1558 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_1_Left_1559 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_1_Left_1560 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_1_Left_1561 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_1_Left_1562 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_1_Left_1563 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_1_Left_1564 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_1_Left_1565 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_1_Left_1566 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_1_Left_1567 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_1_Left_1568 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_1_Left_1569 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_1_Left_1570 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_1_Left_1571 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_1_Left_1572 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_1_Left_1573 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_1_Left_1574 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_1_Left_1575 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_1_Left_1576 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_1_Left_1577 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_1_Left_1578 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_1_Left_1579 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_1_Left_1580 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_1_Left_1581 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_1_Left_1582 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_1_Left_1583 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_1_Left_1584 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_1_Left_1585 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_1_Left_1586 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_1_Left_1587 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_1_Left_1588 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_1_Left_1589 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_1_Left_1590 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_1_Left_1591 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_1_Left_1592 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_1_Left_1593 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_1_Left_1594 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_1_Left_1595 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_1_Left_1596 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_1_Left_1597 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_1_Left_1598 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_1_Left_1599 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_1_Left_1600 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_1_Left_1601 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_178_Left_1602 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_179_Left_1603 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_180_Left_1604 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_181_Left_1605 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_182_Left_1606 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_183_Left_1607 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_184_Left_1608 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_185_Left_1609 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_186_Left_1610 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_187_Left_1611 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_188_Left_1612 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_189_Left_1613 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_1_Left_1614 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_1_Left_1615 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_1_Left_1616 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_1_Left_1617 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_1_Left_1618 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_1_Left_1619 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_1_Left_1620 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_1_Left_1621 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_1_Left_1622 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_1_Left_1623 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_1_Left_1624 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_1_Left_1625 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_1_Left_1626 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_1_Left_1627 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_1_Left_1628 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_1_Left_1629 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_1_Left_1630 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_1_Left_1631 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_1_Left_1632 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_1_Left_1633 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_1_Left_1634 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_1_Left_1635 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_1_Left_1636 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_1_Left_1637 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_1_Left_1638 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_1_Left_1639 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_1_Left_1640 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_1_Left_1641 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_1_Left_1642 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_1_Left_1643 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_1_Left_1644 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_1_Left_1645 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_1_Left_1646 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_1_Left_1647 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_1_Left_1648 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_1_Left_1649 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_1_Left_1650 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_1_Left_1651 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_1_Left_1652 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_1_Left_1653 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_1_Left_1654 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_1_Left_1655 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_1_Left_1656 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_1_Left_1657 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_1_Left_1658 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_1_Left_1659 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_1_Left_1660 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_1_Left_1661 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_1_Left_1662 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_1_Left_1663 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_1_Left_1664 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_1_Left_1665 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_1_Left_1666 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_1_Left_1667 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_1_Left_1668 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_1_Left_1669 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_1_Left_1670 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_1_Left_1671 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_1_Left_1672 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_1_Left_1673 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_1_Left_1674 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_1_Left_1675 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_1_Left_1676 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_1_Left_1677 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_1_Left_1678 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_1_Left_1679 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_1_Left_1680 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_1_Left_1681 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_1_Left_1682 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_1_Left_1683 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_1_Left_1684 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_1_Left_1685 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_1_Left_1686 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_1_Left_1687 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_1_Left_1688 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_1_Left_1689 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_1_Left_1690 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_1_Left_1691 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_1_Left_1692 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_1_Left_1693 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_1_Left_1694 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_1_Left_1695 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_1_Left_1696 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_1_Left_1697 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_1_Left_1698 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_1_Left_1699 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_1_Left_1700 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_1_Left_1701 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_1_Left_1702 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_1_Left_1703 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_1_Left_1704 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_1_Left_1705 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_1_Left_1706 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_1_Left_1707 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_1_Left_1708 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_1_Left_1709 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_1_Left_1710 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_1_Left_1711 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_1_Left_1712 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_1_Left_1713 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_1_Left_1714 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_1_Left_1715 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_1_Left_1716 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_1_Left_1717 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_295_1_Left_1718 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_296_1_Left_1719 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_297_1_Left_1720 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_298_1_Left_1721 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_299_1_Left_1722 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_300_1_Left_1723 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_301_1_Left_1724 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_302_1_Left_1725 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_303_1_Left_1726 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_304_1_Left_1727 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_305_1_Left_1728 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_306_1_Left_1729 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_307_1_Left_1730 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_308_1_Left_1731 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_309_1_Left_1732 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_310_1_Left_1733 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_311_1_Left_1734 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_312_1_Left_1735 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_313_1_Left_1736 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_314_1_Left_1737 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_315_1_Left_1738 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_316_1_Left_1739 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_317_1_Left_1740 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_318_1_Left_1741 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_319_1_Left_1742 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_320_1_Left_1743 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_321_1_Left_1744 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_322_1_Left_1745 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_323_1_Left_1746 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_324_1_Left_1747 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_325_1_Left_1748 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_326_1_Left_1749 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_327_1_Left_1750 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_328_1_Left_1751 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_329_1_Left_1752 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_330_1_Left_1753 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_331_1_Left_1754 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_332_1_Left_1755 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_333_1_Left_1756 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_334_1_Left_1757 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_335_1_Left_1758 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_336_1_Left_1759 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_337_1_Left_1760 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_338_1_Left_1761 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_339_1_Left_1762 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_340_1_Left_1763 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_341_1_Left_1764 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_342_1_Left_1765 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_343_1_Left_1766 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_344_1_Left_1767 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_345_1_Left_1768 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_346_1_Left_1769 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_347_1_Left_1770 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_348_1_Left_1771 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_349_1_Left_1772 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_350_1_Left_1773 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_351_1_Left_1774 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_352_1_Left_1775 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_353_1_Left_1776 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_366_1_Left_1777 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_354_Left_1778 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_355_Left_1779 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_356_Left_1780 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_357_Left_1781 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_358_Left_1782 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_359_Left_1783 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_360_Left_1784 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_361_Left_1785 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_362_Left_1786 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_363_Left_1787 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_364_Left_1788 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_365_Left_1789 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_367_1_Left_1790 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_368_1_Left_1791 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_369_1_Left_1792 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_370_1_Left_1793 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_371_1_Left_1794 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_372_1_Left_1795 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_373_1_Left_1796 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_374_1_Left_1797 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_375_1_Left_1798 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_376_1_Left_1799 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_377_1_Left_1800 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_378_1_Left_1801 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_379_1_Left_1802 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_380_1_Left_1803 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_381_1_Left_1804 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_382_1_Left_1805 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_383_1_Left_1806 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_384_1_Left_1807 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_385_1_Left_1808 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_386_1_Left_1809 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_387_1_Left_1810 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_388_1_Left_1811 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_389_1_Left_1812 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_390_1_Left_1813 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_391_1_Left_1814 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_392_1_Left_1815 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_393_1_Left_1816 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_394_1_Left_1817 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_395_1_Left_1818 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_396_1_Left_1819 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_397_1_Left_1820 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_398_1_Left_1821 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_399_1_Left_1822 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_400_1_Left_1823 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_401_1_Left_1824 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_402_1_Left_1825 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_403_1_Left_1826 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_404_1_Left_1827 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_405_1_Left_1828 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_406_1_Left_1829 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_407_1_Left_1830 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_408_1_Left_1831 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_409_1_Left_1832 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_410_1_Left_1833 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_411_1_Left_1834 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_412_1_Left_1835 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_413_1_Left_1836 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_414_1_Left_1837 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_415_1_Left_1838 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_416_1_Left_1839 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_417_1_Left_1840 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_418_1_Left_1841 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_419_1_Left_1842 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_420_1_Left_1843 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_421_1_Left_1844 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_422_1_Left_1845 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_423_1_Left_1846 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_424_1_Left_1847 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_425_1_Left_1848 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_426_1_Left_1849 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_427_1_Left_1850 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_428_1_Left_1851 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_429_1_Left_1852 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_430_1_Left_1853 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_431_1_Left_1854 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_432_1_Left_1855 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_433_1_Left_1856 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_434_1_Left_1857 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_435_1_Left_1858 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_436_1_Left_1859 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_437_1_Left_1860 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_438_1_Left_1861 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_439_1_Left_1862 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_440_1_Left_1863 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_441_1_Left_1864 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_442_1_Left_1865 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_443_1_Left_1866 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_444_1_Left_1867 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_445_1_Left_1868 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_446_1_Left_1869 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_447_1_Left_1870 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_448_1_Left_1871 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_449_1_Left_1872 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_450_1_Left_1873 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_451_1_Left_1874 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_452_1_Left_1875 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_453_1_Left_1876 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_454_1_Left_1877 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_455_1_Left_1878 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_456_1_Left_1879 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_457_1_Left_1880 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_458_1_Left_1881 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_459_1_Left_1882 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_460_1_Left_1883 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_461_1_Left_1884 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_462_1_Left_1885 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_463_1_Left_1886 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_464_1_Left_1887 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_465_1_Left_1888 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_466_1_Left_1889 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_467_1_Left_1890 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_468_1_Left_1891 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_469_1_Left_1892 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_470_1_Left_1893 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_471_1_Left_1894 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_472_1_Left_1895 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_473_1_Left_1896 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_474_1_Left_1897 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_475_1_Left_1898 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_476_1_Left_1899 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_477_1_Left_1900 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_478_1_Left_1901 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_479_1_Left_1902 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_480_1_Left_1903 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_481_1_Left_1904 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_482_1_Left_1905 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_483_1_Left_1906 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_484_1_Left_1907 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_485_1_Left_1908 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_486_1_Left_1909 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_487_1_Left_1910 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_488_1_Left_1911 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_489_1_Left_1912 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_490_1_Left_1913 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_491_1_Left_1914 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_492_1_Left_1915 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_493_1_Left_1916 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_494_1_Left_1917 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_495_1_Left_1918 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_496_1_Left_1919 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_497_1_Left_1920 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_498_1_Left_1921 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_499_1_Left_1922 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_500_1_Left_1923 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_501_1_Left_1924 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_502_1_Left_1925 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_503_1_Left_1926 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_504_1_Left_1927 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_505_1_Left_1928 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_506_1_Left_1929 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_507_1_Left_1930 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_508_1_Left_1931 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_509_1_Left_1932 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_510_1_Left_1933 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_511_1_Left_1934 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_512_1_Left_1935 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_513_1_Left_1936 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_514_1_Left_1937 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_515_1_Left_1938 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_516_1_Left_1939 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_517_1_Left_1940 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_518_1_Left_1941 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_519_1_Left_1942 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_520_1_Left_1943 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_521_1_Left_1944 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_522_1_Left_1945 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_523_1_Left_1946 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_524_1_Left_1947 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_525_1_Left_1948 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_526_1_Left_1949 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_527_1_Left_1950 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_528_1_Left_1951 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_529_1_Left_1952 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_542_1_Left_1953 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_530_Left_1954 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_531_Left_1955 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_532_Left_1956 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_533_Left_1957 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_534_Left_1958 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_535_Left_1959 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_536_Left_1960 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_537_Left_1961 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_538_Left_1962 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_539_Left_1963 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_540_Left_1964 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_541_Left_1965 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_543_1_Left_1966 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_544_1_Left_1967 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_545_1_Left_1968 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_546_1_Left_1969 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_547_1_Left_1970 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_548_1_Left_1971 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_549_1_Left_1972 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_550_1_Left_1973 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_551_1_Left_1974 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_552_1_Left_1975 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_553_1_Left_1976 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_554_1_Left_1977 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_555_1_Left_1978 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_556_1_Left_1979 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_557_1_Left_1980 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_558_1_Left_1981 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_559_1_Left_1982 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_560_1_Left_1983 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_561_1_Left_1984 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_562_1_Left_1985 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_563_1_Left_1986 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_564_1_Left_1987 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_565_1_Left_1988 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_566_1_Left_1989 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_567_1_Left_1990 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_568_1_Left_1991 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_569_1_Left_1992 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_570_1_Left_1993 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_571_1_Left_1994 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_572_1_Left_1995 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_573_1_Left_1996 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_574_1_Left_1997 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_575_1_Left_1998 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_576_1_Left_1999 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_577_1_Left_2000 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_578_1_Left_2001 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_579_1_Left_2002 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_580_1_Left_2003 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_581_1_Left_2004 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_582_1_Left_2005 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_583_1_Left_2006 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_584_1_Left_2007 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_585_1_Left_2008 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_586_1_Left_2009 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_587_1_Left_2010 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_588_1_Left_2011 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_589_1_Left_2012 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_590_1_Left_2013 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_591_1_Left_2014 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_592_1_Left_2015 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_593_1_Left_2016 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_594_1_Left_2017 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_595_1_Left_2018 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_596_1_Left_2019 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_597_1_Left_2020 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_598_1_Left_2021 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_599_1_Left_2022 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_600_1_Left_2023 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_601_1_Left_2024 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_602_1_Left_2025 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_603_1_Left_2026 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_604_1_Left_2027 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_605_1_Left_2028 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_606_1_Left_2029 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_607_1_Left_2030 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_608_1_Left_2031 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_609_1_Left_2032 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_610_1_Left_2033 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_611_1_Left_2034 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_612_1_Left_2035 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_613_1_Left_2036 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_614_1_Left_2037 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_615_1_Left_2038 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_616_1_Left_2039 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_617_1_Left_2040 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_618_1_Left_2041 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_619_1_Left_2042 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_620_1_Left_2043 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_621_1_Left_2044 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_622_1_Left_2045 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_623_1_Left_2046 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_624_1_Left_2047 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_625_1_Left_2048 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_626_1_Left_2049 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_627_1_Left_2050 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_628_1_Left_2051 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_629_1_Left_2052 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_630_1_Left_2053 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_631_1_Left_2054 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_632_1_Left_2055 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_633_1_Left_2056 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_634_1_Left_2057 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_635_1_Left_2058 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_636_1_Left_2059 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_637_1_Left_2060 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_638_1_Left_2061 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_639_1_Left_2062 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_640_1_Left_2063 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_641_1_Left_2064 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_642_1_Left_2065 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_643_1_Left_2066 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_644_1_Left_2067 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_645_1_Left_2068 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_646_1_Left_2069 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_647_1_Left_2070 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_648_1_Left_2071 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_649_1_Left_2072 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_650_1_Left_2073 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_651_1_Left_2074 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_652_1_Left_2075 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_653_1_Left_2076 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_654_1_Left_2077 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_655_1_Left_2078 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_656_1_Left_2079 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_657_1_Left_2080 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_658_1_Left_2081 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_659_1_Left_2082 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_660_1_Left_2083 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_661_1_Left_2084 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_662_1_Left_2085 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_663_1_Left_2086 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_664_1_Left_2087 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_665_1_Left_2088 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_666_1_Left_2089 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_667_1_Left_2090 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_668_1_Left_2091 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_669_1_Left_2092 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_670_1_Left_2093 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_671_1_Left_2094 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_672_1_Left_2095 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_673_1_Left_2096 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_674_1_Left_2097 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_675_1_Left_2098 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_676_1_Left_2099 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_677_1_Left_2100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_678_1_Left_2101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_679_1_Left_2102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_680_1_Left_2103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_681_1_Left_2104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_682_1_Left_2105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_683_1_Left_2106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_684_1_Left_2107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_685_1_Left_2108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_686_1_Left_2109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_687_1_Left_2110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_688_1_Left_2111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_689_1_Left_2112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_690_1_Left_2113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_691_1_Left_2114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_692_1_Left_2115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_693_1_Left_2116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_694_1_Left_2117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_695_1_Left_2118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_696_1_Left_2119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_697_1_Left_2120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_698_1_Left_2121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_699_1_Left_2122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_700_1_Left_2123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_701_1_Left_2124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_702_1_Left_2125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_703_1_Left_2126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_704_1_Left_2127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_705_1_Left_2128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_718_1_Left_2129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_706_Left_2130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_707_Left_2131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_708_Left_2132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_709_Left_2133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_710_Left_2134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_711_Left_2135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_712_Left_2136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_713_Left_2137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_714_Left_2138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_715_Left_2139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_716_Left_2140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_717_Left_2141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_719_1_Left_2142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_720_1_Left_2143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_721_1_Left_2144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_722_1_Left_2145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_723_1_Left_2146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_724_1_Left_2147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_725_1_Left_2148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_726_1_Left_2149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_727_1_Left_2150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_728_1_Left_2151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_729_1_Left_2152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_730_1_Left_2153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_731_1_Left_2154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_732_1_Left_2155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_733_1_Left_2156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_734_1_Left_2157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_735_1_Left_2158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_736_1_Left_2159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_737_1_Left_2160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_738_1_Left_2161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_739_1_Left_2162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_740_1_Left_2163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_741_1_Left_2164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_742_1_Left_2165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_743_1_Left_2166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_744_1_Left_2167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_745_1_Left_2168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_746_1_Left_2169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_747_1_Left_2170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_748_1_Left_2171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_749_1_Left_2172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_750_1_Left_2173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_751_1_Left_2174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_752_1_Left_2175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_753_1_Left_2176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_754_1_Left_2177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_755_1_Left_2178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_756_1_Left_2179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_757_1_Left_2180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_758_1_Left_2181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_759_1_Left_2182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_760_1_Left_2183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_761_1_Left_2184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_762_1_Left_2185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_763_1_Left_2186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_764_1_Left_2187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_765_1_Left_2188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_766_1_Left_2189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_767_1_Left_2190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_768_1_Left_2191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_769_1_Left_2192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_770_1_Left_2193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_771_1_Left_2194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_772_1_Left_2195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_773_1_Left_2196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_774_1_Left_2197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_775_1_Left_2198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_776_1_Left_2199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_777_1_Left_2200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_778_1_Left_2201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_779_1_Left_2202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_780_1_Left_2203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_781_1_Left_2204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_782_1_Left_2205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_783_1_Left_2206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_784_1_Left_2207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_785_1_Left_2208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_786_1_Left_2209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_787_1_Left_2210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_788_1_Left_2211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_789_1_Left_2212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_790_1_Left_2213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_791_1_Left_2214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_792_1_Left_2215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_793_1_Left_2216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_794_1_Left_2217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_795_1_Left_2218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_796_1_Left_2219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_797_1_Left_2220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_798_1_Left_2221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_799_1_Left_2222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_800_1_Left_2223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_801_1_Left_2224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_802_1_Left_2225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_803_1_Left_2226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_804_1_Left_2227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_805_1_Left_2228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_806_1_Left_2229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_807_1_Left_2230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_808_1_Left_2231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_809_1_Left_2232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_810_1_Left_2233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_811_1_Left_2234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_812_1_Left_2235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_813_1_Left_2236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_814_1_Left_2237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_815_1_Left_2238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_816_1_Left_2239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_817_1_Left_2240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_818_1_Left_2241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_819_1_Left_2242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_820_1_Left_2243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_821_1_Left_2244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_822_1_Left_2245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_823_1_Left_2246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_824_1_Left_2247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_825_1_Left_2248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_826_1_Left_2249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_827_1_Left_2250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_828_1_Left_2251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_829_1_Left_2252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_830_1_Left_2253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_831_1_Left_2254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_832_1_Left_2255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_833_1_Left_2256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_834_1_Left_2257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_835_1_Left_2258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_836_1_Left_2259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_837_1_Left_2260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_838_1_Left_2261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_839_1_Left_2262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_840_1_Left_2263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_841_1_Left_2264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_842_1_Left_2265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_843_1_Left_2266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_844_1_Left_2267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_845_1_Left_2268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_846_1_Left_2269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_847_1_Left_2270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_848_1_Left_2271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_849_1_Left_2272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_850_1_Left_2273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_851_1_Left_2274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_852_1_Left_2275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_853_1_Left_2276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_854_1_Left_2277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_855_1_Left_2278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_856_1_Left_2279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_857_1_Left_2280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_858_1_Left_2281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_859_1_Left_2282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_860_1_Left_2283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_861_1_Left_2284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_862_1_Left_2285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_863_1_Left_2286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_864_1_Left_2287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_865_1_Left_2288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_866_1_Left_2289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_867_1_Left_2290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_868_1_Left_2291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_869_1_Left_2292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_870_1_Left_2293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_871_1_Left_2294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_872_1_Left_2295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_873_1_Left_2296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_874_1_Left_2297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_875_1_Left_2298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_876_1_Left_2299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_877_1_Left_2300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_878_1_Left_2301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_879_1_Left_2302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_880_1_Left_2303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_881_1_Left_2304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_894_1_Left_2305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_882_Left_2306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_883_Left_2307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_884_Left_2308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_885_Left_2309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_886_Left_2310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_887_Left_2311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_888_Left_2312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_889_Left_2313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_890_Left_2314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_891_Left_2315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_892_Left_2316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_893_Left_2317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_895_1_Left_2318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_896_1_Left_2319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_897_1_Left_2320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_898_1_Left_2321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_899_1_Left_2322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_900_1_Left_2323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_901_1_Left_2324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_902_1_Left_2325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_903_1_Left_2326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_904_1_Left_2327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_905_1_Left_2328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_906_1_Left_2329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_907_1_Left_2330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_908_1_Left_2331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_909_1_Left_2332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_910_1_Left_2333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_911_1_Left_2334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_912_1_Left_2335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_913_1_Left_2336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_914_1_Left_2337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_915_1_Left_2338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_916_1_Left_2339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_917_1_Left_2340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_918_1_Left_2341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_919_1_Left_2342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_920_1_Left_2343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_921_1_Left_2344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_922_1_Left_2345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_923_1_Left_2346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_924_1_Left_2347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_925_1_Left_2348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_926_1_Left_2349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_927_1_Left_2350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_928_1_Left_2351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_929_1_Left_2352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_930_1_Left_2353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_931_1_Left_2354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_932_1_Left_2355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_933_1_Left_2356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_934_1_Left_2357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_935_1_Left_2358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_936_1_Left_2359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_937_1_Left_2360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_938_1_Left_2361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_939_1_Left_2362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_940_1_Left_2363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_941_1_Left_2364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_942_1_Left_2365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_943_1_Left_2366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_944_1_Left_2367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_945_1_Left_2368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_946_1_Left_2369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_947_1_Left_2370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_948_1_Left_2371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_949_1_Left_2372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_950_1_Left_2373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_951_1_Left_2374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_952_1_Left_2375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_953_1_Left_2376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_954_1_Left_2377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_955_1_Left_2378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_956_1_Left_2379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_957_1_Left_2380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_958_1_Left_2381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_959_1_Left_2382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_960_1_Left_2383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_961_1_Left_2384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_962_1_Left_2385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_963_1_Left_2386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_964_1_Left_2387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_965_1_Left_2388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_966_1_Left_2389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_967_1_Left_2390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_968_1_Left_2391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_969_1_Left_2392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_970_1_Left_2393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_971_1_Left_2394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_972_1_Left_2395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_973_1_Left_2396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_974_1_Left_2397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_975_1_Left_2398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_976_1_Left_2399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_977_1_Left_2400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_978_1_Left_2401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_979_1_Left_2402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_980_1_Left_2403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_981_1_Left_2404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_982_1_Left_2405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_983_1_Left_2406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_984_1_Left_2407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_985_1_Left_2408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_986_1_Left_2409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_987_1_Left_2410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_988_1_Left_2411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_989_1_Left_2412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_990_1_Left_2413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_991_1_Left_2414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_992_1_Left_2415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_993_1_Left_2416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_994_1_Left_2417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_995_1_Left_2418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_996_1_Left_2419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_997_1_Left_2420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_998_1_Left_2421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_999_1_Left_2422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1000_1_Left_2423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1001_1_Left_2424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1002_1_Left_2425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1003_1_Left_2426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1004_1_Left_2427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1005_1_Left_2428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1006_1_Left_2429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1007_1_Left_2430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1008_1_Left_2431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1009_1_Left_2432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1010_1_Left_2433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1011_1_Left_2434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1012_1_Left_2435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1013_1_Left_2436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1014_1_Left_2437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1015_1_Left_2438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1016_1_Left_2439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1017_1_Left_2440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1018_1_Left_2441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1019_1_Left_2442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1020_1_Left_2443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1021_1_Left_2444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1022_1_Left_2445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1023_1_Left_2446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1024_1_Left_2447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1025_1_Left_2448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1026_1_Left_2449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1027_1_Left_2450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1028_1_Left_2451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1029_1_Left_2452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1030_1_Left_2453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1031_1_Left_2454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1032_1_Left_2455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1033_1_Left_2456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1034_1_Left_2457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1035_1_Left_2458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1036_1_Left_2459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1037_1_Left_2460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1038_1_Left_2461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1039_1_Left_2462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1040_1_Left_2463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1041_1_Left_2464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1042_1_Left_2465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1043_1_Left_2466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1044_1_Left_2467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1045_1_Left_2468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1046_1_Left_2469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1047_1_Left_2470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1048_1_Left_2471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1049_1_Left_2472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1050_1_Left_2473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1051_1_Left_2474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1052_1_Left_2475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1053_1_Left_2476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1054_1_Left_2477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1055_1_Left_2478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1056_1_Left_2479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1057_1_Left_2480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1070_1_Left_2481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1058_Left_2482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1059_Left_2483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1060_Left_2484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1061_Left_2485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1062_Left_2486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1063_Left_2487 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1064_Left_2488 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1065_Left_2489 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1066_Left_2490 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1067_Left_2491 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1068_Left_2492 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1069_Left_2493 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1071_1_Left_2494 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1072_1_Left_2495 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1073_1_Left_2496 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1074_1_Left_2497 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1075_1_Left_2498 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1076_1_Left_2499 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1077_1_Left_2500 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1078_1_Left_2501 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1079_1_Left_2502 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1080_1_Left_2503 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1081_1_Left_2504 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1082_1_Left_2505 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1083_1_Left_2506 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1084_1_Left_2507 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1085_1_Left_2508 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1086_1_Left_2509 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1087_1_Left_2510 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1088_1_Left_2511 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1089_1_Left_2512 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1090_1_Left_2513 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1091_1_Left_2514 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1092_1_Left_2515 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1093_1_Left_2516 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1094_1_Left_2517 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1095_1_Left_2518 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1096_1_Left_2519 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1097_1_Left_2520 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1098_1_Left_2521 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1099_1_Left_2522 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1100_1_Left_2523 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1101_1_Left_2524 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1102_1_Left_2525 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1103_1_Left_2526 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1104_1_Left_2527 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1105_1_Left_2528 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1106_1_Left_2529 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1107_1_Left_2530 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1108_1_Left_2531 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1109_1_Left_2532 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1110_1_Left_2533 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1111_1_Left_2534 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1112_1_Left_2535 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1113_1_Left_2536 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1114_1_Left_2537 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1115_1_Left_2538 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1116_1_Left_2539 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1117_1_Left_2540 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1118_1_Left_2541 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1119_1_Left_2542 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1120_1_Left_2543 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1121_1_Left_2544 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1122_1_Left_2545 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1123_1_Left_2546 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1124_1_Left_2547 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1125_1_Left_2548 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1126_1_Left_2549 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1127_1_Left_2550 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1128_1_Left_2551 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1129_1_Left_2552 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1130_1_Left_2553 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1131_1_Left_2554 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1132_1_Left_2555 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1133_1_Left_2556 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1134_1_Left_2557 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1135_1_Left_2558 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1136_1_Left_2559 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1137_1_Left_2560 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1138_1_Left_2561 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1139_1_Left_2562 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1140_1_Left_2563 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1141_1_Left_2564 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1142_1_Left_2565 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1143_1_Left_2566 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1144_1_Left_2567 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1145_1_Left_2568 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1146_1_Left_2569 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1147_1_Left_2570 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1148_1_Left_2571 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1149_1_Left_2572 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1150_1_Left_2573 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1151_1_Left_2574 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1152_1_Left_2575 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1153_1_Left_2576 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1154_1_Left_2577 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1155_1_Left_2578 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1156_1_Left_2579 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1157_1_Left_2580 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1158_1_Left_2581 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1159_1_Left_2582 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1160_1_Left_2583 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1161_1_Left_2584 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1162_1_Left_2585 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1163_1_Left_2586 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1164_1_Left_2587 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1165_1_Left_2588 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1166_1_Left_2589 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1167_1_Left_2590 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1168_1_Left_2591 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1169_1_Left_2592 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1170_1_Left_2593 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1171_1_Left_2594 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1172_1_Left_2595 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1173_1_Left_2596 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1174_1_Left_2597 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1175_1_Left_2598 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1176_1_Left_2599 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1177_1_Left_2600 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1178_1_Left_2601 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1179_1_Left_2602 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1180_1_Left_2603 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1181_1_Left_2604 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1182_1_Left_2605 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1183_1_Left_2606 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1184_1_Left_2607 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1185_1_Left_2608 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1186_1_Left_2609 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1187_1_Left_2610 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1188_1_Left_2611 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1189_1_Left_2612 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1190_1_Left_2613 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1191_1_Left_2614 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1192_1_Left_2615 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1193_1_Left_2616 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1194_1_Left_2617 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1195_1_Left_2618 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1196_1_Left_2619 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1197_1_Left_2620 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1198_1_Left_2621 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1199_1_Left_2622 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1200_1_Left_2623 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1201_1_Left_2624 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1202_1_Left_2625 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1203_1_Left_2626 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1204_1_Left_2627 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1205_1_Left_2628 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1206_1_Left_2629 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1207_1_Left_2630 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1208_1_Left_2631 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1209_1_Left_2632 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1210_1_Left_2633 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1211_1_Left_2634 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1212_1_Left_2635 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1213_1_Left_2636 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1214_1_Left_2637 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1215_1_Left_2638 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1216_1_Left_2639 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1217_1_Left_2640 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1218_1_Left_2641 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1219_1_Left_2642 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1220_1_Left_2643 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1221_1_Left_2644 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1222_1_Left_2645 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1223_1_Left_2646 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1224_1_Left_2647 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1225_1_Left_2648 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1226_1_Left_2649 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1227_1_Left_2650 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1228_1_Left_2651 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1229_1_Left_2652 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1230_1_Left_2653 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1231_1_Left_2654 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1232_1_Left_2655 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1233_1_Left_2656 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1246_1_Left_2657 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1234_Left_2658 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1235_Left_2659 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1236_Left_2660 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1237_Left_2661 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1238_Left_2662 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1239_Left_2663 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1240_Left_2664 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1241_Left_2665 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1242_Left_2666 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1243_Left_2667 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1244_Left_2668 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1245_Left_2669 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1247_1_Left_2670 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1248_1_Left_2671 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1249_1_Left_2672 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1250_1_Left_2673 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1251_1_Left_2674 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1252_1_Left_2675 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1253_1_Left_2676 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1254_1_Left_2677 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1255_1_Left_2678 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1256_1_Left_2679 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1257_1_Left_2680 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1258_1_Left_2681 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1259_1_Left_2682 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1260_1_Left_2683 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1261_1_Left_2684 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1262_1_Left_2685 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1263_1_Left_2686 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1264_1_Left_2687 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1265_1_Left_2688 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1266_1_Left_2689 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1267_1_Left_2690 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1268_1_Left_2691 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1269_1_Left_2692 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1270_1_Left_2693 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1271_1_Left_2694 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1272_1_Left_2695 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1273_1_Left_2696 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1274_1_Left_2697 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1275_1_Left_2698 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1276_1_Left_2699 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1277_1_Left_2700 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1278_1_Left_2701 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1279_1_Left_2702 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1280_1_Left_2703 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1281_1_Left_2704 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1282_1_Left_2705 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1283_1_Left_2706 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1284_1_Left_2707 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1285_1_Left_2708 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1286_1_Left_2709 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1287_1_Left_2710 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1288_1_Left_2711 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1289_1_Left_2712 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1290_1_Left_2713 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1291_1_Left_2714 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1292_1_Left_2715 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1293_1_Left_2716 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1294_1_Left_2717 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1295_1_Left_2718 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1296_1_Left_2719 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1297_1_Left_2720 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1298_1_Left_2721 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1299_1_Left_2722 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1300_1_Left_2723 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1301_1_Left_2724 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1302_1_Left_2725 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1303_1_Left_2726 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1304_1_Left_2727 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1305_1_Left_2728 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1306_1_Left_2729 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1307_1_Left_2730 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1308_1_Left_2731 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1309_1_Left_2732 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1310_1_Left_2733 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1311_1_Left_2734 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1312_1_Left_2735 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1313_1_Left_2736 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1314_1_Left_2737 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1315_1_Left_2738 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1316_1_Left_2739 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1317_1_Left_2740 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1318_1_Left_2741 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1319_1_Left_2742 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1320_1_Left_2743 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1321_1_Left_2744 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1322_1_Left_2745 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1323_1_Left_2746 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1324_1_Left_2747 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1325_1_Left_2748 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1326_1_Left_2749 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1327_1_Left_2750 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1328_1_Left_2751 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1329_1_Left_2752 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1330_1_Left_2753 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1331_1_Left_2754 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1332_1_Left_2755 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1333_1_Left_2756 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1334_1_Left_2757 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1335_1_Left_2758 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1336_1_Left_2759 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1337_1_Left_2760 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1338_1_Left_2761 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1339_1_Left_2762 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1340_1_Left_2763 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1341_1_Left_2764 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1342_1_Left_2765 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1343_1_Left_2766 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1344_1_Left_2767 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1345_1_Left_2768 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1346_1_Left_2769 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1347_1_Left_2770 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1348_1_Left_2771 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1349_1_Left_2772 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1350_1_Left_2773 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1351_1_Left_2774 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1352_1_Left_2775 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1353_1_Left_2776 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1354_1_Left_2777 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1355_1_Left_2778 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1356_1_Left_2779 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1357_1_Left_2780 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1358_1_Left_2781 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1359_1_Left_2782 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1360_1_Left_2783 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1361_1_Left_2784 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1362_1_Left_2785 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1363_1_Left_2786 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1364_1_Left_2787 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1365_1_Left_2788 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1366_1_Left_2789 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1367_1_Left_2790 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1368_1_Left_2791 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1369_1_Left_2792 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1370_1_Left_2793 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1371_1_Left_2794 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1372_1_Left_2795 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1373_1_Left_2796 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1374_1_Left_2797 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1375_1_Left_2798 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1376_1_Left_2799 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1377_1_Left_2800 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1378_1_Left_2801 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1379_1_Left_2802 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1380_1_Left_2803 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1381_1_Left_2804 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1382_1_Left_2805 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1383_1_Left_2806 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1384_1_Left_2807 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1385_1_Left_2808 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1386_1_Left_2809 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1387_1_Left_2810 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1388_1_Left_2811 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1389_1_Left_2812 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1390_1_Left_2813 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1391_1_Left_2814 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1392_1_Left_2815 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1393_1_Left_2816 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1394_1_Left_2817 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1395_1_Left_2818 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1396_1_Left_2819 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1397_1_Left_2820 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1398_1_Left_2821 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1399_1_Left_2822 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1400_1_Left_2823 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1401_1_Left_2824 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1402_1_Left_2825 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1403_1_Left_2826 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1404_1_Left_2827 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1405_1_Left_2828 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1406_1_Left_2829 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1407_1_Left_2830 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1408_1_Left_2831 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1409_1_Left_2832 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1410_Left_2833 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1411_Left_2834 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1412_Left_2835 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1413_Left_2836 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1414_Left_2837 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1415_Left_2838 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1416_Left_2839 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1417_Left_2840 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1418_Left_2841 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1419_Left_2842 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1420_Left_2843 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1421_Left_2844 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1422_Left_2845 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1423_Left_2846 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_1_Left_2847 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_9_Left_2848 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_9_Left_2849 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_9_Left_2850 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_9_Left_2851 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_9_Left_2852 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_9_Left_2853 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_9_Left_2854 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_9_Left_2855 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_9_Left_2856 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_9_Left_2857 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_9_Left_2858 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_9_Left_2859 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_9_Left_2860 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_9_Left_2861 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_9_Left_2862 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_9_Left_2863 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_9_Left_2864 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_9_Left_2865 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_9_Left_2866 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_9_Left_2867 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_9_Left_2868 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_9_Left_2869 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_9_Left_2870 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_9_Left_2871 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_9_Left_2872 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_9_Left_2873 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_9_Left_2874 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_9_Left_2875 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_9_Left_2876 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_9_Left_2877 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_9_Left_2878 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_9_Left_2879 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_9_Left_2880 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_9_Left_2881 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_9_Left_2882 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_9_Left_2883 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_9_Left_2884 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_9_Left_2885 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_9_Left_2886 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_9_Left_2887 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_9_Left_2888 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_9_Left_2889 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_9_Left_2890 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_9_Left_2891 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_9_Left_2892 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_9_Left_2893 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_9_Left_2894 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_9_Left_2895 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_9_Left_2896 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_9_Left_2897 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_9_Left_2898 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_9_Left_2899 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_9_Left_2900 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_9_Left_2901 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_9_Left_2902 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_9_Left_2903 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_9_Left_2904 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_9_Left_2905 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_9_Left_2906 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_9_Left_2907 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_9_Left_2908 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_9_Left_2909 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_9_Left_2910 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_9_Left_2911 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_9_Left_2912 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_9_Left_2913 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_9_Left_2914 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_9_Left_2915 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_9_Left_2916 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_9_Left_2917 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_9_Left_2918 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_9_Left_2919 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_9_Left_2920 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_9_Left_2921 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_9_Left_2922 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_9_Left_2923 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_9_Left_2924 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_9_Left_2925 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_9_Left_2926 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_9_Left_2927 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_9_Left_2928 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_9_Left_2929 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_9_Left_2930 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_9_Left_2931 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_9_Left_2932 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_9_Left_2933 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_9_Left_2934 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_9_Left_2935 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_9_Left_2936 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_9_Left_2937 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_9_Left_2938 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_9_Left_2939 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_9_Left_2940 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_9_Left_2941 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_9_Left_2942 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_9_Left_2943 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_9_Left_2944 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_9_Left_2945 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_9_Left_2946 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_9_Left_2947 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_9_Left_2948 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_9_Left_2949 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_9_Left_2950 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_9_Left_2951 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_9_Left_2952 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_9_Left_2953 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_9_Left_2954 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_9_Left_2955 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_9_Left_2956 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_9_Left_2957 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_9_Left_2958 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_9_Left_2959 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_9_Left_2960 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_9_Left_2961 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_9_Left_2962 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_9_Left_2963 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_9_Left_2964 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_9_Left_2965 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_9_Left_2966 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_9_Left_2967 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_9_Left_2968 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_9_Left_2969 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_9_Left_2970 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_9_Left_2971 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_9_Left_2972 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_9_Left_2973 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_9_Left_2974 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_9_Left_2975 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_9_Left_2976 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_9_Left_2977 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_9_Left_2978 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_9_Left_2979 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_9_Left_2980 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_9_Left_2981 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_9_Left_2982 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_9_Left_2983 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_9_Left_2984 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_9_Left_2985 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_9_Left_2986 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_9_Left_2987 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_9_Left_2988 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_9_Left_2989 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_9_Left_2990 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_9_Left_2991 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_9_Left_2992 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_9_Left_2993 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_9_Left_2994 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_9_Left_2995 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_9_Left_2996 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_9_Left_2997 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_9_Left_2998 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_9_Left_2999 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_9_Left_3000 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_9_Left_3001 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_9_Left_3002 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_9_Left_3003 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_9_Left_3004 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_9_Left_3005 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_9_Left_3006 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_9_Left_3007 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_9_Left_3008 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_9_Left_3009 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_9_Left_3010 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_9_Left_3011 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_1_Right_3012 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_1_Right_3013 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_1_Right_3014 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_1_Right_3015 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_1_Right_3016 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_1_Right_3017 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_1_Right_3018 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_1_Right_3019 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_1_Right_3020 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_1_Right_3021 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_1_Right_3022 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_1_Right_3023 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_1_Right_3024 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_1_Right_3025 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_1_Right_3026 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_1_Right_3027 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_1_Right_3028 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_1_Right_3029 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_1_Right_3030 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_1_Right_3031 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_1_Right_3032 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_1_Right_3033 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_1_Right_3034 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_1_Right_3035 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_1_Right_3036 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_1_Right_3037 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_1_Right_3038 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_1_Right_3039 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_1_Right_3040 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_1_Right_3041 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_1_Right_3042 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_1_Right_3043 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_1_Right_3044 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_1_Right_3045 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_1_Right_3046 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_1_Right_3047 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_1_Right_3048 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_1_Right_3049 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_1_Right_3050 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_1_Right_3051 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_1_Right_3052 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_1_Right_3053 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_1_Right_3054 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_1_Right_3055 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_1_Right_3056 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_1_Right_3057 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_1_Right_3058 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_1_Right_3059 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_1_Right_3060 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_1_Right_3061 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_1_Right_3062 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_1_Right_3063 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_1_Right_3064 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_1_Right_3065 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_1_Right_3066 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_1_Right_3067 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_1_Right_3068 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_1_Right_3069 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_1_Right_3070 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_1_Right_3071 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_1_Right_3072 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_1_Right_3073 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_1_Right_3074 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_1_Right_3075 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_1_Right_3076 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_1_Right_3077 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_1_Right_3078 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_1_Right_3079 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_1_Right_3080 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_1_Right_3081 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_1_Right_3082 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_1_Right_3083 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_1_Right_3084 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_1_Right_3085 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_1_Right_3086 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_1_Right_3087 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_1_Right_3088 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_1_Right_3089 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_1_Right_3090 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_1_Right_3091 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_1_Right_3092 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_1_Right_3093 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_1_Right_3094 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_1_Right_3095 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_1_Right_3096 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_1_Right_3097 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_1_Right_3098 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_1_Right_3099 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_1_Right_3100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_1_Right_3101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_1_Right_3102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_1_Right_3103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_1_Right_3104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_1_Right_3105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_1_Right_3106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_1_Right_3107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_1_Right_3108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_1_Right_3109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_1_Right_3110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_1_Right_3111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_1_Right_3112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_1_Right_3113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_1_Right_3114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_1_Right_3115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_1_Right_3116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_1_Right_3117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_1_Right_3118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_1_Right_3119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_1_Right_3120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_1_Right_3121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_1_Right_3122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_1_Right_3123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_1_Right_3124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_1_Right_3125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_1_Right_3126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_1_Right_3127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_1_Right_3128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_1_Right_3129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_1_Right_3130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_1_Right_3131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_1_Right_3132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_1_Right_3133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_1_Right_3134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_1_Right_3135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_1_Right_3136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_1_Right_3137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_1_Right_3138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_1_Right_3139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_1_Right_3140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_1_Right_3141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_1_Right_3142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_1_Right_3143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_1_Right_3144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_1_Right_3145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_1_Right_3146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_1_Right_3147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_1_Right_3148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_152_1_Right_3149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_153_1_Right_3150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_154_1_Right_3151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_155_1_Right_3152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_156_1_Right_3153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_157_1_Right_3154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_158_1_Right_3155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_159_1_Right_3156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_160_1_Right_3157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_161_1_Right_3158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_162_1_Right_3159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_163_1_Right_3160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_164_1_Right_3161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_165_1_Right_3162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_166_1_Right_3163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_167_1_Right_3164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_168_1_Right_3165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_169_1_Right_3166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_170_1_Right_3167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_171_1_Right_3168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_172_1_Right_3169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_173_1_Right_3170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_174_1_Right_3171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_175_1_Right_3172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_176_1_Right_3173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_177_1_Right_3174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_1_Right_3175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_9_Left_3176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_9_Left_3177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_9_Left_3178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_9_Left_3179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_9_Left_3180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_9_Left_3181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_9_Left_3182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_9_Left_3183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_9_Left_3184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_9_Left_3185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_9_Left_3186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_9_Left_3187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_9_Left_3188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_9_Left_3189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_9_Left_3190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_9_Left_3191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_9_Left_3192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_9_Left_3193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_9_Left_3194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_9_Left_3195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_9_Left_3196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_9_Left_3197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_9_Left_3198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_9_Left_3199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_9_Left_3200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_9_Left_3201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_9_Left_3202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_9_Left_3203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_9_Left_3204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_9_Left_3205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_9_Left_3206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_9_Left_3207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_9_Left_3208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_9_Left_3209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_9_Left_3210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_9_Left_3211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_9_Left_3212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_9_Left_3213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_9_Left_3214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_9_Left_3215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_9_Left_3216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_9_Left_3217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_9_Left_3218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_9_Left_3219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_9_Left_3220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_9_Left_3221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_9_Left_3222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_9_Left_3223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_9_Left_3224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_9_Left_3225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_9_Left_3226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_9_Left_3227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_9_Left_3228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_9_Left_3229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_9_Left_3230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_9_Left_3231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_9_Left_3232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_9_Left_3233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_9_Left_3234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_9_Left_3235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_9_Left_3236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_9_Left_3237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_9_Left_3238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_9_Left_3239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_9_Left_3240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_9_Left_3241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_9_Left_3242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_9_Left_3243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_9_Left_3244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_9_Left_3245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_9_Left_3246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_9_Left_3247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_9_Left_3248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_9_Left_3249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_9_Left_3250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_9_Left_3251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_9_Left_3252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_9_Left_3253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_9_Left_3254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_9_Left_3255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_9_Left_3256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_9_Left_3257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_9_Left_3258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_9_Left_3259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_9_Left_3260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_9_Left_3261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_9_Left_3262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_9_Left_3263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_9_Left_3264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_9_Left_3265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_9_Left_3266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_9_Left_3267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_9_Left_3268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_9_Left_3269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_9_Left_3270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_9_Left_3271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_9_Left_3272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_9_Left_3273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_9_Left_3274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_9_Left_3275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_9_Left_3276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_9_Left_3277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_9_Left_3278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_9_Left_3279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_9_Left_3280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_295_9_Left_3281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_296_9_Left_3282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_297_9_Left_3283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_298_9_Left_3284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_299_9_Left_3285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_300_9_Left_3286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_301_9_Left_3287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_302_9_Left_3288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_303_9_Left_3289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_304_9_Left_3290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_305_9_Left_3291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_306_9_Left_3292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_307_9_Left_3293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_308_9_Left_3294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_309_9_Left_3295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_310_9_Left_3296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_311_9_Left_3297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_312_9_Left_3298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_313_9_Left_3299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_314_9_Left_3300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_315_9_Left_3301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_316_9_Left_3302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_317_9_Left_3303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_318_9_Left_3304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_319_9_Left_3305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_320_9_Left_3306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_321_9_Left_3307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_322_9_Left_3308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_323_9_Left_3309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_324_9_Left_3310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_325_9_Left_3311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_326_9_Left_3312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_327_9_Left_3313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_328_9_Left_3314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_329_9_Left_3315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_330_9_Left_3316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_331_9_Left_3317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_332_9_Left_3318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_333_9_Left_3319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_334_9_Left_3320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_335_9_Left_3321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_336_9_Left_3322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_337_9_Left_3323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_338_9_Left_3324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_339_9_Left_3325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_340_9_Left_3326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_341_9_Left_3327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_342_9_Left_3328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_343_9_Left_3329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_344_9_Left_3330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_345_9_Left_3331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_346_9_Left_3332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_347_9_Left_3333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_348_9_Left_3334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_349_9_Left_3335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_350_9_Left_3336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_351_9_Left_3337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_352_9_Left_3338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_353_9_Left_3339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_190_1_Right_3340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_191_1_Right_3341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_192_1_Right_3342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_193_1_Right_3343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_194_1_Right_3344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_195_1_Right_3345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_196_1_Right_3346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_197_1_Right_3347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_198_1_Right_3348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_199_1_Right_3349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_200_1_Right_3350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_201_1_Right_3351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_202_1_Right_3352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_203_1_Right_3353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_204_1_Right_3354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_205_1_Right_3355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_206_1_Right_3356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_207_1_Right_3357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_208_1_Right_3358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_209_1_Right_3359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_210_1_Right_3360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_211_1_Right_3361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_212_1_Right_3362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_213_1_Right_3363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_214_1_Right_3364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_215_1_Right_3365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_216_1_Right_3366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_217_1_Right_3367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_218_1_Right_3368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_219_1_Right_3369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_220_1_Right_3370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_221_1_Right_3371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_222_1_Right_3372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_223_1_Right_3373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_224_1_Right_3374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_225_1_Right_3375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_226_1_Right_3376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_227_1_Right_3377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_228_1_Right_3378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_229_1_Right_3379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_230_1_Right_3380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_231_1_Right_3381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_232_1_Right_3382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_233_1_Right_3383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_234_1_Right_3384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_235_1_Right_3385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_236_1_Right_3386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_237_1_Right_3387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_238_1_Right_3388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_239_1_Right_3389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_240_1_Right_3390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_241_1_Right_3391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_242_1_Right_3392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_243_1_Right_3393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_244_1_Right_3394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_245_1_Right_3395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_246_1_Right_3396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_247_1_Right_3397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_248_1_Right_3398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_249_1_Right_3399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_250_1_Right_3400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_251_1_Right_3401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_252_1_Right_3402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_253_1_Right_3403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_254_1_Right_3404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_255_1_Right_3405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_256_1_Right_3406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_257_1_Right_3407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_258_1_Right_3408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_259_1_Right_3409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_260_1_Right_3410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_261_1_Right_3411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_262_1_Right_3412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_263_1_Right_3413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_264_1_Right_3414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_265_1_Right_3415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_266_1_Right_3416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_267_1_Right_3417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_268_1_Right_3418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_269_1_Right_3419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_270_1_Right_3420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_271_1_Right_3421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_272_1_Right_3422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_273_1_Right_3423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_274_1_Right_3424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_275_1_Right_3425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_276_1_Right_3426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_277_1_Right_3427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_278_1_Right_3428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_279_1_Right_3429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_280_1_Right_3430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_281_1_Right_3431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_282_1_Right_3432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_283_1_Right_3433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_284_1_Right_3434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_285_1_Right_3435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_286_1_Right_3436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_287_1_Right_3437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_288_1_Right_3438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_289_1_Right_3439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_290_1_Right_3440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_291_1_Right_3441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_292_1_Right_3442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_293_1_Right_3443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_294_1_Right_3444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_295_1_Right_3445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_296_1_Right_3446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_297_1_Right_3447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_298_1_Right_3448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_299_1_Right_3449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_300_1_Right_3450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_301_1_Right_3451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_302_1_Right_3452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_303_1_Right_3453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_304_1_Right_3454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_305_1_Right_3455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_306_1_Right_3456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_307_1_Right_3457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_308_1_Right_3458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_309_1_Right_3459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_310_1_Right_3460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_311_1_Right_3461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_312_1_Right_3462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_313_1_Right_3463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_314_1_Right_3464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_315_1_Right_3465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_316_1_Right_3466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_317_1_Right_3467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_318_1_Right_3468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_319_1_Right_3469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_320_1_Right_3470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_321_1_Right_3471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_322_1_Right_3472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_323_1_Right_3473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_324_1_Right_3474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_325_1_Right_3475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_326_1_Right_3476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_327_1_Right_3477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_328_1_Right_3478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_329_1_Right_3479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_330_1_Right_3480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_331_1_Right_3481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_332_1_Right_3482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_333_1_Right_3483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_334_1_Right_3484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_335_1_Right_3485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_336_1_Right_3486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_337_1_Right_3487 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_338_1_Right_3488 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_339_1_Right_3489 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_340_1_Right_3490 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_341_1_Right_3491 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_342_1_Right_3492 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_343_1_Right_3493 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_344_1_Right_3494 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_345_1_Right_3495 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_346_1_Right_3496 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_347_1_Right_3497 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_348_1_Right_3498 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_349_1_Right_3499 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_350_1_Right_3500 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_351_1_Right_3501 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_352_1_Right_3502 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_353_1_Right_3503 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_366_9_Left_3504 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_367_9_Left_3505 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_368_9_Left_3506 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_369_9_Left_3507 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_370_9_Left_3508 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_371_9_Left_3509 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_372_9_Left_3510 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_373_9_Left_3511 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_374_9_Left_3512 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_375_9_Left_3513 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_376_9_Left_3514 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_377_9_Left_3515 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_378_9_Left_3516 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_379_9_Left_3517 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_380_9_Left_3518 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_381_9_Left_3519 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_382_9_Left_3520 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_383_9_Left_3521 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_384_9_Left_3522 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_385_9_Left_3523 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_386_9_Left_3524 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_387_9_Left_3525 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_388_9_Left_3526 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_389_9_Left_3527 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_390_9_Left_3528 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_391_9_Left_3529 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_392_9_Left_3530 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_393_9_Left_3531 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_394_9_Left_3532 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_395_9_Left_3533 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_396_9_Left_3534 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_397_9_Left_3535 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_398_9_Left_3536 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_399_9_Left_3537 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_400_9_Left_3538 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_401_9_Left_3539 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_402_9_Left_3540 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_403_9_Left_3541 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_404_9_Left_3542 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_405_9_Left_3543 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_406_9_Left_3544 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_407_9_Left_3545 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_408_9_Left_3546 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_409_9_Left_3547 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_410_9_Left_3548 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_411_9_Left_3549 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_412_9_Left_3550 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_413_9_Left_3551 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_414_9_Left_3552 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_415_9_Left_3553 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_416_9_Left_3554 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_417_9_Left_3555 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_418_9_Left_3556 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_419_9_Left_3557 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_420_9_Left_3558 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_421_9_Left_3559 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_422_9_Left_3560 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_423_9_Left_3561 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_424_9_Left_3562 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_425_9_Left_3563 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_426_9_Left_3564 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_427_9_Left_3565 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_428_9_Left_3566 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_429_9_Left_3567 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_430_9_Left_3568 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_431_9_Left_3569 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_432_9_Left_3570 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_433_9_Left_3571 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_434_9_Left_3572 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_435_9_Left_3573 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_436_9_Left_3574 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_437_9_Left_3575 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_438_9_Left_3576 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_439_9_Left_3577 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_440_9_Left_3578 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_441_9_Left_3579 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_442_9_Left_3580 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_443_9_Left_3581 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_444_9_Left_3582 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_445_9_Left_3583 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_446_9_Left_3584 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_447_9_Left_3585 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_448_9_Left_3586 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_449_9_Left_3587 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_450_9_Left_3588 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_451_9_Left_3589 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_452_9_Left_3590 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_453_9_Left_3591 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_454_9_Left_3592 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_455_9_Left_3593 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_456_9_Left_3594 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_457_9_Left_3595 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_458_9_Left_3596 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_459_9_Left_3597 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_460_9_Left_3598 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_461_9_Left_3599 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_462_9_Left_3600 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_463_9_Left_3601 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_464_9_Left_3602 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_465_9_Left_3603 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_466_9_Left_3604 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_467_9_Left_3605 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_468_9_Left_3606 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_469_9_Left_3607 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_470_9_Left_3608 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_471_9_Left_3609 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_472_9_Left_3610 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_473_9_Left_3611 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_474_9_Left_3612 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_475_9_Left_3613 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_476_9_Left_3614 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_477_9_Left_3615 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_478_9_Left_3616 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_479_9_Left_3617 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_480_9_Left_3618 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_481_9_Left_3619 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_482_9_Left_3620 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_483_9_Left_3621 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_484_9_Left_3622 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_485_9_Left_3623 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_486_9_Left_3624 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_487_9_Left_3625 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_488_9_Left_3626 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_489_9_Left_3627 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_490_9_Left_3628 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_491_9_Left_3629 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_492_9_Left_3630 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_493_9_Left_3631 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_494_9_Left_3632 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_495_9_Left_3633 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_496_9_Left_3634 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_497_9_Left_3635 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_498_9_Left_3636 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_499_9_Left_3637 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_500_9_Left_3638 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_501_9_Left_3639 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_502_9_Left_3640 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_503_9_Left_3641 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_504_9_Left_3642 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_505_9_Left_3643 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_506_9_Left_3644 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_507_9_Left_3645 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_508_9_Left_3646 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_509_9_Left_3647 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_510_9_Left_3648 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_511_9_Left_3649 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_512_9_Left_3650 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_513_9_Left_3651 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_514_9_Left_3652 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_515_9_Left_3653 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_516_9_Left_3654 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_517_9_Left_3655 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_518_9_Left_3656 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_519_9_Left_3657 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_520_9_Left_3658 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_521_9_Left_3659 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_522_9_Left_3660 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_523_9_Left_3661 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_524_9_Left_3662 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_525_9_Left_3663 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_526_9_Left_3664 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_527_9_Left_3665 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_528_9_Left_3666 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_529_9_Left_3667 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_366_1_Right_3668 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_367_1_Right_3669 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_368_1_Right_3670 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_369_1_Right_3671 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_370_1_Right_3672 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_371_1_Right_3673 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_372_1_Right_3674 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_373_1_Right_3675 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_374_1_Right_3676 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_375_1_Right_3677 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_376_1_Right_3678 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_377_1_Right_3679 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_378_1_Right_3680 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_379_1_Right_3681 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_380_1_Right_3682 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_381_1_Right_3683 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_382_1_Right_3684 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_383_1_Right_3685 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_384_1_Right_3686 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_385_1_Right_3687 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_386_1_Right_3688 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_387_1_Right_3689 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_388_1_Right_3690 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_389_1_Right_3691 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_390_1_Right_3692 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_391_1_Right_3693 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_392_1_Right_3694 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_393_1_Right_3695 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_394_1_Right_3696 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_395_1_Right_3697 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_396_1_Right_3698 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_397_1_Right_3699 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_398_1_Right_3700 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_399_1_Right_3701 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_400_1_Right_3702 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_401_1_Right_3703 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_402_1_Right_3704 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_403_1_Right_3705 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_404_1_Right_3706 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_405_1_Right_3707 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_406_1_Right_3708 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_407_1_Right_3709 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_408_1_Right_3710 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_409_1_Right_3711 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_410_1_Right_3712 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_411_1_Right_3713 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_412_1_Right_3714 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_413_1_Right_3715 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_414_1_Right_3716 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_415_1_Right_3717 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_416_1_Right_3718 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_417_1_Right_3719 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_418_1_Right_3720 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_419_1_Right_3721 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_420_1_Right_3722 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_421_1_Right_3723 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_422_1_Right_3724 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_423_1_Right_3725 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_424_1_Right_3726 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_425_1_Right_3727 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_426_1_Right_3728 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_427_1_Right_3729 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_428_1_Right_3730 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_429_1_Right_3731 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_430_1_Right_3732 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_431_1_Right_3733 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_432_1_Right_3734 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_433_1_Right_3735 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_434_1_Right_3736 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_435_1_Right_3737 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_436_1_Right_3738 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_437_1_Right_3739 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_438_1_Right_3740 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_439_1_Right_3741 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_440_1_Right_3742 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_441_1_Right_3743 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_442_1_Right_3744 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_443_1_Right_3745 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_444_1_Right_3746 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_445_1_Right_3747 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_446_1_Right_3748 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_447_1_Right_3749 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_448_1_Right_3750 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_449_1_Right_3751 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_450_1_Right_3752 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_451_1_Right_3753 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_452_1_Right_3754 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_453_1_Right_3755 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_454_1_Right_3756 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_455_1_Right_3757 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_456_1_Right_3758 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_457_1_Right_3759 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_458_1_Right_3760 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_459_1_Right_3761 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_460_1_Right_3762 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_461_1_Right_3763 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_462_1_Right_3764 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_463_1_Right_3765 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_464_1_Right_3766 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_465_1_Right_3767 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_466_1_Right_3768 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_467_1_Right_3769 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_468_1_Right_3770 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_469_1_Right_3771 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_470_1_Right_3772 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_471_1_Right_3773 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_472_1_Right_3774 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_473_1_Right_3775 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_474_1_Right_3776 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_475_1_Right_3777 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_476_1_Right_3778 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_477_1_Right_3779 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_478_1_Right_3780 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_479_1_Right_3781 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_480_1_Right_3782 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_481_1_Right_3783 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_482_1_Right_3784 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_483_1_Right_3785 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_484_1_Right_3786 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_485_1_Right_3787 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_486_1_Right_3788 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_487_1_Right_3789 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_488_1_Right_3790 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_489_1_Right_3791 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_490_1_Right_3792 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_491_1_Right_3793 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_492_1_Right_3794 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_493_1_Right_3795 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_494_1_Right_3796 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_495_1_Right_3797 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_496_1_Right_3798 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_497_1_Right_3799 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_498_1_Right_3800 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_499_1_Right_3801 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_500_1_Right_3802 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_501_1_Right_3803 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_502_1_Right_3804 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_503_1_Right_3805 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_504_1_Right_3806 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_505_1_Right_3807 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_506_1_Right_3808 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_507_1_Right_3809 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_508_1_Right_3810 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_509_1_Right_3811 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_510_1_Right_3812 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_511_1_Right_3813 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_512_1_Right_3814 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_513_1_Right_3815 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_514_1_Right_3816 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_515_1_Right_3817 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_516_1_Right_3818 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_517_1_Right_3819 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_518_1_Right_3820 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_519_1_Right_3821 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_520_1_Right_3822 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_521_1_Right_3823 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_522_1_Right_3824 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_523_1_Right_3825 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_524_1_Right_3826 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_525_1_Right_3827 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_526_1_Right_3828 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_527_1_Right_3829 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_528_1_Right_3830 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_529_1_Right_3831 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_542_9_Left_3832 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_543_9_Left_3833 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_544_9_Left_3834 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_545_9_Left_3835 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_546_9_Left_3836 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_547_9_Left_3837 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_548_9_Left_3838 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_549_9_Left_3839 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_550_9_Left_3840 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_551_9_Left_3841 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_552_9_Left_3842 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_553_9_Left_3843 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_554_9_Left_3844 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_555_9_Left_3845 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_556_9_Left_3846 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_557_9_Left_3847 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_558_9_Left_3848 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_559_9_Left_3849 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_560_9_Left_3850 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_561_9_Left_3851 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_562_9_Left_3852 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_563_9_Left_3853 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_564_9_Left_3854 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_565_9_Left_3855 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_566_9_Left_3856 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_567_9_Left_3857 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_568_9_Left_3858 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_569_9_Left_3859 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_570_9_Left_3860 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_571_9_Left_3861 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_572_9_Left_3862 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_573_9_Left_3863 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_574_9_Left_3864 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_575_9_Left_3865 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_576_9_Left_3866 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_577_9_Left_3867 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_578_9_Left_3868 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_579_9_Left_3869 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_580_9_Left_3870 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_581_9_Left_3871 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_582_9_Left_3872 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_583_9_Left_3873 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_584_9_Left_3874 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_585_9_Left_3875 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_586_9_Left_3876 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_587_9_Left_3877 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_588_9_Left_3878 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_589_9_Left_3879 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_590_9_Left_3880 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_591_9_Left_3881 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_592_9_Left_3882 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_593_9_Left_3883 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_594_9_Left_3884 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_595_9_Left_3885 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_596_9_Left_3886 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_597_9_Left_3887 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_598_9_Left_3888 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_599_9_Left_3889 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_600_9_Left_3890 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_601_9_Left_3891 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_602_9_Left_3892 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_603_9_Left_3893 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_604_9_Left_3894 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_605_9_Left_3895 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_606_9_Left_3896 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_607_9_Left_3897 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_608_9_Left_3898 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_609_9_Left_3899 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_610_9_Left_3900 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_611_9_Left_3901 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_612_9_Left_3902 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_613_9_Left_3903 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_614_9_Left_3904 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_615_9_Left_3905 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_616_9_Left_3906 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_617_9_Left_3907 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_618_9_Left_3908 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_619_9_Left_3909 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_620_9_Left_3910 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_621_9_Left_3911 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_622_9_Left_3912 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_623_9_Left_3913 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_624_9_Left_3914 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_625_9_Left_3915 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_626_9_Left_3916 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_627_9_Left_3917 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_628_9_Left_3918 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_629_9_Left_3919 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_630_9_Left_3920 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_631_9_Left_3921 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_632_9_Left_3922 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_633_9_Left_3923 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_634_9_Left_3924 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_635_9_Left_3925 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_636_9_Left_3926 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_637_9_Left_3927 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_638_9_Left_3928 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_639_9_Left_3929 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_640_9_Left_3930 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_641_9_Left_3931 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_642_9_Left_3932 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_643_9_Left_3933 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_644_9_Left_3934 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_645_9_Left_3935 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_646_9_Left_3936 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_647_9_Left_3937 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_648_9_Left_3938 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_649_9_Left_3939 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_650_9_Left_3940 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_651_9_Left_3941 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_652_9_Left_3942 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_653_9_Left_3943 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_654_9_Left_3944 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_655_9_Left_3945 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_656_9_Left_3946 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_657_9_Left_3947 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_658_9_Left_3948 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_659_9_Left_3949 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_660_9_Left_3950 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_661_9_Left_3951 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_662_9_Left_3952 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_663_9_Left_3953 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_664_9_Left_3954 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_665_9_Left_3955 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_666_9_Left_3956 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_667_9_Left_3957 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_668_9_Left_3958 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_669_9_Left_3959 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_670_9_Left_3960 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_671_9_Left_3961 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_672_9_Left_3962 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_673_9_Left_3963 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_674_9_Left_3964 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_675_9_Left_3965 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_676_9_Left_3966 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_677_9_Left_3967 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_678_9_Left_3968 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_679_9_Left_3969 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_680_9_Left_3970 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_681_9_Left_3971 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_682_9_Left_3972 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_683_9_Left_3973 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_684_9_Left_3974 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_685_9_Left_3975 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_686_9_Left_3976 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_687_9_Left_3977 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_688_9_Left_3978 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_689_9_Left_3979 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_690_9_Left_3980 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_691_9_Left_3981 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_692_9_Left_3982 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_693_9_Left_3983 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_694_9_Left_3984 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_695_9_Left_3985 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_696_9_Left_3986 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_697_9_Left_3987 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_698_9_Left_3988 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_699_9_Left_3989 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_700_9_Left_3990 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_701_9_Left_3991 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_702_9_Left_3992 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_703_9_Left_3993 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_704_9_Left_3994 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_705_9_Left_3995 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_542_1_Right_3996 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_543_1_Right_3997 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_544_1_Right_3998 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_545_1_Right_3999 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_546_1_Right_4000 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_547_1_Right_4001 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_548_1_Right_4002 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_549_1_Right_4003 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_550_1_Right_4004 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_551_1_Right_4005 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_552_1_Right_4006 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_553_1_Right_4007 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_554_1_Right_4008 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_555_1_Right_4009 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_556_1_Right_4010 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_557_1_Right_4011 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_558_1_Right_4012 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_559_1_Right_4013 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_560_1_Right_4014 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_561_1_Right_4015 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_562_1_Right_4016 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_563_1_Right_4017 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_564_1_Right_4018 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_565_1_Right_4019 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_566_1_Right_4020 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_567_1_Right_4021 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_568_1_Right_4022 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_569_1_Right_4023 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_570_1_Right_4024 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_571_1_Right_4025 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_572_1_Right_4026 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_573_1_Right_4027 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_574_1_Right_4028 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_575_1_Right_4029 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_576_1_Right_4030 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_577_1_Right_4031 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_578_1_Right_4032 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_579_1_Right_4033 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_580_1_Right_4034 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_581_1_Right_4035 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_582_1_Right_4036 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_583_1_Right_4037 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_584_1_Right_4038 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_585_1_Right_4039 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_586_1_Right_4040 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_587_1_Right_4041 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_588_1_Right_4042 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_589_1_Right_4043 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_590_1_Right_4044 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_591_1_Right_4045 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_592_1_Right_4046 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_593_1_Right_4047 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_594_1_Right_4048 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_595_1_Right_4049 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_596_1_Right_4050 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_597_1_Right_4051 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_598_1_Right_4052 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_599_1_Right_4053 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_600_1_Right_4054 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_601_1_Right_4055 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_602_1_Right_4056 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_603_1_Right_4057 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_604_1_Right_4058 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_605_1_Right_4059 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_606_1_Right_4060 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_607_1_Right_4061 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_608_1_Right_4062 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_609_1_Right_4063 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_610_1_Right_4064 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_611_1_Right_4065 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_612_1_Right_4066 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_613_1_Right_4067 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_614_1_Right_4068 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_615_1_Right_4069 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_616_1_Right_4070 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_617_1_Right_4071 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_618_1_Right_4072 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_619_1_Right_4073 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_620_1_Right_4074 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_621_1_Right_4075 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_622_1_Right_4076 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_623_1_Right_4077 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_624_1_Right_4078 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_625_1_Right_4079 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_626_1_Right_4080 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_627_1_Right_4081 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_628_1_Right_4082 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_629_1_Right_4083 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_630_1_Right_4084 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_631_1_Right_4085 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_632_1_Right_4086 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_633_1_Right_4087 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_634_1_Right_4088 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_635_1_Right_4089 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_636_1_Right_4090 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_637_1_Right_4091 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_638_1_Right_4092 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_639_1_Right_4093 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_640_1_Right_4094 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_641_1_Right_4095 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_642_1_Right_4096 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_643_1_Right_4097 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_644_1_Right_4098 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_645_1_Right_4099 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_646_1_Right_4100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_647_1_Right_4101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_648_1_Right_4102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_649_1_Right_4103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_650_1_Right_4104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_651_1_Right_4105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_652_1_Right_4106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_653_1_Right_4107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_654_1_Right_4108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_655_1_Right_4109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_656_1_Right_4110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_657_1_Right_4111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_658_1_Right_4112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_659_1_Right_4113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_660_1_Right_4114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_661_1_Right_4115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_662_1_Right_4116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_663_1_Right_4117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_664_1_Right_4118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_665_1_Right_4119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_666_1_Right_4120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_667_1_Right_4121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_668_1_Right_4122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_669_1_Right_4123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_670_1_Right_4124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_671_1_Right_4125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_672_1_Right_4126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_673_1_Right_4127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_674_1_Right_4128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_675_1_Right_4129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_676_1_Right_4130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_677_1_Right_4131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_678_1_Right_4132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_679_1_Right_4133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_680_1_Right_4134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_681_1_Right_4135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_682_1_Right_4136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_683_1_Right_4137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_684_1_Right_4138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_685_1_Right_4139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_686_1_Right_4140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_687_1_Right_4141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_688_1_Right_4142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_689_1_Right_4143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_690_1_Right_4144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_691_1_Right_4145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_692_1_Right_4146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_693_1_Right_4147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_694_1_Right_4148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_695_1_Right_4149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_696_1_Right_4150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_697_1_Right_4151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_698_1_Right_4152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_699_1_Right_4153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_700_1_Right_4154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_701_1_Right_4155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_702_1_Right_4156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_703_1_Right_4157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_704_1_Right_4158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_705_1_Right_4159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_718_9_Left_4160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_719_9_Left_4161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_720_9_Left_4162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_721_9_Left_4163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_722_9_Left_4164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_723_9_Left_4165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_724_9_Left_4166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_725_9_Left_4167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_726_9_Left_4168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_727_9_Left_4169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_728_9_Left_4170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_729_9_Left_4171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_730_9_Left_4172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_731_9_Left_4173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_732_9_Left_4174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_733_9_Left_4175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_734_9_Left_4176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_735_9_Left_4177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_736_9_Left_4178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_737_9_Left_4179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_738_9_Left_4180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_739_9_Left_4181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_740_9_Left_4182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_741_9_Left_4183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_742_9_Left_4184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_743_9_Left_4185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_744_9_Left_4186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_745_9_Left_4187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_746_9_Left_4188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_747_9_Left_4189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_748_9_Left_4190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_749_9_Left_4191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_750_9_Left_4192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_751_9_Left_4193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_752_9_Left_4194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_753_9_Left_4195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_754_9_Left_4196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_755_9_Left_4197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_756_9_Left_4198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_757_9_Left_4199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_758_9_Left_4200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_759_9_Left_4201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_760_9_Left_4202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_761_9_Left_4203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_762_9_Left_4204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_763_9_Left_4205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_764_9_Left_4206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_765_9_Left_4207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_766_9_Left_4208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_767_9_Left_4209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_768_9_Left_4210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_769_9_Left_4211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_770_9_Left_4212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_771_9_Left_4213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_772_9_Left_4214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_773_9_Left_4215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_774_9_Left_4216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_775_9_Left_4217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_776_9_Left_4218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_777_9_Left_4219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_778_9_Left_4220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_779_9_Left_4221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_780_9_Left_4222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_781_9_Left_4223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_782_9_Left_4224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_783_9_Left_4225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_784_9_Left_4226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_785_9_Left_4227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_786_9_Left_4228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_787_9_Left_4229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_788_9_Left_4230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_789_9_Left_4231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_790_9_Left_4232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_791_9_Left_4233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_792_9_Left_4234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_793_9_Left_4235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_794_9_Left_4236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_795_9_Left_4237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_796_9_Left_4238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_797_9_Left_4239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_798_9_Left_4240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_799_9_Left_4241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_800_9_Left_4242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_801_9_Left_4243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_802_9_Left_4244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_803_9_Left_4245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_804_9_Left_4246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_805_9_Left_4247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_806_9_Left_4248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_807_9_Left_4249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_808_9_Left_4250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_809_9_Left_4251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_810_9_Left_4252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_811_9_Left_4253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_812_9_Left_4254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_813_9_Left_4255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_814_9_Left_4256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_815_9_Left_4257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_816_9_Left_4258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_817_9_Left_4259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_818_9_Left_4260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_819_9_Left_4261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_820_9_Left_4262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_821_9_Left_4263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_822_9_Left_4264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_823_9_Left_4265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_824_9_Left_4266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_825_9_Left_4267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_826_9_Left_4268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_827_9_Left_4269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_828_9_Left_4270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_829_9_Left_4271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_830_9_Left_4272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_831_9_Left_4273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_832_9_Left_4274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_833_9_Left_4275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_834_9_Left_4276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_835_9_Left_4277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_836_9_Left_4278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_837_9_Left_4279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_838_9_Left_4280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_839_9_Left_4281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_840_9_Left_4282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_841_9_Left_4283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_842_9_Left_4284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_843_9_Left_4285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_844_9_Left_4286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_845_9_Left_4287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_846_9_Left_4288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_847_9_Left_4289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_848_9_Left_4290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_849_9_Left_4291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_850_9_Left_4292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_851_9_Left_4293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_852_9_Left_4294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_853_9_Left_4295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_854_9_Left_4296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_855_9_Left_4297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_856_9_Left_4298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_857_9_Left_4299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_858_9_Left_4300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_859_9_Left_4301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_860_9_Left_4302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_861_9_Left_4303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_862_9_Left_4304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_863_9_Left_4305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_864_9_Left_4306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_865_9_Left_4307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_866_9_Left_4308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_867_9_Left_4309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_868_9_Left_4310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_869_9_Left_4311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_870_9_Left_4312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_871_9_Left_4313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_872_9_Left_4314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_873_9_Left_4315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_874_9_Left_4316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_875_9_Left_4317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_876_9_Left_4318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_877_9_Left_4319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_878_9_Left_4320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_879_9_Left_4321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_880_9_Left_4322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_881_9_Left_4323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_718_1_Right_4324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_719_1_Right_4325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_720_1_Right_4326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_721_1_Right_4327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_722_1_Right_4328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_723_1_Right_4329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_724_1_Right_4330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_725_1_Right_4331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_726_1_Right_4332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_727_1_Right_4333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_728_1_Right_4334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_729_1_Right_4335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_730_1_Right_4336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_731_1_Right_4337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_732_1_Right_4338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_733_1_Right_4339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_734_1_Right_4340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_735_1_Right_4341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_736_1_Right_4342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_737_1_Right_4343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_738_1_Right_4344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_739_1_Right_4345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_740_1_Right_4346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_741_1_Right_4347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_742_1_Right_4348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_743_1_Right_4349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_744_1_Right_4350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_745_1_Right_4351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_746_1_Right_4352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_747_1_Right_4353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_748_1_Right_4354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_749_1_Right_4355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_750_1_Right_4356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_751_1_Right_4357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_752_1_Right_4358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_753_1_Right_4359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_754_1_Right_4360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_755_1_Right_4361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_756_1_Right_4362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_757_1_Right_4363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_758_1_Right_4364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_759_1_Right_4365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_760_1_Right_4366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_761_1_Right_4367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_762_1_Right_4368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_763_1_Right_4369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_764_1_Right_4370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_765_1_Right_4371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_766_1_Right_4372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_767_1_Right_4373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_768_1_Right_4374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_769_1_Right_4375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_770_1_Right_4376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_771_1_Right_4377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_772_1_Right_4378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_773_1_Right_4379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_774_1_Right_4380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_775_1_Right_4381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_776_1_Right_4382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_777_1_Right_4383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_778_1_Right_4384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_779_1_Right_4385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_780_1_Right_4386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_781_1_Right_4387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_782_1_Right_4388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_783_1_Right_4389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_784_1_Right_4390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_785_1_Right_4391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_786_1_Right_4392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_787_1_Right_4393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_788_1_Right_4394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_789_1_Right_4395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_790_1_Right_4396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_791_1_Right_4397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_792_1_Right_4398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_793_1_Right_4399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_794_1_Right_4400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_795_1_Right_4401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_796_1_Right_4402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_797_1_Right_4403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_798_1_Right_4404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_799_1_Right_4405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_800_1_Right_4406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_801_1_Right_4407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_802_1_Right_4408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_803_1_Right_4409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_804_1_Right_4410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_805_1_Right_4411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_806_1_Right_4412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_807_1_Right_4413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_808_1_Right_4414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_809_1_Right_4415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_810_1_Right_4416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_811_1_Right_4417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_812_1_Right_4418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_813_1_Right_4419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_814_1_Right_4420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_815_1_Right_4421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_816_1_Right_4422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_817_1_Right_4423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_818_1_Right_4424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_819_1_Right_4425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_820_1_Right_4426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_821_1_Right_4427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_822_1_Right_4428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_823_1_Right_4429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_824_1_Right_4430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_825_1_Right_4431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_826_1_Right_4432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_827_1_Right_4433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_828_1_Right_4434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_829_1_Right_4435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_830_1_Right_4436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_831_1_Right_4437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_832_1_Right_4438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_833_1_Right_4439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_834_1_Right_4440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_835_1_Right_4441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_836_1_Right_4442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_837_1_Right_4443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_838_1_Right_4444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_839_1_Right_4445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_840_1_Right_4446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_841_1_Right_4447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_842_1_Right_4448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_843_1_Right_4449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_844_1_Right_4450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_845_1_Right_4451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_846_1_Right_4452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_847_1_Right_4453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_848_1_Right_4454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_849_1_Right_4455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_850_1_Right_4456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_851_1_Right_4457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_852_1_Right_4458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_853_1_Right_4459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_854_1_Right_4460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_855_1_Right_4461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_856_1_Right_4462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_857_1_Right_4463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_858_1_Right_4464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_859_1_Right_4465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_860_1_Right_4466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_861_1_Right_4467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_862_1_Right_4468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_863_1_Right_4469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_864_1_Right_4470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_865_1_Right_4471 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_866_1_Right_4472 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_867_1_Right_4473 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_868_1_Right_4474 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_869_1_Right_4475 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_870_1_Right_4476 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_871_1_Right_4477 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_872_1_Right_4478 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_873_1_Right_4479 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_874_1_Right_4480 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_875_1_Right_4481 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_876_1_Right_4482 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_877_1_Right_4483 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_878_1_Right_4484 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_879_1_Right_4485 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_880_1_Right_4486 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_881_1_Right_4487 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_894_9_Left_4488 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_895_9_Left_4489 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_896_9_Left_4490 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_897_9_Left_4491 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_898_9_Left_4492 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_899_9_Left_4493 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_900_9_Left_4494 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_901_9_Left_4495 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_902_9_Left_4496 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_903_9_Left_4497 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_904_9_Left_4498 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_905_9_Left_4499 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_906_9_Left_4500 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_907_9_Left_4501 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_908_9_Left_4502 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_909_9_Left_4503 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_910_9_Left_4504 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_911_9_Left_4505 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_912_9_Left_4506 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_913_9_Left_4507 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_914_9_Left_4508 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_915_9_Left_4509 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_916_9_Left_4510 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_917_9_Left_4511 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_918_9_Left_4512 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_919_9_Left_4513 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_920_9_Left_4514 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_921_9_Left_4515 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_922_9_Left_4516 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_923_9_Left_4517 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_924_9_Left_4518 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_925_9_Left_4519 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_926_9_Left_4520 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_927_9_Left_4521 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_928_9_Left_4522 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_929_9_Left_4523 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_930_9_Left_4524 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_931_9_Left_4525 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_932_9_Left_4526 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_933_9_Left_4527 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_934_9_Left_4528 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_935_9_Left_4529 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_936_9_Left_4530 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_937_9_Left_4531 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_938_9_Left_4532 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_939_9_Left_4533 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_940_9_Left_4534 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_941_9_Left_4535 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_942_9_Left_4536 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_943_9_Left_4537 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_944_9_Left_4538 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_945_9_Left_4539 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_946_9_Left_4540 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_947_9_Left_4541 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_948_9_Left_4542 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_949_9_Left_4543 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_950_9_Left_4544 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_951_9_Left_4545 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_952_9_Left_4546 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_953_9_Left_4547 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_954_9_Left_4548 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_955_9_Left_4549 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_956_9_Left_4550 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_957_9_Left_4551 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_958_9_Left_4552 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_959_9_Left_4553 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_960_9_Left_4554 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_961_9_Left_4555 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_962_9_Left_4556 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_963_9_Left_4557 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_964_9_Left_4558 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_965_9_Left_4559 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_966_9_Left_4560 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_967_9_Left_4561 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_968_9_Left_4562 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_969_9_Left_4563 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_970_9_Left_4564 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_971_9_Left_4565 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_972_9_Left_4566 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_973_9_Left_4567 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_974_9_Left_4568 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_975_9_Left_4569 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_976_9_Left_4570 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_977_9_Left_4571 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_978_9_Left_4572 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_979_9_Left_4573 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_980_9_Left_4574 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_981_9_Left_4575 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_982_9_Left_4576 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_983_9_Left_4577 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_984_9_Left_4578 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_985_9_Left_4579 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_986_9_Left_4580 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_987_9_Left_4581 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_988_9_Left_4582 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_989_9_Left_4583 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_990_9_Left_4584 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_991_9_Left_4585 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_992_9_Left_4586 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_993_9_Left_4587 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_994_9_Left_4588 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_995_9_Left_4589 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_996_9_Left_4590 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_997_9_Left_4591 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_998_9_Left_4592 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_999_9_Left_4593 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1000_9_Left_4594 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1001_9_Left_4595 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1002_9_Left_4596 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1003_9_Left_4597 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1004_9_Left_4598 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1005_9_Left_4599 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1006_9_Left_4600 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1007_9_Left_4601 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1008_9_Left_4602 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1009_9_Left_4603 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1010_9_Left_4604 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1011_9_Left_4605 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1012_9_Left_4606 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1013_9_Left_4607 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1014_9_Left_4608 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1015_9_Left_4609 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1016_9_Left_4610 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1017_9_Left_4611 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1018_9_Left_4612 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1019_9_Left_4613 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1020_9_Left_4614 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1021_9_Left_4615 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1022_9_Left_4616 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1023_9_Left_4617 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1024_9_Left_4618 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1025_9_Left_4619 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1026_9_Left_4620 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1027_9_Left_4621 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1028_9_Left_4622 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1029_9_Left_4623 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1030_9_Left_4624 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1031_9_Left_4625 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1032_9_Left_4626 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1033_9_Left_4627 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1034_9_Left_4628 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1035_9_Left_4629 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1036_9_Left_4630 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1037_9_Left_4631 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1038_9_Left_4632 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1039_9_Left_4633 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1040_9_Left_4634 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1041_9_Left_4635 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1042_9_Left_4636 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1043_9_Left_4637 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1044_9_Left_4638 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1045_9_Left_4639 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1046_9_Left_4640 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1047_9_Left_4641 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1048_9_Left_4642 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1049_9_Left_4643 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1050_9_Left_4644 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1051_9_Left_4645 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1052_9_Left_4646 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1053_9_Left_4647 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1054_9_Left_4648 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1055_9_Left_4649 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1056_9_Left_4650 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1057_9_Left_4651 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_894_1_Right_4652 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_895_1_Right_4653 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_896_1_Right_4654 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_897_1_Right_4655 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_898_1_Right_4656 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_899_1_Right_4657 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_900_1_Right_4658 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_901_1_Right_4659 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_902_1_Right_4660 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_903_1_Right_4661 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_904_1_Right_4662 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_905_1_Right_4663 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_906_1_Right_4664 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_907_1_Right_4665 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_908_1_Right_4666 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_909_1_Right_4667 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_910_1_Right_4668 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_911_1_Right_4669 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_912_1_Right_4670 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_913_1_Right_4671 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_914_1_Right_4672 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_915_1_Right_4673 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_916_1_Right_4674 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_917_1_Right_4675 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_918_1_Right_4676 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_919_1_Right_4677 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_920_1_Right_4678 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_921_1_Right_4679 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_922_1_Right_4680 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_923_1_Right_4681 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_924_1_Right_4682 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_925_1_Right_4683 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_926_1_Right_4684 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_927_1_Right_4685 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_928_1_Right_4686 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_929_1_Right_4687 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_930_1_Right_4688 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_931_1_Right_4689 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_932_1_Right_4690 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_933_1_Right_4691 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_934_1_Right_4692 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_935_1_Right_4693 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_936_1_Right_4694 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_937_1_Right_4695 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_938_1_Right_4696 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_939_1_Right_4697 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_940_1_Right_4698 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_941_1_Right_4699 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_942_1_Right_4700 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_943_1_Right_4701 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_944_1_Right_4702 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_945_1_Right_4703 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_946_1_Right_4704 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_947_1_Right_4705 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_948_1_Right_4706 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_949_1_Right_4707 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_950_1_Right_4708 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_951_1_Right_4709 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_952_1_Right_4710 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_953_1_Right_4711 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_954_1_Right_4712 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_955_1_Right_4713 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_956_1_Right_4714 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_957_1_Right_4715 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_958_1_Right_4716 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_959_1_Right_4717 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_960_1_Right_4718 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_961_1_Right_4719 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_962_1_Right_4720 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_963_1_Right_4721 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_964_1_Right_4722 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_965_1_Right_4723 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_966_1_Right_4724 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_967_1_Right_4725 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_968_1_Right_4726 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_969_1_Right_4727 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_970_1_Right_4728 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_971_1_Right_4729 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_972_1_Right_4730 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_973_1_Right_4731 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_974_1_Right_4732 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_975_1_Right_4733 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_976_1_Right_4734 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_977_1_Right_4735 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_978_1_Right_4736 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_979_1_Right_4737 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_980_1_Right_4738 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_981_1_Right_4739 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_982_1_Right_4740 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_983_1_Right_4741 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_984_1_Right_4742 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_985_1_Right_4743 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_986_1_Right_4744 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_987_1_Right_4745 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_988_1_Right_4746 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_989_1_Right_4747 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_990_1_Right_4748 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_991_1_Right_4749 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_992_1_Right_4750 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_993_1_Right_4751 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_994_1_Right_4752 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_995_1_Right_4753 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_996_1_Right_4754 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_997_1_Right_4755 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_998_1_Right_4756 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_999_1_Right_4757 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1000_1_Right_4758 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1001_1_Right_4759 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1002_1_Right_4760 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1003_1_Right_4761 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1004_1_Right_4762 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1005_1_Right_4763 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1006_1_Right_4764 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1007_1_Right_4765 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1008_1_Right_4766 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1009_1_Right_4767 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1010_1_Right_4768 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1011_1_Right_4769 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1012_1_Right_4770 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1013_1_Right_4771 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1014_1_Right_4772 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1015_1_Right_4773 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1016_1_Right_4774 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1017_1_Right_4775 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1018_1_Right_4776 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1019_1_Right_4777 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1020_1_Right_4778 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1021_1_Right_4779 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1022_1_Right_4780 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1023_1_Right_4781 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1024_1_Right_4782 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1025_1_Right_4783 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1026_1_Right_4784 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1027_1_Right_4785 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1028_1_Right_4786 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1029_1_Right_4787 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1030_1_Right_4788 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1031_1_Right_4789 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1032_1_Right_4790 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1033_1_Right_4791 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1034_1_Right_4792 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1035_1_Right_4793 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1036_1_Right_4794 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1037_1_Right_4795 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1038_1_Right_4796 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1039_1_Right_4797 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1040_1_Right_4798 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1041_1_Right_4799 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1042_1_Right_4800 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1043_1_Right_4801 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1044_1_Right_4802 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1045_1_Right_4803 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1046_1_Right_4804 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1047_1_Right_4805 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1048_1_Right_4806 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1049_1_Right_4807 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1050_1_Right_4808 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1051_1_Right_4809 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1052_1_Right_4810 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1053_1_Right_4811 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1054_1_Right_4812 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1055_1_Right_4813 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1056_1_Right_4814 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1057_1_Right_4815 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1070_9_Left_4816 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1071_9_Left_4817 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1072_9_Left_4818 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1073_9_Left_4819 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1074_9_Left_4820 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1075_9_Left_4821 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1076_9_Left_4822 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1077_9_Left_4823 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1078_9_Left_4824 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1079_9_Left_4825 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1080_9_Left_4826 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1081_9_Left_4827 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1082_9_Left_4828 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1083_9_Left_4829 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1084_9_Left_4830 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1085_9_Left_4831 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1086_9_Left_4832 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1087_9_Left_4833 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1088_9_Left_4834 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1089_9_Left_4835 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1090_9_Left_4836 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1091_9_Left_4837 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1092_9_Left_4838 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1093_9_Left_4839 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1094_9_Left_4840 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1095_9_Left_4841 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1096_9_Left_4842 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1097_9_Left_4843 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1098_9_Left_4844 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1099_9_Left_4845 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1100_9_Left_4846 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1101_9_Left_4847 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1102_9_Left_4848 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1103_9_Left_4849 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1104_9_Left_4850 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1105_9_Left_4851 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1106_9_Left_4852 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1107_9_Left_4853 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1108_9_Left_4854 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1109_9_Left_4855 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1110_9_Left_4856 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1111_9_Left_4857 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1112_9_Left_4858 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1113_9_Left_4859 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1114_9_Left_4860 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1115_9_Left_4861 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1116_9_Left_4862 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1117_9_Left_4863 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1118_9_Left_4864 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1119_9_Left_4865 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1120_9_Left_4866 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1121_9_Left_4867 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1122_9_Left_4868 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1123_9_Left_4869 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1124_9_Left_4870 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1125_9_Left_4871 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1126_9_Left_4872 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1127_9_Left_4873 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1128_9_Left_4874 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1129_9_Left_4875 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1130_9_Left_4876 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1131_9_Left_4877 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1132_9_Left_4878 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1133_9_Left_4879 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1134_9_Left_4880 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1135_9_Left_4881 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1136_9_Left_4882 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1137_9_Left_4883 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1138_9_Left_4884 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1139_9_Left_4885 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1140_9_Left_4886 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1141_9_Left_4887 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1142_9_Left_4888 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1143_9_Left_4889 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1144_9_Left_4890 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1145_9_Left_4891 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1146_9_Left_4892 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1147_9_Left_4893 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1148_9_Left_4894 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1149_9_Left_4895 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1150_9_Left_4896 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1151_9_Left_4897 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1152_9_Left_4898 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1153_9_Left_4899 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1154_9_Left_4900 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1155_9_Left_4901 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1156_9_Left_4902 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1157_9_Left_4903 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1158_9_Left_4904 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1159_9_Left_4905 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1160_9_Left_4906 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1161_9_Left_4907 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1162_9_Left_4908 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1163_9_Left_4909 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1164_9_Left_4910 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1165_9_Left_4911 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1166_9_Left_4912 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1167_9_Left_4913 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1168_9_Left_4914 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1169_9_Left_4915 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1170_9_Left_4916 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1171_9_Left_4917 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1172_9_Left_4918 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1173_9_Left_4919 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1174_9_Left_4920 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1175_9_Left_4921 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1176_9_Left_4922 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1177_9_Left_4923 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1178_9_Left_4924 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1179_9_Left_4925 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1180_9_Left_4926 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1181_9_Left_4927 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1182_9_Left_4928 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1183_9_Left_4929 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1184_9_Left_4930 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1185_9_Left_4931 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1186_9_Left_4932 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1187_9_Left_4933 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1188_9_Left_4934 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1189_9_Left_4935 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1190_9_Left_4936 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1191_9_Left_4937 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1192_9_Left_4938 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1193_9_Left_4939 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1194_9_Left_4940 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1195_9_Left_4941 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1196_9_Left_4942 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1197_9_Left_4943 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1198_9_Left_4944 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1199_9_Left_4945 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1200_9_Left_4946 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1201_9_Left_4947 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1202_9_Left_4948 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1203_9_Left_4949 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1204_9_Left_4950 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1205_9_Left_4951 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1206_9_Left_4952 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1207_9_Left_4953 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1208_9_Left_4954 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1209_9_Left_4955 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1210_9_Left_4956 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1211_9_Left_4957 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1212_9_Left_4958 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1213_9_Left_4959 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1214_9_Left_4960 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1215_9_Left_4961 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1216_9_Left_4962 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1217_9_Left_4963 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1218_9_Left_4964 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1219_9_Left_4965 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1220_9_Left_4966 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1221_9_Left_4967 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1222_9_Left_4968 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1223_9_Left_4969 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1224_9_Left_4970 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1225_9_Left_4971 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1226_9_Left_4972 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1227_9_Left_4973 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1228_9_Left_4974 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1229_9_Left_4975 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1230_9_Left_4976 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1231_9_Left_4977 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1232_9_Left_4978 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1233_9_Left_4979 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1070_1_Right_4980 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1071_1_Right_4981 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1072_1_Right_4982 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1073_1_Right_4983 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1074_1_Right_4984 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1075_1_Right_4985 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1076_1_Right_4986 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1077_1_Right_4987 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1078_1_Right_4988 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1079_1_Right_4989 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1080_1_Right_4990 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1081_1_Right_4991 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1082_1_Right_4992 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1083_1_Right_4993 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1084_1_Right_4994 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1085_1_Right_4995 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1086_1_Right_4996 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1087_1_Right_4997 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1088_1_Right_4998 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1089_1_Right_4999 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1090_1_Right_5000 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1091_1_Right_5001 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1092_1_Right_5002 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1093_1_Right_5003 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1094_1_Right_5004 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1095_1_Right_5005 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1096_1_Right_5006 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1097_1_Right_5007 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1098_1_Right_5008 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1099_1_Right_5009 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1100_1_Right_5010 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1101_1_Right_5011 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1102_1_Right_5012 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1103_1_Right_5013 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1104_1_Right_5014 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1105_1_Right_5015 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1106_1_Right_5016 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1107_1_Right_5017 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1108_1_Right_5018 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1109_1_Right_5019 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1110_1_Right_5020 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1111_1_Right_5021 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1112_1_Right_5022 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1113_1_Right_5023 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1114_1_Right_5024 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1115_1_Right_5025 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1116_1_Right_5026 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1117_1_Right_5027 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1118_1_Right_5028 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1119_1_Right_5029 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1120_1_Right_5030 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1121_1_Right_5031 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1122_1_Right_5032 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1123_1_Right_5033 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1124_1_Right_5034 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1125_1_Right_5035 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1126_1_Right_5036 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1127_1_Right_5037 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1128_1_Right_5038 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1129_1_Right_5039 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1130_1_Right_5040 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1131_1_Right_5041 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1132_1_Right_5042 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1133_1_Right_5043 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1134_1_Right_5044 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1135_1_Right_5045 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1136_1_Right_5046 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1137_1_Right_5047 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1138_1_Right_5048 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1139_1_Right_5049 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1140_1_Right_5050 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1141_1_Right_5051 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1142_1_Right_5052 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1143_1_Right_5053 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1144_1_Right_5054 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1145_1_Right_5055 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1146_1_Right_5056 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1147_1_Right_5057 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1148_1_Right_5058 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1149_1_Right_5059 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1150_1_Right_5060 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1151_1_Right_5061 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1152_1_Right_5062 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1153_1_Right_5063 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1154_1_Right_5064 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1155_1_Right_5065 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1156_1_Right_5066 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1157_1_Right_5067 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1158_1_Right_5068 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1159_1_Right_5069 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1160_1_Right_5070 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1161_1_Right_5071 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1162_1_Right_5072 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1163_1_Right_5073 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1164_1_Right_5074 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1165_1_Right_5075 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1166_1_Right_5076 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1167_1_Right_5077 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1168_1_Right_5078 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1169_1_Right_5079 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1170_1_Right_5080 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1171_1_Right_5081 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1172_1_Right_5082 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1173_1_Right_5083 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1174_1_Right_5084 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1175_1_Right_5085 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1176_1_Right_5086 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1177_1_Right_5087 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1178_1_Right_5088 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1179_1_Right_5089 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1180_1_Right_5090 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1181_1_Right_5091 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1182_1_Right_5092 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1183_1_Right_5093 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1184_1_Right_5094 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1185_1_Right_5095 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1186_1_Right_5096 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1187_1_Right_5097 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1188_1_Right_5098 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1189_1_Right_5099 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1190_1_Right_5100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1191_1_Right_5101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1192_1_Right_5102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1193_1_Right_5103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1194_1_Right_5104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1195_1_Right_5105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1196_1_Right_5106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1197_1_Right_5107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1198_1_Right_5108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1199_1_Right_5109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1200_1_Right_5110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1201_1_Right_5111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1202_1_Right_5112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1203_1_Right_5113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1204_1_Right_5114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1205_1_Right_5115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1206_1_Right_5116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1207_1_Right_5117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1208_1_Right_5118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1209_1_Right_5119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1210_1_Right_5120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1211_1_Right_5121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1212_1_Right_5122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1213_1_Right_5123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1214_1_Right_5124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1215_1_Right_5125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1216_1_Right_5126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1217_1_Right_5127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1218_1_Right_5128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1219_1_Right_5129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1220_1_Right_5130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1221_1_Right_5131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1222_1_Right_5132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1223_1_Right_5133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1224_1_Right_5134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1225_1_Right_5135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1226_1_Right_5136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1227_1_Right_5137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1228_1_Right_5138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1229_1_Right_5139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1230_1_Right_5140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1231_1_Right_5141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1232_1_Right_5142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1233_1_Right_5143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1246_9_Left_5144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1247_9_Left_5145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1248_9_Left_5146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1249_9_Left_5147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1250_9_Left_5148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1251_9_Left_5149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1252_9_Left_5150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1253_9_Left_5151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1254_9_Left_5152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1255_9_Left_5153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1256_9_Left_5154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1257_9_Left_5155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1258_9_Left_5156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1259_9_Left_5157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1260_9_Left_5158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1261_9_Left_5159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1262_9_Left_5160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1263_9_Left_5161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1264_9_Left_5162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1265_9_Left_5163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1266_9_Left_5164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1267_9_Left_5165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1268_9_Left_5166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1269_9_Left_5167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1270_9_Left_5168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1271_9_Left_5169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1272_9_Left_5170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1273_9_Left_5171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1274_9_Left_5172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1275_9_Left_5173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1276_9_Left_5174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1277_9_Left_5175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1278_9_Left_5176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1279_9_Left_5177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1280_9_Left_5178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1281_9_Left_5179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1282_9_Left_5180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1283_9_Left_5181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1284_9_Left_5182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1285_9_Left_5183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1286_9_Left_5184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1287_9_Left_5185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1288_9_Left_5186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1289_9_Left_5187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1290_9_Left_5188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1291_9_Left_5189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1292_9_Left_5190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1293_9_Left_5191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1294_9_Left_5192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1295_9_Left_5193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1296_9_Left_5194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1297_9_Left_5195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1298_9_Left_5196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1299_9_Left_5197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1300_9_Left_5198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1301_9_Left_5199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1302_9_Left_5200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1303_9_Left_5201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1304_9_Left_5202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1305_9_Left_5203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1306_9_Left_5204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1307_9_Left_5205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1308_9_Left_5206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1309_9_Left_5207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1310_9_Left_5208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1311_9_Left_5209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1312_9_Left_5210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1313_9_Left_5211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1314_9_Left_5212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1315_9_Left_5213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1316_9_Left_5214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1317_9_Left_5215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1318_9_Left_5216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1319_9_Left_5217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1320_9_Left_5218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1321_9_Left_5219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1322_9_Left_5220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1323_9_Left_5221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1324_9_Left_5222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1325_9_Left_5223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1326_9_Left_5224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1327_9_Left_5225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1328_9_Left_5226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1329_9_Left_5227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1330_9_Left_5228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1331_9_Left_5229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1332_9_Left_5230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1333_9_Left_5231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1334_9_Left_5232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1335_9_Left_5233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1336_9_Left_5234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1337_9_Left_5235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1338_9_Left_5236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1339_9_Left_5237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1340_9_Left_5238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1341_9_Left_5239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1342_9_Left_5240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1343_9_Left_5241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1344_9_Left_5242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1345_9_Left_5243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1346_9_Left_5244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1347_9_Left_5245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1348_9_Left_5246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1349_9_Left_5247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1350_9_Left_5248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1351_9_Left_5249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1352_9_Left_5250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1353_9_Left_5251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1354_9_Left_5252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1355_9_Left_5253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1356_9_Left_5254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1357_9_Left_5255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1358_9_Left_5256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1359_9_Left_5257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1360_9_Left_5258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1361_9_Left_5259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1362_9_Left_5260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1363_9_Left_5261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1364_9_Left_5262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1365_9_Left_5263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1366_9_Left_5264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1367_9_Left_5265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1368_9_Left_5266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1369_9_Left_5267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1370_9_Left_5268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1371_9_Left_5269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1372_9_Left_5270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1373_9_Left_5271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1374_9_Left_5272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1375_9_Left_5273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1376_9_Left_5274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1377_9_Left_5275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1378_9_Left_5276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1379_9_Left_5277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1380_9_Left_5278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1381_9_Left_5279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1382_9_Left_5280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1383_9_Left_5281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1384_9_Left_5282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1385_9_Left_5283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1386_9_Left_5284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1387_9_Left_5285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1388_9_Left_5286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1389_9_Left_5287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1390_9_Left_5288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1391_9_Left_5289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1392_9_Left_5290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1393_9_Left_5291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1394_9_Left_5292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1395_9_Left_5293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1396_9_Left_5294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1397_9_Left_5295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1398_9_Left_5296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1399_9_Left_5297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1400_9_Left_5298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1401_9_Left_5299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1402_9_Left_5300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1403_9_Left_5301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1404_9_Left_5302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1405_9_Left_5303 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1406_9_Left_5304 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1407_9_Left_5305 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1408_9_Left_5306 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1409_9_Left_5307 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1246_1_Right_5308 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1247_1_Right_5309 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1248_1_Right_5310 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1249_1_Right_5311 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1250_1_Right_5312 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1251_1_Right_5313 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1252_1_Right_5314 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1253_1_Right_5315 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1254_1_Right_5316 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1255_1_Right_5317 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1256_1_Right_5318 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1257_1_Right_5319 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1258_1_Right_5320 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1259_1_Right_5321 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1260_1_Right_5322 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1261_1_Right_5323 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1262_1_Right_5324 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1263_1_Right_5325 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1264_1_Right_5326 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1265_1_Right_5327 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1266_1_Right_5328 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1267_1_Right_5329 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1268_1_Right_5330 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1269_1_Right_5331 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1270_1_Right_5332 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1271_1_Right_5333 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1272_1_Right_5334 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1273_1_Right_5335 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1274_1_Right_5336 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1275_1_Right_5337 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1276_1_Right_5338 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1277_1_Right_5339 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1278_1_Right_5340 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1279_1_Right_5341 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1280_1_Right_5342 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1281_1_Right_5343 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1282_1_Right_5344 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1283_1_Right_5345 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1284_1_Right_5346 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1285_1_Right_5347 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1286_1_Right_5348 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1287_1_Right_5349 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1288_1_Right_5350 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1289_1_Right_5351 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1290_1_Right_5352 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1291_1_Right_5353 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1292_1_Right_5354 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1293_1_Right_5355 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1294_1_Right_5356 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1295_1_Right_5357 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1296_1_Right_5358 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1297_1_Right_5359 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1298_1_Right_5360 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1299_1_Right_5361 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1300_1_Right_5362 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1301_1_Right_5363 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1302_1_Right_5364 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1303_1_Right_5365 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1304_1_Right_5366 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1305_1_Right_5367 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1306_1_Right_5368 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1307_1_Right_5369 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1308_1_Right_5370 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1309_1_Right_5371 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1310_1_Right_5372 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1311_1_Right_5373 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1312_1_Right_5374 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1313_1_Right_5375 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1314_1_Right_5376 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1315_1_Right_5377 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1316_1_Right_5378 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1317_1_Right_5379 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1318_1_Right_5380 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1319_1_Right_5381 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1320_1_Right_5382 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1321_1_Right_5383 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1322_1_Right_5384 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1323_1_Right_5385 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1324_1_Right_5386 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1325_1_Right_5387 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1326_1_Right_5388 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1327_1_Right_5389 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1328_1_Right_5390 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1329_1_Right_5391 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1330_1_Right_5392 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1331_1_Right_5393 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1332_1_Right_5394 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1333_1_Right_5395 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1334_1_Right_5396 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1335_1_Right_5397 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1336_1_Right_5398 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1337_1_Right_5399 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1338_1_Right_5400 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1339_1_Right_5401 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1340_1_Right_5402 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1341_1_Right_5403 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1342_1_Right_5404 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1343_1_Right_5405 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1344_1_Right_5406 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1345_1_Right_5407 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1346_1_Right_5408 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1347_1_Right_5409 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1348_1_Right_5410 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1349_1_Right_5411 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1350_1_Right_5412 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1351_1_Right_5413 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1352_1_Right_5414 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1353_1_Right_5415 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1354_1_Right_5416 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1355_1_Right_5417 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1356_1_Right_5418 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1357_1_Right_5419 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1358_1_Right_5420 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1359_1_Right_5421 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1360_1_Right_5422 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1361_1_Right_5423 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1362_1_Right_5424 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1363_1_Right_5425 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1364_1_Right_5426 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1365_1_Right_5427 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1366_1_Right_5428 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1367_1_Right_5429 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1368_1_Right_5430 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1369_1_Right_5431 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1370_1_Right_5432 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1371_1_Right_5433 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1372_1_Right_5434 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1373_1_Right_5435 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1374_1_Right_5436 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1375_1_Right_5437 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1376_1_Right_5438 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1377_1_Right_5439 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1378_1_Right_5440 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1379_1_Right_5441 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1380_1_Right_5442 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1381_1_Right_5443 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1382_1_Right_5444 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1383_1_Right_5445 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1384_1_Right_5446 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1385_1_Right_5447 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1386_1_Right_5448 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1387_1_Right_5449 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1388_1_Right_5450 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1389_1_Right_5451 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1390_1_Right_5452 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1391_1_Right_5453 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1392_1_Right_5454 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1393_1_Right_5455 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1394_1_Right_5456 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1395_1_Right_5457 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1396_1_Right_5458 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1397_1_Right_5459 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1398_1_Right_5460 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1399_1_Right_5461 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1400_1_Right_5462 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1401_1_Right_5463 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1402_1_Right_5464 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1403_1_Right_5465 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1404_1_Right_5466 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1405_1_Right_5467 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1406_1_Right_5468 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1407_1_Right_5469 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1408_1_Right_5470 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1409_1_Right_5471 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5472 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5473 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5474 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5475 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5476 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5477 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5478 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5479 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5480 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5481 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5482 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5483 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5484 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_5485 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_5486 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_5487 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_5488 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_5489 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_5490 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_5491 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1_5492 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_5493 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_5494 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_5495 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_5496 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_5497 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_5498 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_5499 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_5500 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_5501 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_5502 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_5503 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_5504 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_5505 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_3_5506 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_5507 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_5508 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_5509 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_5510 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_5511 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_5512 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_5513 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_5514 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_5515 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_5516 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_5517 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_5518 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_5519 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_5_5520 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_5521 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_5522 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_5523 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_5524 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_5525 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_5526 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_5527 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_5528 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_5529 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_5530 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_5531 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_5532 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_5533 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_7_5534 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_5535 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_5536 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_5537 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_5538 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_5539 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_5540 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_5541 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_5542 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_5543 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_5544 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_5545 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_5546 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_5547 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_9_5548 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_5549 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_5550 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_5551 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_5552 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_5553 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_5554 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_5555 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_5556 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_5557 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_5558 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_5559 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_5560 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_5561 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_11_5562 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_5563 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_5564 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_5565 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_5566 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_5567 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_5568 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_5569 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5570 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5571 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5572 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5573 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5574 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5575 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5576 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5577 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5578 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5579 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5580 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5581 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5582 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_13_5583 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5584 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5585 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5586 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5587 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5588 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5589 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5590 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5591 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5592 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5593 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5594 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5595 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5596 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_178_5597 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_5598 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_5599 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_5600 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_5601 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_5602 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_5603 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_179_5604 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_5605 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_5606 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_5607 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_5608 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_5609 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_5610 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_180_5611 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_5612 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_5613 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_5614 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_5615 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_5616 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_5617 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_181_5618 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_5619 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_5620 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_5621 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_5622 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_5623 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_5624 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_182_5625 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_5626 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_5627 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_5628 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_5629 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_5630 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_5631 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_183_5632 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_5633 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_5634 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_5635 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_5636 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_5637 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_5638 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_184_5639 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_5640 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_5641 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_5642 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_5643 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_5644 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_5645 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_185_5646 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_5647 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_5648 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_5649 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_5650 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_5651 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_5652 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_186_5653 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_5654 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_5655 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_5656 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_5657 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_5658 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_5659 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_187_5660 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_5661 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_5662 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_5663 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_5664 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_5665 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_5666 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_188_5667 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5668 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5669 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5670 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5671 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5672 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5673 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5674 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5675 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5676 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5677 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5678 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5679 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5680 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_189_5681 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5682 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5683 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5684 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5685 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5686 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5687 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5688 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5689 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5690 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5691 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5692 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5693 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5694 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_354_5695 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_355_5696 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_355_5697 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_355_5698 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_355_5699 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_355_5700 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_355_5701 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_355_5702 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_356_5703 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_356_5704 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_356_5705 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_356_5706 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_356_5707 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_356_5708 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_356_5709 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_357_5710 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_357_5711 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_357_5712 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_357_5713 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_357_5714 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_357_5715 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_357_5716 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_358_5717 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_358_5718 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_358_5719 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_358_5720 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_358_5721 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_358_5722 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_358_5723 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_359_5724 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_359_5725 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_359_5726 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_359_5727 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_359_5728 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_359_5729 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_359_5730 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_360_5731 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_360_5732 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_360_5733 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_360_5734 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_360_5735 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_360_5736 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_360_5737 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_361_5738 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_361_5739 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_361_5740 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_361_5741 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_361_5742 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_361_5743 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_361_5744 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_362_5745 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_362_5746 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_362_5747 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_362_5748 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_362_5749 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_362_5750 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_362_5751 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_363_5752 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_363_5753 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_363_5754 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_363_5755 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_363_5756 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_363_5757 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_363_5758 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_364_5759 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_364_5760 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_364_5761 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_364_5762 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_364_5763 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_364_5764 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_364_5765 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5766 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5767 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5768 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5769 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5770 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5771 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5772 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5773 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5774 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5775 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5776 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5777 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5778 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_365_5779 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5780 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5781 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5782 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5783 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5784 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5785 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5786 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5787 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5788 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5789 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5790 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5791 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5792 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_530_5793 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_531_5794 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_531_5795 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_531_5796 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_531_5797 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_531_5798 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_531_5799 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_531_5800 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_532_5801 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_532_5802 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_532_5803 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_532_5804 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_532_5805 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_532_5806 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_532_5807 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_533_5808 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_533_5809 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_533_5810 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_533_5811 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_533_5812 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_533_5813 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_533_5814 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_534_5815 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_534_5816 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_534_5817 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_534_5818 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_534_5819 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_534_5820 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_534_5821 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_535_5822 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_535_5823 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_535_5824 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_535_5825 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_535_5826 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_535_5827 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_535_5828 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_536_5829 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_536_5830 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_536_5831 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_536_5832 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_536_5833 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_536_5834 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_536_5835 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_537_5836 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_537_5837 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_537_5838 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_537_5839 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_537_5840 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_537_5841 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_537_5842 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_538_5843 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_538_5844 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_538_5845 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_538_5846 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_538_5847 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_538_5848 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_538_5849 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_539_5850 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_539_5851 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_539_5852 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_539_5853 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_539_5854 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_539_5855 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_539_5856 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_540_5857 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_540_5858 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_540_5859 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_540_5860 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_540_5861 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_540_5862 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_540_5863 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5864 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5865 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5866 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5867 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5868 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5869 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5870 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5871 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5872 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5873 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5874 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5875 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5876 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_541_5877 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5878 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5879 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5880 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5881 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5882 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5883 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5884 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5885 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5886 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5887 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5888 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5889 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5890 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_706_5891 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_707_5892 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_707_5893 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_707_5894 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_707_5895 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_707_5896 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_707_5897 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_707_5898 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_708_5899 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_708_5900 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_708_5901 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_708_5902 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_708_5903 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_708_5904 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_708_5905 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_709_5906 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_709_5907 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_709_5908 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_709_5909 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_709_5910 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_709_5911 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_709_5912 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_710_5913 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_710_5914 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_710_5915 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_710_5916 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_710_5917 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_710_5918 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_710_5919 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_711_5920 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_711_5921 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_711_5922 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_711_5923 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_711_5924 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_711_5925 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_711_5926 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_712_5927 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_712_5928 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_712_5929 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_712_5930 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_712_5931 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_712_5932 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_712_5933 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_713_5934 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_713_5935 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_713_5936 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_713_5937 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_713_5938 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_713_5939 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_713_5940 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_714_5941 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_714_5942 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_714_5943 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_714_5944 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_714_5945 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_714_5946 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_714_5947 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_715_5948 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_715_5949 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_715_5950 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_715_5951 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_715_5952 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_715_5953 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_715_5954 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_716_5955 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_716_5956 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_716_5957 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_716_5958 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_716_5959 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_716_5960 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_716_5961 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5962 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5963 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5964 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5965 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5966 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5967 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5968 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5969 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5970 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5971 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5972 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5973 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5974 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_717_5975 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5976 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5977 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5978 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5979 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5980 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5981 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5982 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5983 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5984 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5985 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5986 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5987 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5988 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_882_5989 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_883_5990 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_883_5991 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_883_5992 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_883_5993 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_883_5994 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_883_5995 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_883_5996 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_884_5997 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_884_5998 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_884_5999 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_884_6000 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_884_6001 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_884_6002 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_884_6003 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_885_6004 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_885_6005 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_885_6006 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_885_6007 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_885_6008 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_885_6009 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_885_6010 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_886_6011 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_886_6012 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_886_6013 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_886_6014 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_886_6015 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_886_6016 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_886_6017 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_887_6018 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_887_6019 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_887_6020 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_887_6021 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_887_6022 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_887_6023 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_887_6024 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_888_6025 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_888_6026 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_888_6027 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_888_6028 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_888_6029 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_888_6030 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_888_6031 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_889_6032 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_889_6033 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_889_6034 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_889_6035 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_889_6036 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_889_6037 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_889_6038 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_890_6039 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_890_6040 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_890_6041 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_890_6042 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_890_6043 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_890_6044 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_890_6045 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_891_6046 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_891_6047 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_891_6048 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_891_6049 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_891_6050 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_891_6051 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_891_6052 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_892_6053 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_892_6054 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_892_6055 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_892_6056 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_892_6057 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_892_6058 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_892_6059 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6060 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6061 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6062 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6063 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6064 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6065 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6066 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6067 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6068 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6069 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6070 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6071 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6072 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_893_6073 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6074 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6075 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6076 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6077 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6078 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6079 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6080 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6081 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6082 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6083 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6084 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6085 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6086 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1058_6087 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1059_6088 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1059_6089 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1059_6090 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1059_6091 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1059_6092 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1059_6093 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1059_6094 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1060_6095 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1060_6096 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1060_6097 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1060_6098 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1060_6099 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1060_6100 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1060_6101 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1061_6102 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1061_6103 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1061_6104 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1061_6105 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1061_6106 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1061_6107 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1061_6108 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1062_6109 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1062_6110 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1062_6111 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1062_6112 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1062_6113 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1062_6114 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1062_6115 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1063_6116 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1063_6117 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1063_6118 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1063_6119 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1063_6120 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1063_6121 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1063_6122 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1064_6123 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1064_6124 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1064_6125 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1064_6126 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1064_6127 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1064_6128 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1064_6129 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1065_6130 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1065_6131 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1065_6132 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1065_6133 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1065_6134 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1065_6135 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1065_6136 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1066_6137 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1066_6138 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1066_6139 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1066_6140 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1066_6141 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1066_6142 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1066_6143 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1067_6144 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1067_6145 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1067_6146 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1067_6147 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1067_6148 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1067_6149 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1067_6150 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1068_6151 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1068_6152 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1068_6153 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1068_6154 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1068_6155 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1068_6156 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1068_6157 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6158 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6159 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6160 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6161 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6162 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6163 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6164 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6165 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6166 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6167 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6168 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6169 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6170 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1069_6171 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6172 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6173 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6174 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6175 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6176 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6177 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6178 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6179 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6180 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6181 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6182 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6183 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6184 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1234_6185 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1235_6186 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1235_6187 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1235_6188 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1235_6189 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1235_6190 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1235_6191 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1235_6192 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1236_6193 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1236_6194 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1236_6195 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1236_6196 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1236_6197 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1236_6198 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1236_6199 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1237_6200 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1237_6201 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1237_6202 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1237_6203 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1237_6204 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1237_6205 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1237_6206 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1238_6207 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1238_6208 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1238_6209 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1238_6210 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1238_6211 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1238_6212 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1238_6213 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1239_6214 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1239_6215 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1239_6216 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1239_6217 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1239_6218 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1239_6219 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1239_6220 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1240_6221 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1240_6222 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1240_6223 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1240_6224 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1240_6225 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1240_6226 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1240_6227 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1241_6228 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1241_6229 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1241_6230 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1241_6231 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1241_6232 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1241_6233 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1241_6234 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1242_6235 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1242_6236 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1242_6237 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1242_6238 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1242_6239 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1242_6240 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1242_6241 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1243_6242 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1243_6243 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1243_6244 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1243_6245 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1243_6246 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1243_6247 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1243_6248 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1244_6249 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1244_6250 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1244_6251 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1244_6252 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1244_6253 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1244_6254 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1244_6255 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6256 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6257 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6258 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6259 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6260 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6261 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6262 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6263 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6264 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6265 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6266 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6267 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6268 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1245_6269 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6270 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6271 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6272 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6273 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6274 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6275 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6276 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6277 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6278 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6279 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6280 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6281 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6282 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1410_6283 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1411_6284 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1411_6285 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1411_6286 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1411_6287 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1411_6288 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1411_6289 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1411_6290 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1412_6291 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1412_6292 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1412_6293 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1412_6294 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1412_6295 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1412_6296 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1412_6297 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1413_6298 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1413_6299 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1413_6300 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1413_6301 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1413_6302 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1413_6303 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1413_6304 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1414_6305 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1414_6306 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1414_6307 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1414_6308 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1414_6309 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1414_6310 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1414_6311 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1415_6312 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1415_6313 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1415_6314 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1415_6315 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1415_6316 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1415_6317 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1415_6318 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1416_6319 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1416_6320 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1416_6321 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1416_6322 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1416_6323 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1416_6324 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1416_6325 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1417_6326 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1417_6327 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1417_6328 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1417_6329 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1417_6330 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1417_6331 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1417_6332 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1418_6333 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1418_6334 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1418_6335 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1418_6336 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1418_6337 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1418_6338 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1418_6339 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1419_6340 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1419_6341 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1419_6342 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1419_6343 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1419_6344 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1419_6345 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1419_6346 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1420_6347 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1420_6348 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1420_6349 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1420_6350 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1420_6351 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1420_6352 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1420_6353 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1421_6354 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1421_6355 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1421_6356 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1421_6357 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1421_6358 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1421_6359 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1421_6360 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1422_6361 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1422_6362 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1422_6363 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1422_6364 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1422_6365 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1422_6366 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1422_6367 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6368 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6369 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6370 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6371 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6372 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6373 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6374 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6375 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6376 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6377 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6378 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6379 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6380 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_1423_6381 ();
 BUFx2_ASAP7_75t_R input1 (.A(io_ins_down_0[0]),
    .Y(net1));
 BUFx2_ASAP7_75t_R input2 (.A(io_ins_down_0[10]),
    .Y(net2));
 BUFx2_ASAP7_75t_R input3 (.A(io_ins_down_0[11]),
    .Y(net3));
 BUFx2_ASAP7_75t_R input4 (.A(io_ins_down_0[12]),
    .Y(net4));
 BUFx2_ASAP7_75t_R input5 (.A(io_ins_down_0[13]),
    .Y(net5));
 BUFx2_ASAP7_75t_R input6 (.A(io_ins_down_0[14]),
    .Y(net6));
 BUFx2_ASAP7_75t_R input7 (.A(io_ins_down_0[15]),
    .Y(net7));
 BUFx2_ASAP7_75t_R input8 (.A(io_ins_down_0[16]),
    .Y(net8));
 BUFx2_ASAP7_75t_R input9 (.A(io_ins_down_0[17]),
    .Y(net9));
 BUFx2_ASAP7_75t_R input10 (.A(io_ins_down_0[18]),
    .Y(net10));
 BUFx2_ASAP7_75t_R input11 (.A(io_ins_down_0[19]),
    .Y(net11));
 BUFx2_ASAP7_75t_R input12 (.A(io_ins_down_0[1]),
    .Y(net12));
 BUFx2_ASAP7_75t_R input13 (.A(io_ins_down_0[20]),
    .Y(net13));
 BUFx2_ASAP7_75t_R input14 (.A(io_ins_down_0[21]),
    .Y(net14));
 BUFx2_ASAP7_75t_R input15 (.A(io_ins_down_0[22]),
    .Y(net15));
 BUFx2_ASAP7_75t_R input16 (.A(io_ins_down_0[23]),
    .Y(net16));
 BUFx2_ASAP7_75t_R input17 (.A(io_ins_down_0[24]),
    .Y(net17));
 BUFx2_ASAP7_75t_R input18 (.A(io_ins_down_0[25]),
    .Y(net18));
 BUFx2_ASAP7_75t_R input19 (.A(io_ins_down_0[26]),
    .Y(net19));
 BUFx2_ASAP7_75t_R input20 (.A(io_ins_down_0[27]),
    .Y(net20));
 BUFx2_ASAP7_75t_R input21 (.A(io_ins_down_0[28]),
    .Y(net21));
 BUFx2_ASAP7_75t_R input22 (.A(io_ins_down_0[29]),
    .Y(net22));
 BUFx2_ASAP7_75t_R input23 (.A(io_ins_down_0[2]),
    .Y(net23));
 BUFx2_ASAP7_75t_R input24 (.A(io_ins_down_0[30]),
    .Y(net24));
 BUFx2_ASAP7_75t_R input25 (.A(io_ins_down_0[31]),
    .Y(net25));
 BUFx2_ASAP7_75t_R input26 (.A(io_ins_down_0[32]),
    .Y(net26));
 BUFx2_ASAP7_75t_R input27 (.A(io_ins_down_0[33]),
    .Y(net27));
 BUFx2_ASAP7_75t_R input28 (.A(io_ins_down_0[34]),
    .Y(net28));
 BUFx2_ASAP7_75t_R input29 (.A(io_ins_down_0[35]),
    .Y(net29));
 BUFx2_ASAP7_75t_R input30 (.A(io_ins_down_0[36]),
    .Y(net30));
 BUFx2_ASAP7_75t_R input31 (.A(io_ins_down_0[37]),
    .Y(net31));
 BUFx2_ASAP7_75t_R input32 (.A(io_ins_down_0[38]),
    .Y(net32));
 BUFx2_ASAP7_75t_R input33 (.A(io_ins_down_0[39]),
    .Y(net33));
 BUFx2_ASAP7_75t_R input34 (.A(io_ins_down_0[3]),
    .Y(net34));
 BUFx2_ASAP7_75t_R input35 (.A(io_ins_down_0[40]),
    .Y(net35));
 BUFx2_ASAP7_75t_R input36 (.A(io_ins_down_0[41]),
    .Y(net36));
 BUFx2_ASAP7_75t_R input37 (.A(io_ins_down_0[42]),
    .Y(net37));
 BUFx2_ASAP7_75t_R input38 (.A(io_ins_down_0[43]),
    .Y(net38));
 BUFx2_ASAP7_75t_R input39 (.A(io_ins_down_0[44]),
    .Y(net39));
 BUFx2_ASAP7_75t_R input40 (.A(io_ins_down_0[45]),
    .Y(net40));
 BUFx2_ASAP7_75t_R input41 (.A(io_ins_down_0[46]),
    .Y(net41));
 BUFx2_ASAP7_75t_R input42 (.A(io_ins_down_0[47]),
    .Y(net42));
 BUFx2_ASAP7_75t_R input43 (.A(io_ins_down_0[48]),
    .Y(net43));
 BUFx2_ASAP7_75t_R input44 (.A(io_ins_down_0[49]),
    .Y(net44));
 BUFx2_ASAP7_75t_R input45 (.A(io_ins_down_0[4]),
    .Y(net45));
 BUFx2_ASAP7_75t_R input46 (.A(io_ins_down_0[50]),
    .Y(net46));
 BUFx2_ASAP7_75t_R input47 (.A(io_ins_down_0[51]),
    .Y(net47));
 BUFx2_ASAP7_75t_R input48 (.A(io_ins_down_0[52]),
    .Y(net48));
 BUFx2_ASAP7_75t_R input49 (.A(io_ins_down_0[53]),
    .Y(net49));
 BUFx2_ASAP7_75t_R input50 (.A(io_ins_down_0[54]),
    .Y(net50));
 BUFx2_ASAP7_75t_R input51 (.A(io_ins_down_0[55]),
    .Y(net51));
 BUFx2_ASAP7_75t_R input52 (.A(io_ins_down_0[56]),
    .Y(net52));
 BUFx2_ASAP7_75t_R input53 (.A(io_ins_down_0[57]),
    .Y(net53));
 BUFx2_ASAP7_75t_R input54 (.A(io_ins_down_0[58]),
    .Y(net54));
 BUFx2_ASAP7_75t_R input55 (.A(io_ins_down_0[59]),
    .Y(net55));
 BUFx2_ASAP7_75t_R input56 (.A(io_ins_down_0[5]),
    .Y(net56));
 BUFx2_ASAP7_75t_R input57 (.A(io_ins_down_0[60]),
    .Y(net57));
 BUFx2_ASAP7_75t_R input58 (.A(io_ins_down_0[61]),
    .Y(net58));
 BUFx2_ASAP7_75t_R input59 (.A(io_ins_down_0[62]),
    .Y(net59));
 BUFx2_ASAP7_75t_R input60 (.A(io_ins_down_0[63]),
    .Y(net60));
 BUFx2_ASAP7_75t_R input61 (.A(io_ins_down_0[6]),
    .Y(net61));
 BUFx2_ASAP7_75t_R input62 (.A(io_ins_down_0[7]),
    .Y(net62));
 BUFx2_ASAP7_75t_R input63 (.A(io_ins_down_0[8]),
    .Y(net63));
 BUFx2_ASAP7_75t_R input64 (.A(io_ins_down_0[9]),
    .Y(net64));
 BUFx2_ASAP7_75t_R input65 (.A(io_ins_down_1[0]),
    .Y(net65));
 BUFx2_ASAP7_75t_R input66 (.A(io_ins_down_1[10]),
    .Y(net66));
 BUFx2_ASAP7_75t_R input67 (.A(io_ins_down_1[11]),
    .Y(net67));
 BUFx2_ASAP7_75t_R input68 (.A(io_ins_down_1[12]),
    .Y(net68));
 BUFx2_ASAP7_75t_R input69 (.A(io_ins_down_1[13]),
    .Y(net69));
 BUFx2_ASAP7_75t_R input70 (.A(io_ins_down_1[14]),
    .Y(net70));
 BUFx2_ASAP7_75t_R input71 (.A(io_ins_down_1[15]),
    .Y(net71));
 BUFx2_ASAP7_75t_R input72 (.A(io_ins_down_1[16]),
    .Y(net72));
 BUFx2_ASAP7_75t_R input73 (.A(io_ins_down_1[17]),
    .Y(net73));
 BUFx2_ASAP7_75t_R input74 (.A(io_ins_down_1[18]),
    .Y(net74));
 BUFx2_ASAP7_75t_R input75 (.A(io_ins_down_1[19]),
    .Y(net75));
 BUFx2_ASAP7_75t_R input76 (.A(io_ins_down_1[1]),
    .Y(net76));
 BUFx2_ASAP7_75t_R input77 (.A(io_ins_down_1[20]),
    .Y(net77));
 BUFx2_ASAP7_75t_R input78 (.A(io_ins_down_1[21]),
    .Y(net78));
 BUFx2_ASAP7_75t_R input79 (.A(io_ins_down_1[22]),
    .Y(net79));
 BUFx2_ASAP7_75t_R input80 (.A(io_ins_down_1[23]),
    .Y(net80));
 BUFx2_ASAP7_75t_R input81 (.A(io_ins_down_1[24]),
    .Y(net81));
 BUFx2_ASAP7_75t_R input82 (.A(io_ins_down_1[25]),
    .Y(net82));
 BUFx2_ASAP7_75t_R input83 (.A(io_ins_down_1[26]),
    .Y(net83));
 BUFx2_ASAP7_75t_R input84 (.A(io_ins_down_1[27]),
    .Y(net84));
 BUFx2_ASAP7_75t_R input85 (.A(io_ins_down_1[28]),
    .Y(net85));
 BUFx2_ASAP7_75t_R input86 (.A(io_ins_down_1[29]),
    .Y(net86));
 BUFx2_ASAP7_75t_R input87 (.A(io_ins_down_1[2]),
    .Y(net87));
 BUFx2_ASAP7_75t_R input88 (.A(io_ins_down_1[30]),
    .Y(net88));
 BUFx2_ASAP7_75t_R input89 (.A(io_ins_down_1[31]),
    .Y(net89));
 BUFx2_ASAP7_75t_R input90 (.A(io_ins_down_1[32]),
    .Y(net90));
 BUFx2_ASAP7_75t_R input91 (.A(io_ins_down_1[33]),
    .Y(net91));
 BUFx2_ASAP7_75t_R input92 (.A(io_ins_down_1[34]),
    .Y(net92));
 BUFx2_ASAP7_75t_R input93 (.A(io_ins_down_1[35]),
    .Y(net93));
 BUFx2_ASAP7_75t_R input94 (.A(io_ins_down_1[36]),
    .Y(net94));
 BUFx2_ASAP7_75t_R input95 (.A(io_ins_down_1[37]),
    .Y(net95));
 BUFx2_ASAP7_75t_R input96 (.A(io_ins_down_1[38]),
    .Y(net96));
 BUFx2_ASAP7_75t_R input97 (.A(io_ins_down_1[39]),
    .Y(net97));
 BUFx2_ASAP7_75t_R input98 (.A(io_ins_down_1[3]),
    .Y(net98));
 BUFx2_ASAP7_75t_R input99 (.A(io_ins_down_1[40]),
    .Y(net99));
 BUFx2_ASAP7_75t_R input100 (.A(io_ins_down_1[41]),
    .Y(net100));
 BUFx2_ASAP7_75t_R input101 (.A(io_ins_down_1[42]),
    .Y(net101));
 BUFx2_ASAP7_75t_R input102 (.A(io_ins_down_1[43]),
    .Y(net102));
 BUFx2_ASAP7_75t_R input103 (.A(io_ins_down_1[44]),
    .Y(net103));
 BUFx2_ASAP7_75t_R input104 (.A(io_ins_down_1[45]),
    .Y(net104));
 BUFx2_ASAP7_75t_R input105 (.A(io_ins_down_1[46]),
    .Y(net105));
 BUFx2_ASAP7_75t_R input106 (.A(io_ins_down_1[47]),
    .Y(net106));
 BUFx2_ASAP7_75t_R input107 (.A(io_ins_down_1[48]),
    .Y(net107));
 BUFx2_ASAP7_75t_R input108 (.A(io_ins_down_1[49]),
    .Y(net108));
 BUFx2_ASAP7_75t_R input109 (.A(io_ins_down_1[4]),
    .Y(net109));
 BUFx2_ASAP7_75t_R input110 (.A(io_ins_down_1[50]),
    .Y(net110));
 BUFx2_ASAP7_75t_R input111 (.A(io_ins_down_1[51]),
    .Y(net111));
 BUFx2_ASAP7_75t_R input112 (.A(io_ins_down_1[52]),
    .Y(net112));
 BUFx2_ASAP7_75t_R input113 (.A(io_ins_down_1[53]),
    .Y(net113));
 BUFx2_ASAP7_75t_R input114 (.A(io_ins_down_1[54]),
    .Y(net114));
 BUFx2_ASAP7_75t_R input115 (.A(io_ins_down_1[55]),
    .Y(net115));
 BUFx2_ASAP7_75t_R input116 (.A(io_ins_down_1[56]),
    .Y(net116));
 BUFx2_ASAP7_75t_R input117 (.A(io_ins_down_1[57]),
    .Y(net117));
 BUFx2_ASAP7_75t_R input118 (.A(io_ins_down_1[58]),
    .Y(net118));
 BUFx2_ASAP7_75t_R input119 (.A(io_ins_down_1[59]),
    .Y(net119));
 BUFx2_ASAP7_75t_R input120 (.A(io_ins_down_1[5]),
    .Y(net120));
 BUFx2_ASAP7_75t_R input121 (.A(io_ins_down_1[60]),
    .Y(net121));
 BUFx2_ASAP7_75t_R input122 (.A(io_ins_down_1[61]),
    .Y(net122));
 BUFx2_ASAP7_75t_R input123 (.A(io_ins_down_1[62]),
    .Y(net123));
 BUFx2_ASAP7_75t_R input124 (.A(io_ins_down_1[63]),
    .Y(net124));
 BUFx2_ASAP7_75t_R input125 (.A(io_ins_down_1[6]),
    .Y(net125));
 BUFx2_ASAP7_75t_R input126 (.A(io_ins_down_1[7]),
    .Y(net126));
 BUFx2_ASAP7_75t_R input127 (.A(io_ins_down_1[8]),
    .Y(net127));
 BUFx2_ASAP7_75t_R input128 (.A(io_ins_down_1[9]),
    .Y(net128));
 BUFx2_ASAP7_75t_R input129 (.A(io_ins_down_2[0]),
    .Y(net129));
 BUFx2_ASAP7_75t_R input130 (.A(io_ins_down_2[10]),
    .Y(net130));
 BUFx2_ASAP7_75t_R input131 (.A(io_ins_down_2[11]),
    .Y(net131));
 BUFx2_ASAP7_75t_R input132 (.A(io_ins_down_2[12]),
    .Y(net132));
 BUFx2_ASAP7_75t_R input133 (.A(io_ins_down_2[13]),
    .Y(net133));
 BUFx2_ASAP7_75t_R input134 (.A(io_ins_down_2[14]),
    .Y(net134));
 BUFx2_ASAP7_75t_R input135 (.A(io_ins_down_2[15]),
    .Y(net135));
 BUFx2_ASAP7_75t_R input136 (.A(io_ins_down_2[16]),
    .Y(net136));
 BUFx2_ASAP7_75t_R input137 (.A(io_ins_down_2[17]),
    .Y(net137));
 BUFx2_ASAP7_75t_R input138 (.A(io_ins_down_2[18]),
    .Y(net138));
 BUFx2_ASAP7_75t_R input139 (.A(io_ins_down_2[19]),
    .Y(net139));
 BUFx2_ASAP7_75t_R input140 (.A(io_ins_down_2[1]),
    .Y(net140));
 BUFx2_ASAP7_75t_R input141 (.A(io_ins_down_2[20]),
    .Y(net141));
 BUFx2_ASAP7_75t_R input142 (.A(io_ins_down_2[21]),
    .Y(net142));
 BUFx2_ASAP7_75t_R input143 (.A(io_ins_down_2[22]),
    .Y(net143));
 BUFx2_ASAP7_75t_R input144 (.A(io_ins_down_2[23]),
    .Y(net144));
 BUFx2_ASAP7_75t_R input145 (.A(io_ins_down_2[24]),
    .Y(net145));
 BUFx2_ASAP7_75t_R input146 (.A(io_ins_down_2[25]),
    .Y(net146));
 BUFx2_ASAP7_75t_R input147 (.A(io_ins_down_2[26]),
    .Y(net147));
 BUFx2_ASAP7_75t_R input148 (.A(io_ins_down_2[27]),
    .Y(net148));
 BUFx2_ASAP7_75t_R input149 (.A(io_ins_down_2[28]),
    .Y(net149));
 BUFx2_ASAP7_75t_R input150 (.A(io_ins_down_2[29]),
    .Y(net150));
 BUFx2_ASAP7_75t_R input151 (.A(io_ins_down_2[2]),
    .Y(net151));
 BUFx2_ASAP7_75t_R input152 (.A(io_ins_down_2[30]),
    .Y(net152));
 BUFx2_ASAP7_75t_R input153 (.A(io_ins_down_2[31]),
    .Y(net153));
 BUFx2_ASAP7_75t_R input154 (.A(io_ins_down_2[32]),
    .Y(net154));
 BUFx2_ASAP7_75t_R input155 (.A(io_ins_down_2[33]),
    .Y(net155));
 BUFx2_ASAP7_75t_R input156 (.A(io_ins_down_2[34]),
    .Y(net156));
 BUFx2_ASAP7_75t_R input157 (.A(io_ins_down_2[35]),
    .Y(net157));
 BUFx2_ASAP7_75t_R input158 (.A(io_ins_down_2[36]),
    .Y(net158));
 BUFx2_ASAP7_75t_R input159 (.A(io_ins_down_2[37]),
    .Y(net159));
 BUFx2_ASAP7_75t_R input160 (.A(io_ins_down_2[38]),
    .Y(net160));
 BUFx2_ASAP7_75t_R input161 (.A(io_ins_down_2[39]),
    .Y(net161));
 BUFx2_ASAP7_75t_R input162 (.A(io_ins_down_2[3]),
    .Y(net162));
 BUFx2_ASAP7_75t_R input163 (.A(io_ins_down_2[40]),
    .Y(net163));
 BUFx2_ASAP7_75t_R input164 (.A(io_ins_down_2[41]),
    .Y(net164));
 BUFx2_ASAP7_75t_R input165 (.A(io_ins_down_2[42]),
    .Y(net165));
 BUFx2_ASAP7_75t_R input166 (.A(io_ins_down_2[43]),
    .Y(net166));
 BUFx2_ASAP7_75t_R input167 (.A(io_ins_down_2[44]),
    .Y(net167));
 BUFx2_ASAP7_75t_R input168 (.A(io_ins_down_2[45]),
    .Y(net168));
 BUFx2_ASAP7_75t_R input169 (.A(io_ins_down_2[46]),
    .Y(net169));
 BUFx2_ASAP7_75t_R input170 (.A(io_ins_down_2[47]),
    .Y(net170));
 BUFx2_ASAP7_75t_R input171 (.A(io_ins_down_2[48]),
    .Y(net171));
 BUFx2_ASAP7_75t_R input172 (.A(io_ins_down_2[49]),
    .Y(net172));
 BUFx2_ASAP7_75t_R input173 (.A(io_ins_down_2[4]),
    .Y(net173));
 BUFx2_ASAP7_75t_R input174 (.A(io_ins_down_2[50]),
    .Y(net174));
 BUFx2_ASAP7_75t_R input175 (.A(io_ins_down_2[51]),
    .Y(net175));
 BUFx2_ASAP7_75t_R input176 (.A(io_ins_down_2[52]),
    .Y(net176));
 BUFx2_ASAP7_75t_R input177 (.A(io_ins_down_2[53]),
    .Y(net177));
 BUFx2_ASAP7_75t_R input178 (.A(io_ins_down_2[54]),
    .Y(net178));
 BUFx2_ASAP7_75t_R input179 (.A(io_ins_down_2[55]),
    .Y(net179));
 BUFx2_ASAP7_75t_R input180 (.A(io_ins_down_2[56]),
    .Y(net180));
 BUFx2_ASAP7_75t_R input181 (.A(io_ins_down_2[57]),
    .Y(net181));
 BUFx2_ASAP7_75t_R input182 (.A(io_ins_down_2[58]),
    .Y(net182));
 BUFx2_ASAP7_75t_R input183 (.A(io_ins_down_2[59]),
    .Y(net183));
 BUFx2_ASAP7_75t_R input184 (.A(io_ins_down_2[5]),
    .Y(net184));
 BUFx2_ASAP7_75t_R input185 (.A(io_ins_down_2[60]),
    .Y(net185));
 BUFx2_ASAP7_75t_R input186 (.A(io_ins_down_2[61]),
    .Y(net186));
 BUFx2_ASAP7_75t_R input187 (.A(io_ins_down_2[62]),
    .Y(net187));
 BUFx2_ASAP7_75t_R input188 (.A(io_ins_down_2[63]),
    .Y(net188));
 BUFx2_ASAP7_75t_R input189 (.A(io_ins_down_2[6]),
    .Y(net189));
 BUFx2_ASAP7_75t_R input190 (.A(io_ins_down_2[7]),
    .Y(net190));
 BUFx2_ASAP7_75t_R input191 (.A(io_ins_down_2[8]),
    .Y(net191));
 BUFx2_ASAP7_75t_R input192 (.A(io_ins_down_2[9]),
    .Y(net192));
 BUFx2_ASAP7_75t_R input193 (.A(io_ins_down_3[0]),
    .Y(net193));
 BUFx2_ASAP7_75t_R input194 (.A(io_ins_down_3[10]),
    .Y(net194));
 BUFx2_ASAP7_75t_R input195 (.A(io_ins_down_3[11]),
    .Y(net195));
 BUFx2_ASAP7_75t_R input196 (.A(io_ins_down_3[12]),
    .Y(net196));
 BUFx2_ASAP7_75t_R input197 (.A(io_ins_down_3[13]),
    .Y(net197));
 BUFx2_ASAP7_75t_R input198 (.A(io_ins_down_3[14]),
    .Y(net198));
 BUFx2_ASAP7_75t_R input199 (.A(io_ins_down_3[15]),
    .Y(net199));
 BUFx2_ASAP7_75t_R input200 (.A(io_ins_down_3[16]),
    .Y(net200));
 BUFx2_ASAP7_75t_R input201 (.A(io_ins_down_3[17]),
    .Y(net201));
 BUFx2_ASAP7_75t_R input202 (.A(io_ins_down_3[18]),
    .Y(net202));
 BUFx2_ASAP7_75t_R input203 (.A(io_ins_down_3[19]),
    .Y(net203));
 BUFx2_ASAP7_75t_R input204 (.A(io_ins_down_3[1]),
    .Y(net204));
 BUFx2_ASAP7_75t_R input205 (.A(io_ins_down_3[20]),
    .Y(net205));
 BUFx2_ASAP7_75t_R input206 (.A(io_ins_down_3[21]),
    .Y(net206));
 BUFx2_ASAP7_75t_R input207 (.A(io_ins_down_3[22]),
    .Y(net207));
 BUFx2_ASAP7_75t_R input208 (.A(io_ins_down_3[23]),
    .Y(net208));
 BUFx2_ASAP7_75t_R input209 (.A(io_ins_down_3[24]),
    .Y(net209));
 BUFx2_ASAP7_75t_R input210 (.A(io_ins_down_3[25]),
    .Y(net210));
 BUFx2_ASAP7_75t_R input211 (.A(io_ins_down_3[26]),
    .Y(net211));
 BUFx2_ASAP7_75t_R input212 (.A(io_ins_down_3[27]),
    .Y(net212));
 BUFx2_ASAP7_75t_R input213 (.A(io_ins_down_3[28]),
    .Y(net213));
 BUFx2_ASAP7_75t_R input214 (.A(io_ins_down_3[29]),
    .Y(net214));
 BUFx2_ASAP7_75t_R input215 (.A(io_ins_down_3[2]),
    .Y(net215));
 BUFx2_ASAP7_75t_R input216 (.A(io_ins_down_3[30]),
    .Y(net216));
 BUFx2_ASAP7_75t_R input217 (.A(io_ins_down_3[31]),
    .Y(net217));
 BUFx2_ASAP7_75t_R input218 (.A(io_ins_down_3[32]),
    .Y(net218));
 BUFx2_ASAP7_75t_R input219 (.A(io_ins_down_3[33]),
    .Y(net219));
 BUFx2_ASAP7_75t_R input220 (.A(io_ins_down_3[34]),
    .Y(net220));
 BUFx2_ASAP7_75t_R input221 (.A(io_ins_down_3[35]),
    .Y(net221));
 BUFx2_ASAP7_75t_R input222 (.A(io_ins_down_3[36]),
    .Y(net222));
 BUFx2_ASAP7_75t_R input223 (.A(io_ins_down_3[37]),
    .Y(net223));
 BUFx2_ASAP7_75t_R input224 (.A(io_ins_down_3[38]),
    .Y(net224));
 BUFx2_ASAP7_75t_R input225 (.A(io_ins_down_3[39]),
    .Y(net225));
 BUFx2_ASAP7_75t_R input226 (.A(io_ins_down_3[3]),
    .Y(net226));
 BUFx2_ASAP7_75t_R input227 (.A(io_ins_down_3[40]),
    .Y(net227));
 BUFx2_ASAP7_75t_R input228 (.A(io_ins_down_3[41]),
    .Y(net228));
 BUFx2_ASAP7_75t_R input229 (.A(io_ins_down_3[42]),
    .Y(net229));
 BUFx2_ASAP7_75t_R input230 (.A(io_ins_down_3[43]),
    .Y(net230));
 BUFx2_ASAP7_75t_R input231 (.A(io_ins_down_3[44]),
    .Y(net231));
 BUFx2_ASAP7_75t_R input232 (.A(io_ins_down_3[45]),
    .Y(net232));
 BUFx2_ASAP7_75t_R input233 (.A(io_ins_down_3[46]),
    .Y(net233));
 BUFx2_ASAP7_75t_R input234 (.A(io_ins_down_3[47]),
    .Y(net234));
 BUFx2_ASAP7_75t_R input235 (.A(io_ins_down_3[48]),
    .Y(net235));
 BUFx2_ASAP7_75t_R input236 (.A(io_ins_down_3[49]),
    .Y(net236));
 BUFx2_ASAP7_75t_R input237 (.A(io_ins_down_3[4]),
    .Y(net237));
 BUFx2_ASAP7_75t_R input238 (.A(io_ins_down_3[50]),
    .Y(net238));
 BUFx2_ASAP7_75t_R input239 (.A(io_ins_down_3[51]),
    .Y(net239));
 BUFx2_ASAP7_75t_R input240 (.A(io_ins_down_3[52]),
    .Y(net240));
 BUFx2_ASAP7_75t_R input241 (.A(io_ins_down_3[53]),
    .Y(net241));
 BUFx2_ASAP7_75t_R input242 (.A(io_ins_down_3[54]),
    .Y(net242));
 BUFx2_ASAP7_75t_R input243 (.A(io_ins_down_3[55]),
    .Y(net243));
 BUFx2_ASAP7_75t_R input244 (.A(io_ins_down_3[56]),
    .Y(net244));
 BUFx2_ASAP7_75t_R input245 (.A(io_ins_down_3[57]),
    .Y(net245));
 BUFx2_ASAP7_75t_R input246 (.A(io_ins_down_3[58]),
    .Y(net246));
 BUFx2_ASAP7_75t_R input247 (.A(io_ins_down_3[59]),
    .Y(net247));
 BUFx2_ASAP7_75t_R input248 (.A(io_ins_down_3[5]),
    .Y(net248));
 BUFx2_ASAP7_75t_R input249 (.A(io_ins_down_3[60]),
    .Y(net249));
 BUFx2_ASAP7_75t_R input250 (.A(io_ins_down_3[61]),
    .Y(net250));
 BUFx2_ASAP7_75t_R input251 (.A(io_ins_down_3[62]),
    .Y(net251));
 BUFx2_ASAP7_75t_R input252 (.A(io_ins_down_3[63]),
    .Y(net252));
 BUFx2_ASAP7_75t_R input253 (.A(io_ins_down_3[6]),
    .Y(net253));
 BUFx2_ASAP7_75t_R input254 (.A(io_ins_down_3[7]),
    .Y(net254));
 BUFx2_ASAP7_75t_R input255 (.A(io_ins_down_3[8]),
    .Y(net255));
 BUFx2_ASAP7_75t_R input256 (.A(io_ins_down_3[9]),
    .Y(net256));
 BUFx2_ASAP7_75t_R input257 (.A(io_ins_down_4[0]),
    .Y(net257));
 BUFx2_ASAP7_75t_R input258 (.A(io_ins_down_4[10]),
    .Y(net258));
 BUFx2_ASAP7_75t_R input259 (.A(io_ins_down_4[11]),
    .Y(net259));
 BUFx2_ASAP7_75t_R input260 (.A(io_ins_down_4[12]),
    .Y(net260));
 BUFx2_ASAP7_75t_R input261 (.A(io_ins_down_4[13]),
    .Y(net261));
 BUFx2_ASAP7_75t_R input262 (.A(io_ins_down_4[14]),
    .Y(net262));
 BUFx2_ASAP7_75t_R input263 (.A(io_ins_down_4[15]),
    .Y(net263));
 BUFx2_ASAP7_75t_R input264 (.A(io_ins_down_4[16]),
    .Y(net264));
 BUFx2_ASAP7_75t_R input265 (.A(io_ins_down_4[17]),
    .Y(net265));
 BUFx2_ASAP7_75t_R input266 (.A(io_ins_down_4[18]),
    .Y(net266));
 BUFx2_ASAP7_75t_R input267 (.A(io_ins_down_4[19]),
    .Y(net267));
 BUFx2_ASAP7_75t_R input268 (.A(io_ins_down_4[1]),
    .Y(net268));
 BUFx2_ASAP7_75t_R input269 (.A(io_ins_down_4[20]),
    .Y(net269));
 BUFx2_ASAP7_75t_R input270 (.A(io_ins_down_4[21]),
    .Y(net270));
 BUFx2_ASAP7_75t_R input271 (.A(io_ins_down_4[22]),
    .Y(net271));
 BUFx2_ASAP7_75t_R input272 (.A(io_ins_down_4[23]),
    .Y(net272));
 BUFx2_ASAP7_75t_R input273 (.A(io_ins_down_4[24]),
    .Y(net273));
 BUFx2_ASAP7_75t_R input274 (.A(io_ins_down_4[25]),
    .Y(net274));
 BUFx2_ASAP7_75t_R input275 (.A(io_ins_down_4[26]),
    .Y(net275));
 BUFx2_ASAP7_75t_R input276 (.A(io_ins_down_4[27]),
    .Y(net276));
 BUFx2_ASAP7_75t_R input277 (.A(io_ins_down_4[28]),
    .Y(net277));
 BUFx2_ASAP7_75t_R input278 (.A(io_ins_down_4[29]),
    .Y(net278));
 BUFx2_ASAP7_75t_R input279 (.A(io_ins_down_4[2]),
    .Y(net279));
 BUFx2_ASAP7_75t_R input280 (.A(io_ins_down_4[30]),
    .Y(net280));
 BUFx2_ASAP7_75t_R input281 (.A(io_ins_down_4[31]),
    .Y(net281));
 BUFx2_ASAP7_75t_R input282 (.A(io_ins_down_4[32]),
    .Y(net282));
 BUFx2_ASAP7_75t_R input283 (.A(io_ins_down_4[33]),
    .Y(net283));
 BUFx2_ASAP7_75t_R input284 (.A(io_ins_down_4[34]),
    .Y(net284));
 BUFx2_ASAP7_75t_R input285 (.A(io_ins_down_4[35]),
    .Y(net285));
 BUFx2_ASAP7_75t_R input286 (.A(io_ins_down_4[36]),
    .Y(net286));
 BUFx2_ASAP7_75t_R input287 (.A(io_ins_down_4[37]),
    .Y(net287));
 BUFx2_ASAP7_75t_R input288 (.A(io_ins_down_4[38]),
    .Y(net288));
 BUFx2_ASAP7_75t_R input289 (.A(io_ins_down_4[39]),
    .Y(net289));
 BUFx2_ASAP7_75t_R input290 (.A(io_ins_down_4[3]),
    .Y(net290));
 BUFx2_ASAP7_75t_R input291 (.A(io_ins_down_4[40]),
    .Y(net291));
 BUFx2_ASAP7_75t_R input292 (.A(io_ins_down_4[41]),
    .Y(net292));
 BUFx2_ASAP7_75t_R input293 (.A(io_ins_down_4[42]),
    .Y(net293));
 BUFx2_ASAP7_75t_R input294 (.A(io_ins_down_4[43]),
    .Y(net294));
 BUFx2_ASAP7_75t_R input295 (.A(io_ins_down_4[44]),
    .Y(net295));
 BUFx2_ASAP7_75t_R input296 (.A(io_ins_down_4[45]),
    .Y(net296));
 BUFx2_ASAP7_75t_R input297 (.A(io_ins_down_4[46]),
    .Y(net297));
 BUFx2_ASAP7_75t_R input298 (.A(io_ins_down_4[47]),
    .Y(net298));
 BUFx2_ASAP7_75t_R input299 (.A(io_ins_down_4[48]),
    .Y(net299));
 BUFx2_ASAP7_75t_R input300 (.A(io_ins_down_4[49]),
    .Y(net300));
 BUFx2_ASAP7_75t_R input301 (.A(io_ins_down_4[4]),
    .Y(net301));
 BUFx2_ASAP7_75t_R input302 (.A(io_ins_down_4[50]),
    .Y(net302));
 BUFx2_ASAP7_75t_R input303 (.A(io_ins_down_4[51]),
    .Y(net303));
 BUFx2_ASAP7_75t_R input304 (.A(io_ins_down_4[52]),
    .Y(net304));
 BUFx2_ASAP7_75t_R input305 (.A(io_ins_down_4[53]),
    .Y(net305));
 BUFx2_ASAP7_75t_R input306 (.A(io_ins_down_4[54]),
    .Y(net306));
 BUFx2_ASAP7_75t_R input307 (.A(io_ins_down_4[55]),
    .Y(net307));
 BUFx2_ASAP7_75t_R input308 (.A(io_ins_down_4[56]),
    .Y(net308));
 BUFx2_ASAP7_75t_R input309 (.A(io_ins_down_4[57]),
    .Y(net309));
 BUFx2_ASAP7_75t_R input310 (.A(io_ins_down_4[58]),
    .Y(net310));
 BUFx2_ASAP7_75t_R input311 (.A(io_ins_down_4[59]),
    .Y(net311));
 BUFx2_ASAP7_75t_R input312 (.A(io_ins_down_4[5]),
    .Y(net312));
 BUFx2_ASAP7_75t_R input313 (.A(io_ins_down_4[60]),
    .Y(net313));
 BUFx2_ASAP7_75t_R input314 (.A(io_ins_down_4[61]),
    .Y(net314));
 BUFx2_ASAP7_75t_R input315 (.A(io_ins_down_4[62]),
    .Y(net315));
 BUFx2_ASAP7_75t_R input316 (.A(io_ins_down_4[63]),
    .Y(net316));
 BUFx2_ASAP7_75t_R input317 (.A(io_ins_down_4[6]),
    .Y(net317));
 BUFx2_ASAP7_75t_R input318 (.A(io_ins_down_4[7]),
    .Y(net318));
 BUFx2_ASAP7_75t_R input319 (.A(io_ins_down_4[8]),
    .Y(net319));
 BUFx2_ASAP7_75t_R input320 (.A(io_ins_down_4[9]),
    .Y(net320));
 BUFx2_ASAP7_75t_R input321 (.A(io_ins_down_5[0]),
    .Y(net321));
 BUFx2_ASAP7_75t_R input322 (.A(io_ins_down_5[10]),
    .Y(net322));
 BUFx2_ASAP7_75t_R input323 (.A(io_ins_down_5[11]),
    .Y(net323));
 BUFx2_ASAP7_75t_R input324 (.A(io_ins_down_5[12]),
    .Y(net324));
 BUFx2_ASAP7_75t_R input325 (.A(io_ins_down_5[13]),
    .Y(net325));
 BUFx2_ASAP7_75t_R input326 (.A(io_ins_down_5[14]),
    .Y(net326));
 BUFx2_ASAP7_75t_R input327 (.A(io_ins_down_5[15]),
    .Y(net327));
 BUFx2_ASAP7_75t_R input328 (.A(io_ins_down_5[16]),
    .Y(net328));
 BUFx2_ASAP7_75t_R input329 (.A(io_ins_down_5[17]),
    .Y(net329));
 BUFx2_ASAP7_75t_R input330 (.A(io_ins_down_5[18]),
    .Y(net330));
 BUFx2_ASAP7_75t_R input331 (.A(io_ins_down_5[19]),
    .Y(net331));
 BUFx2_ASAP7_75t_R input332 (.A(io_ins_down_5[1]),
    .Y(net332));
 BUFx2_ASAP7_75t_R input333 (.A(io_ins_down_5[20]),
    .Y(net333));
 BUFx2_ASAP7_75t_R input334 (.A(io_ins_down_5[21]),
    .Y(net334));
 BUFx2_ASAP7_75t_R input335 (.A(io_ins_down_5[22]),
    .Y(net335));
 BUFx2_ASAP7_75t_R input336 (.A(io_ins_down_5[23]),
    .Y(net336));
 BUFx2_ASAP7_75t_R input337 (.A(io_ins_down_5[24]),
    .Y(net337));
 BUFx2_ASAP7_75t_R input338 (.A(io_ins_down_5[25]),
    .Y(net338));
 BUFx2_ASAP7_75t_R input339 (.A(io_ins_down_5[26]),
    .Y(net339));
 BUFx2_ASAP7_75t_R input340 (.A(io_ins_down_5[27]),
    .Y(net340));
 BUFx2_ASAP7_75t_R input341 (.A(io_ins_down_5[28]),
    .Y(net341));
 BUFx2_ASAP7_75t_R input342 (.A(io_ins_down_5[29]),
    .Y(net342));
 BUFx2_ASAP7_75t_R input343 (.A(io_ins_down_5[2]),
    .Y(net343));
 BUFx2_ASAP7_75t_R input344 (.A(io_ins_down_5[30]),
    .Y(net344));
 BUFx2_ASAP7_75t_R input345 (.A(io_ins_down_5[31]),
    .Y(net345));
 BUFx2_ASAP7_75t_R input346 (.A(io_ins_down_5[32]),
    .Y(net346));
 BUFx2_ASAP7_75t_R input347 (.A(io_ins_down_5[33]),
    .Y(net347));
 BUFx2_ASAP7_75t_R input348 (.A(io_ins_down_5[34]),
    .Y(net348));
 BUFx2_ASAP7_75t_R input349 (.A(io_ins_down_5[35]),
    .Y(net349));
 BUFx2_ASAP7_75t_R input350 (.A(io_ins_down_5[36]),
    .Y(net350));
 BUFx2_ASAP7_75t_R input351 (.A(io_ins_down_5[37]),
    .Y(net351));
 BUFx2_ASAP7_75t_R input352 (.A(io_ins_down_5[38]),
    .Y(net352));
 BUFx2_ASAP7_75t_R input353 (.A(io_ins_down_5[39]),
    .Y(net353));
 BUFx2_ASAP7_75t_R input354 (.A(io_ins_down_5[3]),
    .Y(net354));
 BUFx2_ASAP7_75t_R input355 (.A(io_ins_down_5[40]),
    .Y(net355));
 BUFx2_ASAP7_75t_R input356 (.A(io_ins_down_5[41]),
    .Y(net356));
 BUFx2_ASAP7_75t_R input357 (.A(io_ins_down_5[42]),
    .Y(net357));
 BUFx2_ASAP7_75t_R input358 (.A(io_ins_down_5[43]),
    .Y(net358));
 BUFx2_ASAP7_75t_R input359 (.A(io_ins_down_5[44]),
    .Y(net359));
 BUFx2_ASAP7_75t_R input360 (.A(io_ins_down_5[45]),
    .Y(net360));
 BUFx2_ASAP7_75t_R input361 (.A(io_ins_down_5[46]),
    .Y(net361));
 BUFx2_ASAP7_75t_R input362 (.A(io_ins_down_5[47]),
    .Y(net362));
 BUFx2_ASAP7_75t_R input363 (.A(io_ins_down_5[48]),
    .Y(net363));
 BUFx2_ASAP7_75t_R input364 (.A(io_ins_down_5[49]),
    .Y(net364));
 BUFx2_ASAP7_75t_R input365 (.A(io_ins_down_5[4]),
    .Y(net365));
 BUFx2_ASAP7_75t_R input366 (.A(io_ins_down_5[50]),
    .Y(net366));
 BUFx2_ASAP7_75t_R input367 (.A(io_ins_down_5[51]),
    .Y(net367));
 BUFx2_ASAP7_75t_R input368 (.A(io_ins_down_5[52]),
    .Y(net368));
 BUFx2_ASAP7_75t_R input369 (.A(io_ins_down_5[53]),
    .Y(net369));
 BUFx2_ASAP7_75t_R input370 (.A(io_ins_down_5[54]),
    .Y(net370));
 BUFx2_ASAP7_75t_R input371 (.A(io_ins_down_5[55]),
    .Y(net371));
 BUFx2_ASAP7_75t_R input372 (.A(io_ins_down_5[56]),
    .Y(net372));
 BUFx2_ASAP7_75t_R input373 (.A(io_ins_down_5[57]),
    .Y(net373));
 BUFx2_ASAP7_75t_R input374 (.A(io_ins_down_5[58]),
    .Y(net374));
 BUFx2_ASAP7_75t_R input375 (.A(io_ins_down_5[59]),
    .Y(net375));
 BUFx2_ASAP7_75t_R input376 (.A(io_ins_down_5[5]),
    .Y(net376));
 BUFx2_ASAP7_75t_R input377 (.A(io_ins_down_5[60]),
    .Y(net377));
 BUFx2_ASAP7_75t_R input378 (.A(io_ins_down_5[61]),
    .Y(net378));
 BUFx2_ASAP7_75t_R input379 (.A(io_ins_down_5[62]),
    .Y(net379));
 BUFx2_ASAP7_75t_R input380 (.A(io_ins_down_5[63]),
    .Y(net380));
 BUFx2_ASAP7_75t_R input381 (.A(io_ins_down_5[6]),
    .Y(net381));
 BUFx2_ASAP7_75t_R input382 (.A(io_ins_down_5[7]),
    .Y(net382));
 BUFx2_ASAP7_75t_R input383 (.A(io_ins_down_5[8]),
    .Y(net383));
 BUFx2_ASAP7_75t_R input384 (.A(io_ins_down_5[9]),
    .Y(net384));
 BUFx2_ASAP7_75t_R input385 (.A(io_ins_down_6[0]),
    .Y(net385));
 BUFx2_ASAP7_75t_R input386 (.A(io_ins_down_6[10]),
    .Y(net386));
 BUFx2_ASAP7_75t_R input387 (.A(io_ins_down_6[11]),
    .Y(net387));
 BUFx2_ASAP7_75t_R input388 (.A(io_ins_down_6[12]),
    .Y(net388));
 BUFx2_ASAP7_75t_R input389 (.A(io_ins_down_6[13]),
    .Y(net389));
 BUFx2_ASAP7_75t_R input390 (.A(io_ins_down_6[14]),
    .Y(net390));
 BUFx2_ASAP7_75t_R input391 (.A(io_ins_down_6[15]),
    .Y(net391));
 BUFx2_ASAP7_75t_R input392 (.A(io_ins_down_6[16]),
    .Y(net392));
 BUFx2_ASAP7_75t_R input393 (.A(io_ins_down_6[17]),
    .Y(net393));
 BUFx2_ASAP7_75t_R input394 (.A(io_ins_down_6[18]),
    .Y(net394));
 BUFx2_ASAP7_75t_R input395 (.A(io_ins_down_6[19]),
    .Y(net395));
 BUFx2_ASAP7_75t_R input396 (.A(io_ins_down_6[1]),
    .Y(net396));
 BUFx2_ASAP7_75t_R input397 (.A(io_ins_down_6[20]),
    .Y(net397));
 BUFx2_ASAP7_75t_R input398 (.A(io_ins_down_6[21]),
    .Y(net398));
 BUFx2_ASAP7_75t_R input399 (.A(io_ins_down_6[22]),
    .Y(net399));
 BUFx2_ASAP7_75t_R input400 (.A(io_ins_down_6[23]),
    .Y(net400));
 BUFx2_ASAP7_75t_R input401 (.A(io_ins_down_6[24]),
    .Y(net401));
 BUFx2_ASAP7_75t_R input402 (.A(io_ins_down_6[25]),
    .Y(net402));
 BUFx2_ASAP7_75t_R input403 (.A(io_ins_down_6[26]),
    .Y(net403));
 BUFx2_ASAP7_75t_R input404 (.A(io_ins_down_6[27]),
    .Y(net404));
 BUFx2_ASAP7_75t_R input405 (.A(io_ins_down_6[28]),
    .Y(net405));
 BUFx2_ASAP7_75t_R input406 (.A(io_ins_down_6[29]),
    .Y(net406));
 BUFx2_ASAP7_75t_R input407 (.A(io_ins_down_6[2]),
    .Y(net407));
 BUFx2_ASAP7_75t_R input408 (.A(io_ins_down_6[30]),
    .Y(net408));
 BUFx2_ASAP7_75t_R input409 (.A(io_ins_down_6[31]),
    .Y(net409));
 BUFx2_ASAP7_75t_R input410 (.A(io_ins_down_6[32]),
    .Y(net410));
 BUFx2_ASAP7_75t_R input411 (.A(io_ins_down_6[33]),
    .Y(net411));
 BUFx2_ASAP7_75t_R input412 (.A(io_ins_down_6[34]),
    .Y(net412));
 BUFx2_ASAP7_75t_R input413 (.A(io_ins_down_6[35]),
    .Y(net413));
 BUFx2_ASAP7_75t_R input414 (.A(io_ins_down_6[36]),
    .Y(net414));
 BUFx2_ASAP7_75t_R input415 (.A(io_ins_down_6[37]),
    .Y(net415));
 BUFx2_ASAP7_75t_R input416 (.A(io_ins_down_6[38]),
    .Y(net416));
 BUFx2_ASAP7_75t_R input417 (.A(io_ins_down_6[39]),
    .Y(net417));
 BUFx2_ASAP7_75t_R input418 (.A(io_ins_down_6[3]),
    .Y(net418));
 BUFx2_ASAP7_75t_R input419 (.A(io_ins_down_6[40]),
    .Y(net419));
 BUFx2_ASAP7_75t_R input420 (.A(io_ins_down_6[41]),
    .Y(net420));
 BUFx2_ASAP7_75t_R input421 (.A(io_ins_down_6[42]),
    .Y(net421));
 BUFx2_ASAP7_75t_R input422 (.A(io_ins_down_6[43]),
    .Y(net422));
 BUFx2_ASAP7_75t_R input423 (.A(io_ins_down_6[44]),
    .Y(net423));
 BUFx2_ASAP7_75t_R input424 (.A(io_ins_down_6[45]),
    .Y(net424));
 BUFx2_ASAP7_75t_R input425 (.A(io_ins_down_6[46]),
    .Y(net425));
 BUFx2_ASAP7_75t_R input426 (.A(io_ins_down_6[47]),
    .Y(net426));
 BUFx2_ASAP7_75t_R input427 (.A(io_ins_down_6[48]),
    .Y(net427));
 BUFx2_ASAP7_75t_R input428 (.A(io_ins_down_6[49]),
    .Y(net428));
 BUFx2_ASAP7_75t_R input429 (.A(io_ins_down_6[4]),
    .Y(net429));
 BUFx2_ASAP7_75t_R input430 (.A(io_ins_down_6[50]),
    .Y(net430));
 BUFx2_ASAP7_75t_R input431 (.A(io_ins_down_6[51]),
    .Y(net431));
 BUFx2_ASAP7_75t_R input432 (.A(io_ins_down_6[52]),
    .Y(net432));
 BUFx2_ASAP7_75t_R input433 (.A(io_ins_down_6[53]),
    .Y(net433));
 BUFx2_ASAP7_75t_R input434 (.A(io_ins_down_6[54]),
    .Y(net434));
 BUFx2_ASAP7_75t_R input435 (.A(io_ins_down_6[55]),
    .Y(net435));
 BUFx2_ASAP7_75t_R input436 (.A(io_ins_down_6[56]),
    .Y(net436));
 BUFx2_ASAP7_75t_R input437 (.A(io_ins_down_6[57]),
    .Y(net437));
 BUFx2_ASAP7_75t_R input438 (.A(io_ins_down_6[58]),
    .Y(net438));
 BUFx2_ASAP7_75t_R input439 (.A(io_ins_down_6[59]),
    .Y(net439));
 BUFx2_ASAP7_75t_R input440 (.A(io_ins_down_6[5]),
    .Y(net440));
 BUFx2_ASAP7_75t_R input441 (.A(io_ins_down_6[60]),
    .Y(net441));
 BUFx2_ASAP7_75t_R input442 (.A(io_ins_down_6[61]),
    .Y(net442));
 BUFx2_ASAP7_75t_R input443 (.A(io_ins_down_6[62]),
    .Y(net443));
 BUFx2_ASAP7_75t_R input444 (.A(io_ins_down_6[63]),
    .Y(net444));
 BUFx2_ASAP7_75t_R input445 (.A(io_ins_down_6[6]),
    .Y(net445));
 BUFx2_ASAP7_75t_R input446 (.A(io_ins_down_6[7]),
    .Y(net446));
 BUFx2_ASAP7_75t_R input447 (.A(io_ins_down_6[8]),
    .Y(net447));
 BUFx2_ASAP7_75t_R input448 (.A(io_ins_down_6[9]),
    .Y(net448));
 BUFx2_ASAP7_75t_R input449 (.A(io_ins_down_7[0]),
    .Y(net449));
 BUFx2_ASAP7_75t_R input450 (.A(io_ins_down_7[10]),
    .Y(net450));
 BUFx2_ASAP7_75t_R input451 (.A(io_ins_down_7[11]),
    .Y(net451));
 BUFx2_ASAP7_75t_R input452 (.A(io_ins_down_7[12]),
    .Y(net452));
 BUFx2_ASAP7_75t_R input453 (.A(io_ins_down_7[13]),
    .Y(net453));
 BUFx2_ASAP7_75t_R input454 (.A(io_ins_down_7[14]),
    .Y(net454));
 BUFx2_ASAP7_75t_R input455 (.A(io_ins_down_7[15]),
    .Y(net455));
 BUFx2_ASAP7_75t_R input456 (.A(io_ins_down_7[16]),
    .Y(net456));
 BUFx2_ASAP7_75t_R input457 (.A(io_ins_down_7[17]),
    .Y(net457));
 BUFx2_ASAP7_75t_R input458 (.A(io_ins_down_7[18]),
    .Y(net458));
 BUFx2_ASAP7_75t_R input459 (.A(io_ins_down_7[19]),
    .Y(net459));
 BUFx2_ASAP7_75t_R input460 (.A(io_ins_down_7[1]),
    .Y(net460));
 BUFx2_ASAP7_75t_R input461 (.A(io_ins_down_7[20]),
    .Y(net461));
 BUFx2_ASAP7_75t_R input462 (.A(io_ins_down_7[21]),
    .Y(net462));
 BUFx2_ASAP7_75t_R input463 (.A(io_ins_down_7[22]),
    .Y(net463));
 BUFx2_ASAP7_75t_R input464 (.A(io_ins_down_7[23]),
    .Y(net464));
 BUFx2_ASAP7_75t_R input465 (.A(io_ins_down_7[24]),
    .Y(net465));
 BUFx2_ASAP7_75t_R input466 (.A(io_ins_down_7[25]),
    .Y(net466));
 BUFx2_ASAP7_75t_R input467 (.A(io_ins_down_7[26]),
    .Y(net467));
 BUFx2_ASAP7_75t_R input468 (.A(io_ins_down_7[27]),
    .Y(net468));
 BUFx2_ASAP7_75t_R input469 (.A(io_ins_down_7[28]),
    .Y(net469));
 BUFx2_ASAP7_75t_R input470 (.A(io_ins_down_7[29]),
    .Y(net470));
 BUFx2_ASAP7_75t_R input471 (.A(io_ins_down_7[2]),
    .Y(net471));
 BUFx2_ASAP7_75t_R input472 (.A(io_ins_down_7[30]),
    .Y(net472));
 BUFx2_ASAP7_75t_R input473 (.A(io_ins_down_7[31]),
    .Y(net473));
 BUFx2_ASAP7_75t_R input474 (.A(io_ins_down_7[32]),
    .Y(net474));
 BUFx2_ASAP7_75t_R input475 (.A(io_ins_down_7[33]),
    .Y(net475));
 BUFx2_ASAP7_75t_R input476 (.A(io_ins_down_7[34]),
    .Y(net476));
 BUFx2_ASAP7_75t_R input477 (.A(io_ins_down_7[35]),
    .Y(net477));
 BUFx2_ASAP7_75t_R input478 (.A(io_ins_down_7[36]),
    .Y(net478));
 BUFx2_ASAP7_75t_R input479 (.A(io_ins_down_7[37]),
    .Y(net479));
 BUFx2_ASAP7_75t_R input480 (.A(io_ins_down_7[38]),
    .Y(net480));
 BUFx2_ASAP7_75t_R input481 (.A(io_ins_down_7[39]),
    .Y(net481));
 BUFx2_ASAP7_75t_R input482 (.A(io_ins_down_7[3]),
    .Y(net482));
 BUFx2_ASAP7_75t_R input483 (.A(io_ins_down_7[40]),
    .Y(net483));
 BUFx2_ASAP7_75t_R input484 (.A(io_ins_down_7[41]),
    .Y(net484));
 BUFx2_ASAP7_75t_R input485 (.A(io_ins_down_7[42]),
    .Y(net485));
 BUFx2_ASAP7_75t_R input486 (.A(io_ins_down_7[43]),
    .Y(net486));
 BUFx2_ASAP7_75t_R input487 (.A(io_ins_down_7[44]),
    .Y(net487));
 BUFx2_ASAP7_75t_R input488 (.A(io_ins_down_7[45]),
    .Y(net488));
 BUFx2_ASAP7_75t_R input489 (.A(io_ins_down_7[46]),
    .Y(net489));
 BUFx2_ASAP7_75t_R input490 (.A(io_ins_down_7[47]),
    .Y(net490));
 BUFx2_ASAP7_75t_R input491 (.A(io_ins_down_7[48]),
    .Y(net491));
 BUFx2_ASAP7_75t_R input492 (.A(io_ins_down_7[49]),
    .Y(net492));
 BUFx2_ASAP7_75t_R input493 (.A(io_ins_down_7[4]),
    .Y(net493));
 BUFx2_ASAP7_75t_R input494 (.A(io_ins_down_7[50]),
    .Y(net494));
 BUFx2_ASAP7_75t_R input495 (.A(io_ins_down_7[51]),
    .Y(net495));
 BUFx2_ASAP7_75t_R input496 (.A(io_ins_down_7[52]),
    .Y(net496));
 BUFx2_ASAP7_75t_R input497 (.A(io_ins_down_7[53]),
    .Y(net497));
 BUFx2_ASAP7_75t_R input498 (.A(io_ins_down_7[54]),
    .Y(net498));
 BUFx2_ASAP7_75t_R input499 (.A(io_ins_down_7[55]),
    .Y(net499));
 BUFx2_ASAP7_75t_R input500 (.A(io_ins_down_7[56]),
    .Y(net500));
 BUFx2_ASAP7_75t_R input501 (.A(io_ins_down_7[57]),
    .Y(net501));
 BUFx2_ASAP7_75t_R input502 (.A(io_ins_down_7[58]),
    .Y(net502));
 BUFx2_ASAP7_75t_R input503 (.A(io_ins_down_7[59]),
    .Y(net503));
 BUFx2_ASAP7_75t_R input504 (.A(io_ins_down_7[5]),
    .Y(net504));
 BUFx2_ASAP7_75t_R input505 (.A(io_ins_down_7[60]),
    .Y(net505));
 BUFx2_ASAP7_75t_R input506 (.A(io_ins_down_7[61]),
    .Y(net506));
 BUFx2_ASAP7_75t_R input507 (.A(io_ins_down_7[62]),
    .Y(net507));
 BUFx2_ASAP7_75t_R input508 (.A(io_ins_down_7[63]),
    .Y(net508));
 BUFx2_ASAP7_75t_R input509 (.A(io_ins_down_7[6]),
    .Y(net509));
 BUFx2_ASAP7_75t_R input510 (.A(io_ins_down_7[7]),
    .Y(net510));
 BUFx2_ASAP7_75t_R input511 (.A(io_ins_down_7[8]),
    .Y(net511));
 BUFx2_ASAP7_75t_R input512 (.A(io_ins_down_7[9]),
    .Y(net512));
 BUFx2_ASAP7_75t_R input513 (.A(io_ins_left_0[0]),
    .Y(net513));
 BUFx2_ASAP7_75t_R input514 (.A(io_ins_left_0[10]),
    .Y(net514));
 BUFx2_ASAP7_75t_R input515 (.A(io_ins_left_0[11]),
    .Y(net515));
 BUFx2_ASAP7_75t_R input516 (.A(io_ins_left_0[12]),
    .Y(net516));
 BUFx2_ASAP7_75t_R input517 (.A(io_ins_left_0[13]),
    .Y(net517));
 BUFx2_ASAP7_75t_R input518 (.A(io_ins_left_0[14]),
    .Y(net518));
 BUFx2_ASAP7_75t_R input519 (.A(io_ins_left_0[15]),
    .Y(net519));
 BUFx2_ASAP7_75t_R input520 (.A(io_ins_left_0[16]),
    .Y(net520));
 BUFx2_ASAP7_75t_R input521 (.A(io_ins_left_0[17]),
    .Y(net521));
 BUFx2_ASAP7_75t_R input522 (.A(io_ins_left_0[18]),
    .Y(net522));
 BUFx2_ASAP7_75t_R input523 (.A(io_ins_left_0[19]),
    .Y(net523));
 BUFx2_ASAP7_75t_R input524 (.A(io_ins_left_0[1]),
    .Y(net524));
 BUFx2_ASAP7_75t_R input525 (.A(io_ins_left_0[20]),
    .Y(net525));
 BUFx2_ASAP7_75t_R input526 (.A(io_ins_left_0[21]),
    .Y(net526));
 BUFx2_ASAP7_75t_R input527 (.A(io_ins_left_0[22]),
    .Y(net527));
 BUFx2_ASAP7_75t_R input528 (.A(io_ins_left_0[23]),
    .Y(net528));
 BUFx2_ASAP7_75t_R input529 (.A(io_ins_left_0[24]),
    .Y(net529));
 BUFx2_ASAP7_75t_R input530 (.A(io_ins_left_0[25]),
    .Y(net530));
 BUFx2_ASAP7_75t_R input531 (.A(io_ins_left_0[26]),
    .Y(net531));
 BUFx2_ASAP7_75t_R input532 (.A(io_ins_left_0[27]),
    .Y(net532));
 BUFx2_ASAP7_75t_R input533 (.A(io_ins_left_0[28]),
    .Y(net533));
 BUFx2_ASAP7_75t_R input534 (.A(io_ins_left_0[29]),
    .Y(net534));
 BUFx2_ASAP7_75t_R input535 (.A(io_ins_left_0[2]),
    .Y(net535));
 BUFx2_ASAP7_75t_R input536 (.A(io_ins_left_0[30]),
    .Y(net536));
 BUFx2_ASAP7_75t_R input537 (.A(io_ins_left_0[31]),
    .Y(net537));
 BUFx2_ASAP7_75t_R input538 (.A(io_ins_left_0[32]),
    .Y(net538));
 BUFx2_ASAP7_75t_R input539 (.A(io_ins_left_0[33]),
    .Y(net539));
 BUFx2_ASAP7_75t_R input540 (.A(io_ins_left_0[34]),
    .Y(net540));
 BUFx2_ASAP7_75t_R input541 (.A(io_ins_left_0[35]),
    .Y(net541));
 BUFx2_ASAP7_75t_R input542 (.A(io_ins_left_0[36]),
    .Y(net542));
 BUFx2_ASAP7_75t_R input543 (.A(io_ins_left_0[37]),
    .Y(net543));
 BUFx2_ASAP7_75t_R input544 (.A(io_ins_left_0[38]),
    .Y(net544));
 BUFx2_ASAP7_75t_R input545 (.A(io_ins_left_0[39]),
    .Y(net545));
 BUFx2_ASAP7_75t_R input546 (.A(io_ins_left_0[3]),
    .Y(net546));
 BUFx2_ASAP7_75t_R input547 (.A(io_ins_left_0[40]),
    .Y(net547));
 BUFx2_ASAP7_75t_R input548 (.A(io_ins_left_0[41]),
    .Y(net548));
 BUFx2_ASAP7_75t_R input549 (.A(io_ins_left_0[42]),
    .Y(net549));
 BUFx2_ASAP7_75t_R input550 (.A(io_ins_left_0[43]),
    .Y(net550));
 BUFx2_ASAP7_75t_R input551 (.A(io_ins_left_0[44]),
    .Y(net551));
 BUFx2_ASAP7_75t_R input552 (.A(io_ins_left_0[45]),
    .Y(net552));
 BUFx2_ASAP7_75t_R input553 (.A(io_ins_left_0[46]),
    .Y(net553));
 BUFx2_ASAP7_75t_R input554 (.A(io_ins_left_0[47]),
    .Y(net554));
 BUFx2_ASAP7_75t_R input555 (.A(io_ins_left_0[48]),
    .Y(net555));
 BUFx2_ASAP7_75t_R input556 (.A(io_ins_left_0[49]),
    .Y(net556));
 BUFx2_ASAP7_75t_R input557 (.A(io_ins_left_0[4]),
    .Y(net557));
 BUFx2_ASAP7_75t_R input558 (.A(io_ins_left_0[50]),
    .Y(net558));
 BUFx2_ASAP7_75t_R input559 (.A(io_ins_left_0[51]),
    .Y(net559));
 BUFx2_ASAP7_75t_R input560 (.A(io_ins_left_0[52]),
    .Y(net560));
 BUFx2_ASAP7_75t_R input561 (.A(io_ins_left_0[53]),
    .Y(net561));
 BUFx2_ASAP7_75t_R input562 (.A(io_ins_left_0[54]),
    .Y(net562));
 BUFx2_ASAP7_75t_R input563 (.A(io_ins_left_0[55]),
    .Y(net563));
 BUFx2_ASAP7_75t_R input564 (.A(io_ins_left_0[56]),
    .Y(net564));
 BUFx2_ASAP7_75t_R input565 (.A(io_ins_left_0[57]),
    .Y(net565));
 BUFx2_ASAP7_75t_R input566 (.A(io_ins_left_0[58]),
    .Y(net566));
 BUFx2_ASAP7_75t_R input567 (.A(io_ins_left_0[59]),
    .Y(net567));
 BUFx2_ASAP7_75t_R input568 (.A(io_ins_left_0[5]),
    .Y(net568));
 BUFx2_ASAP7_75t_R input569 (.A(io_ins_left_0[60]),
    .Y(net569));
 BUFx2_ASAP7_75t_R input570 (.A(io_ins_left_0[61]),
    .Y(net570));
 BUFx2_ASAP7_75t_R input571 (.A(io_ins_left_0[62]),
    .Y(net571));
 BUFx2_ASAP7_75t_R input572 (.A(io_ins_left_0[63]),
    .Y(net572));
 BUFx2_ASAP7_75t_R input573 (.A(io_ins_left_0[6]),
    .Y(net573));
 BUFx2_ASAP7_75t_R input574 (.A(io_ins_left_0[7]),
    .Y(net574));
 BUFx2_ASAP7_75t_R input575 (.A(io_ins_left_0[8]),
    .Y(net575));
 BUFx2_ASAP7_75t_R input576 (.A(io_ins_left_0[9]),
    .Y(net576));
 BUFx2_ASAP7_75t_R input577 (.A(io_ins_left_1[0]),
    .Y(net577));
 BUFx2_ASAP7_75t_R input578 (.A(io_ins_left_1[10]),
    .Y(net578));
 BUFx2_ASAP7_75t_R input579 (.A(io_ins_left_1[11]),
    .Y(net579));
 BUFx2_ASAP7_75t_R input580 (.A(io_ins_left_1[12]),
    .Y(net580));
 BUFx2_ASAP7_75t_R input581 (.A(io_ins_left_1[13]),
    .Y(net581));
 BUFx2_ASAP7_75t_R input582 (.A(io_ins_left_1[14]),
    .Y(net582));
 BUFx2_ASAP7_75t_R input583 (.A(io_ins_left_1[15]),
    .Y(net583));
 BUFx2_ASAP7_75t_R input584 (.A(io_ins_left_1[16]),
    .Y(net584));
 BUFx2_ASAP7_75t_R input585 (.A(io_ins_left_1[17]),
    .Y(net585));
 BUFx2_ASAP7_75t_R input586 (.A(io_ins_left_1[18]),
    .Y(net586));
 BUFx2_ASAP7_75t_R input587 (.A(io_ins_left_1[19]),
    .Y(net587));
 BUFx2_ASAP7_75t_R input588 (.A(io_ins_left_1[1]),
    .Y(net588));
 BUFx2_ASAP7_75t_R input589 (.A(io_ins_left_1[20]),
    .Y(net589));
 BUFx2_ASAP7_75t_R input590 (.A(io_ins_left_1[21]),
    .Y(net590));
 BUFx2_ASAP7_75t_R input591 (.A(io_ins_left_1[22]),
    .Y(net591));
 BUFx2_ASAP7_75t_R input592 (.A(io_ins_left_1[23]),
    .Y(net592));
 BUFx2_ASAP7_75t_R input593 (.A(io_ins_left_1[24]),
    .Y(net593));
 BUFx2_ASAP7_75t_R input594 (.A(io_ins_left_1[25]),
    .Y(net594));
 BUFx2_ASAP7_75t_R input595 (.A(io_ins_left_1[26]),
    .Y(net595));
 BUFx2_ASAP7_75t_R input596 (.A(io_ins_left_1[27]),
    .Y(net596));
 BUFx2_ASAP7_75t_R input597 (.A(io_ins_left_1[28]),
    .Y(net597));
 BUFx2_ASAP7_75t_R input598 (.A(io_ins_left_1[29]),
    .Y(net598));
 BUFx2_ASAP7_75t_R input599 (.A(io_ins_left_1[2]),
    .Y(net599));
 BUFx2_ASAP7_75t_R input600 (.A(io_ins_left_1[30]),
    .Y(net600));
 BUFx2_ASAP7_75t_R input601 (.A(io_ins_left_1[31]),
    .Y(net601));
 BUFx2_ASAP7_75t_R input602 (.A(io_ins_left_1[32]),
    .Y(net602));
 BUFx2_ASAP7_75t_R input603 (.A(io_ins_left_1[33]),
    .Y(net603));
 BUFx2_ASAP7_75t_R input604 (.A(io_ins_left_1[34]),
    .Y(net604));
 BUFx2_ASAP7_75t_R input605 (.A(io_ins_left_1[35]),
    .Y(net605));
 BUFx2_ASAP7_75t_R input606 (.A(io_ins_left_1[36]),
    .Y(net606));
 BUFx2_ASAP7_75t_R input607 (.A(io_ins_left_1[37]),
    .Y(net607));
 BUFx2_ASAP7_75t_R input608 (.A(io_ins_left_1[38]),
    .Y(net608));
 BUFx2_ASAP7_75t_R input609 (.A(io_ins_left_1[39]),
    .Y(net609));
 BUFx2_ASAP7_75t_R input610 (.A(io_ins_left_1[3]),
    .Y(net610));
 BUFx2_ASAP7_75t_R input611 (.A(io_ins_left_1[40]),
    .Y(net611));
 BUFx2_ASAP7_75t_R input612 (.A(io_ins_left_1[41]),
    .Y(net612));
 BUFx2_ASAP7_75t_R input613 (.A(io_ins_left_1[42]),
    .Y(net613));
 BUFx2_ASAP7_75t_R input614 (.A(io_ins_left_1[43]),
    .Y(net614));
 BUFx2_ASAP7_75t_R input615 (.A(io_ins_left_1[44]),
    .Y(net615));
 BUFx2_ASAP7_75t_R input616 (.A(io_ins_left_1[45]),
    .Y(net616));
 BUFx2_ASAP7_75t_R input617 (.A(io_ins_left_1[46]),
    .Y(net617));
 BUFx2_ASAP7_75t_R input618 (.A(io_ins_left_1[47]),
    .Y(net618));
 BUFx2_ASAP7_75t_R input619 (.A(io_ins_left_1[48]),
    .Y(net619));
 BUFx2_ASAP7_75t_R input620 (.A(io_ins_left_1[49]),
    .Y(net620));
 BUFx2_ASAP7_75t_R input621 (.A(io_ins_left_1[4]),
    .Y(net621));
 BUFx2_ASAP7_75t_R input622 (.A(io_ins_left_1[50]),
    .Y(net622));
 BUFx2_ASAP7_75t_R input623 (.A(io_ins_left_1[51]),
    .Y(net623));
 BUFx2_ASAP7_75t_R input624 (.A(io_ins_left_1[52]),
    .Y(net624));
 BUFx2_ASAP7_75t_R input625 (.A(io_ins_left_1[53]),
    .Y(net625));
 BUFx2_ASAP7_75t_R input626 (.A(io_ins_left_1[54]),
    .Y(net626));
 BUFx2_ASAP7_75t_R input627 (.A(io_ins_left_1[55]),
    .Y(net627));
 BUFx2_ASAP7_75t_R input628 (.A(io_ins_left_1[56]),
    .Y(net628));
 BUFx2_ASAP7_75t_R input629 (.A(io_ins_left_1[57]),
    .Y(net629));
 BUFx2_ASAP7_75t_R input630 (.A(io_ins_left_1[58]),
    .Y(net630));
 BUFx2_ASAP7_75t_R input631 (.A(io_ins_left_1[59]),
    .Y(net631));
 BUFx2_ASAP7_75t_R input632 (.A(io_ins_left_1[5]),
    .Y(net632));
 BUFx2_ASAP7_75t_R input633 (.A(io_ins_left_1[60]),
    .Y(net633));
 BUFx2_ASAP7_75t_R input634 (.A(io_ins_left_1[61]),
    .Y(net634));
 BUFx2_ASAP7_75t_R input635 (.A(io_ins_left_1[62]),
    .Y(net635));
 BUFx2_ASAP7_75t_R input636 (.A(io_ins_left_1[63]),
    .Y(net636));
 BUFx2_ASAP7_75t_R input637 (.A(io_ins_left_1[6]),
    .Y(net637));
 BUFx2_ASAP7_75t_R input638 (.A(io_ins_left_1[7]),
    .Y(net638));
 BUFx2_ASAP7_75t_R input639 (.A(io_ins_left_1[8]),
    .Y(net639));
 BUFx2_ASAP7_75t_R input640 (.A(io_ins_left_1[9]),
    .Y(net640));
 BUFx2_ASAP7_75t_R input641 (.A(io_ins_left_2[0]),
    .Y(net641));
 BUFx2_ASAP7_75t_R input642 (.A(io_ins_left_2[10]),
    .Y(net642));
 BUFx2_ASAP7_75t_R input643 (.A(io_ins_left_2[11]),
    .Y(net643));
 BUFx2_ASAP7_75t_R input644 (.A(io_ins_left_2[12]),
    .Y(net644));
 BUFx2_ASAP7_75t_R input645 (.A(io_ins_left_2[13]),
    .Y(net645));
 BUFx2_ASAP7_75t_R input646 (.A(io_ins_left_2[14]),
    .Y(net646));
 BUFx2_ASAP7_75t_R input647 (.A(io_ins_left_2[15]),
    .Y(net647));
 BUFx2_ASAP7_75t_R input648 (.A(io_ins_left_2[16]),
    .Y(net648));
 BUFx2_ASAP7_75t_R input649 (.A(io_ins_left_2[17]),
    .Y(net649));
 BUFx2_ASAP7_75t_R input650 (.A(io_ins_left_2[18]),
    .Y(net650));
 BUFx2_ASAP7_75t_R input651 (.A(io_ins_left_2[19]),
    .Y(net651));
 BUFx2_ASAP7_75t_R input652 (.A(io_ins_left_2[1]),
    .Y(net652));
 BUFx2_ASAP7_75t_R input653 (.A(io_ins_left_2[20]),
    .Y(net653));
 BUFx2_ASAP7_75t_R input654 (.A(io_ins_left_2[21]),
    .Y(net654));
 BUFx2_ASAP7_75t_R input655 (.A(io_ins_left_2[22]),
    .Y(net655));
 BUFx2_ASAP7_75t_R input656 (.A(io_ins_left_2[23]),
    .Y(net656));
 BUFx2_ASAP7_75t_R input657 (.A(io_ins_left_2[24]),
    .Y(net657));
 BUFx2_ASAP7_75t_R input658 (.A(io_ins_left_2[25]),
    .Y(net658));
 BUFx2_ASAP7_75t_R input659 (.A(io_ins_left_2[26]),
    .Y(net659));
 BUFx2_ASAP7_75t_R input660 (.A(io_ins_left_2[27]),
    .Y(net660));
 BUFx2_ASAP7_75t_R input661 (.A(io_ins_left_2[28]),
    .Y(net661));
 BUFx2_ASAP7_75t_R input662 (.A(io_ins_left_2[29]),
    .Y(net662));
 BUFx2_ASAP7_75t_R input663 (.A(io_ins_left_2[2]),
    .Y(net663));
 BUFx2_ASAP7_75t_R input664 (.A(io_ins_left_2[30]),
    .Y(net664));
 BUFx2_ASAP7_75t_R input665 (.A(io_ins_left_2[31]),
    .Y(net665));
 BUFx2_ASAP7_75t_R input666 (.A(io_ins_left_2[32]),
    .Y(net666));
 BUFx2_ASAP7_75t_R input667 (.A(io_ins_left_2[33]),
    .Y(net667));
 BUFx2_ASAP7_75t_R input668 (.A(io_ins_left_2[34]),
    .Y(net668));
 BUFx2_ASAP7_75t_R input669 (.A(io_ins_left_2[35]),
    .Y(net669));
 BUFx2_ASAP7_75t_R input670 (.A(io_ins_left_2[36]),
    .Y(net670));
 BUFx2_ASAP7_75t_R input671 (.A(io_ins_left_2[37]),
    .Y(net671));
 BUFx2_ASAP7_75t_R input672 (.A(io_ins_left_2[38]),
    .Y(net672));
 BUFx2_ASAP7_75t_R input673 (.A(io_ins_left_2[39]),
    .Y(net673));
 BUFx2_ASAP7_75t_R input674 (.A(io_ins_left_2[3]),
    .Y(net674));
 BUFx2_ASAP7_75t_R input675 (.A(io_ins_left_2[40]),
    .Y(net675));
 BUFx2_ASAP7_75t_R input676 (.A(io_ins_left_2[41]),
    .Y(net676));
 BUFx2_ASAP7_75t_R input677 (.A(io_ins_left_2[42]),
    .Y(net677));
 BUFx2_ASAP7_75t_R input678 (.A(io_ins_left_2[43]),
    .Y(net678));
 BUFx2_ASAP7_75t_R input679 (.A(io_ins_left_2[44]),
    .Y(net679));
 BUFx2_ASAP7_75t_R input680 (.A(io_ins_left_2[45]),
    .Y(net680));
 BUFx2_ASAP7_75t_R input681 (.A(io_ins_left_2[46]),
    .Y(net681));
 BUFx2_ASAP7_75t_R input682 (.A(io_ins_left_2[47]),
    .Y(net682));
 BUFx2_ASAP7_75t_R input683 (.A(io_ins_left_2[48]),
    .Y(net683));
 BUFx2_ASAP7_75t_R input684 (.A(io_ins_left_2[49]),
    .Y(net684));
 BUFx2_ASAP7_75t_R input685 (.A(io_ins_left_2[4]),
    .Y(net685));
 BUFx2_ASAP7_75t_R input686 (.A(io_ins_left_2[50]),
    .Y(net686));
 BUFx2_ASAP7_75t_R input687 (.A(io_ins_left_2[51]),
    .Y(net687));
 BUFx2_ASAP7_75t_R input688 (.A(io_ins_left_2[52]),
    .Y(net688));
 BUFx2_ASAP7_75t_R input689 (.A(io_ins_left_2[53]),
    .Y(net689));
 BUFx2_ASAP7_75t_R input690 (.A(io_ins_left_2[54]),
    .Y(net690));
 BUFx2_ASAP7_75t_R input691 (.A(io_ins_left_2[55]),
    .Y(net691));
 BUFx2_ASAP7_75t_R input692 (.A(io_ins_left_2[56]),
    .Y(net692));
 BUFx2_ASAP7_75t_R input693 (.A(io_ins_left_2[57]),
    .Y(net693));
 BUFx2_ASAP7_75t_R input694 (.A(io_ins_left_2[58]),
    .Y(net694));
 BUFx2_ASAP7_75t_R input695 (.A(io_ins_left_2[59]),
    .Y(net695));
 BUFx2_ASAP7_75t_R input696 (.A(io_ins_left_2[5]),
    .Y(net696));
 BUFx2_ASAP7_75t_R input697 (.A(io_ins_left_2[60]),
    .Y(net697));
 BUFx2_ASAP7_75t_R input698 (.A(io_ins_left_2[61]),
    .Y(net698));
 BUFx2_ASAP7_75t_R input699 (.A(io_ins_left_2[62]),
    .Y(net699));
 BUFx2_ASAP7_75t_R input700 (.A(io_ins_left_2[63]),
    .Y(net700));
 BUFx2_ASAP7_75t_R input701 (.A(io_ins_left_2[6]),
    .Y(net701));
 BUFx2_ASAP7_75t_R input702 (.A(io_ins_left_2[7]),
    .Y(net702));
 BUFx2_ASAP7_75t_R input703 (.A(io_ins_left_2[8]),
    .Y(net703));
 BUFx2_ASAP7_75t_R input704 (.A(io_ins_left_2[9]),
    .Y(net704));
 BUFx2_ASAP7_75t_R input705 (.A(io_ins_left_3[0]),
    .Y(net705));
 BUFx2_ASAP7_75t_R input706 (.A(io_ins_left_3[10]),
    .Y(net706));
 BUFx2_ASAP7_75t_R input707 (.A(io_ins_left_3[11]),
    .Y(net707));
 BUFx2_ASAP7_75t_R input708 (.A(io_ins_left_3[12]),
    .Y(net708));
 BUFx2_ASAP7_75t_R input709 (.A(io_ins_left_3[13]),
    .Y(net709));
 BUFx2_ASAP7_75t_R input710 (.A(io_ins_left_3[14]),
    .Y(net710));
 BUFx2_ASAP7_75t_R input711 (.A(io_ins_left_3[15]),
    .Y(net711));
 BUFx2_ASAP7_75t_R input712 (.A(io_ins_left_3[16]),
    .Y(net712));
 BUFx2_ASAP7_75t_R input713 (.A(io_ins_left_3[17]),
    .Y(net713));
 BUFx2_ASAP7_75t_R input714 (.A(io_ins_left_3[18]),
    .Y(net714));
 BUFx2_ASAP7_75t_R input715 (.A(io_ins_left_3[19]),
    .Y(net715));
 BUFx2_ASAP7_75t_R input716 (.A(io_ins_left_3[1]),
    .Y(net716));
 BUFx2_ASAP7_75t_R input717 (.A(io_ins_left_3[20]),
    .Y(net717));
 BUFx2_ASAP7_75t_R input718 (.A(io_ins_left_3[21]),
    .Y(net718));
 BUFx2_ASAP7_75t_R input719 (.A(io_ins_left_3[22]),
    .Y(net719));
 BUFx2_ASAP7_75t_R input720 (.A(io_ins_left_3[23]),
    .Y(net720));
 BUFx2_ASAP7_75t_R input721 (.A(io_ins_left_3[24]),
    .Y(net721));
 BUFx2_ASAP7_75t_R input722 (.A(io_ins_left_3[25]),
    .Y(net722));
 BUFx2_ASAP7_75t_R input723 (.A(io_ins_left_3[26]),
    .Y(net723));
 BUFx2_ASAP7_75t_R input724 (.A(io_ins_left_3[27]),
    .Y(net724));
 BUFx2_ASAP7_75t_R input725 (.A(io_ins_left_3[28]),
    .Y(net725));
 BUFx2_ASAP7_75t_R input726 (.A(io_ins_left_3[29]),
    .Y(net726));
 BUFx2_ASAP7_75t_R input727 (.A(io_ins_left_3[2]),
    .Y(net727));
 BUFx2_ASAP7_75t_R input728 (.A(io_ins_left_3[30]),
    .Y(net728));
 BUFx2_ASAP7_75t_R input729 (.A(io_ins_left_3[31]),
    .Y(net729));
 BUFx2_ASAP7_75t_R input730 (.A(io_ins_left_3[32]),
    .Y(net730));
 BUFx2_ASAP7_75t_R input731 (.A(io_ins_left_3[33]),
    .Y(net731));
 BUFx2_ASAP7_75t_R input732 (.A(io_ins_left_3[34]),
    .Y(net732));
 BUFx2_ASAP7_75t_R input733 (.A(io_ins_left_3[35]),
    .Y(net733));
 BUFx2_ASAP7_75t_R input734 (.A(io_ins_left_3[36]),
    .Y(net734));
 BUFx2_ASAP7_75t_R input735 (.A(io_ins_left_3[37]),
    .Y(net735));
 BUFx2_ASAP7_75t_R input736 (.A(io_ins_left_3[38]),
    .Y(net736));
 BUFx2_ASAP7_75t_R input737 (.A(io_ins_left_3[39]),
    .Y(net737));
 BUFx2_ASAP7_75t_R input738 (.A(io_ins_left_3[3]),
    .Y(net738));
 BUFx2_ASAP7_75t_R input739 (.A(io_ins_left_3[40]),
    .Y(net739));
 BUFx2_ASAP7_75t_R input740 (.A(io_ins_left_3[41]),
    .Y(net740));
 BUFx2_ASAP7_75t_R input741 (.A(io_ins_left_3[42]),
    .Y(net741));
 BUFx2_ASAP7_75t_R input742 (.A(io_ins_left_3[43]),
    .Y(net742));
 BUFx2_ASAP7_75t_R input743 (.A(io_ins_left_3[44]),
    .Y(net743));
 BUFx2_ASAP7_75t_R input744 (.A(io_ins_left_3[45]),
    .Y(net744));
 BUFx2_ASAP7_75t_R input745 (.A(io_ins_left_3[46]),
    .Y(net745));
 BUFx2_ASAP7_75t_R input746 (.A(io_ins_left_3[47]),
    .Y(net746));
 BUFx2_ASAP7_75t_R input747 (.A(io_ins_left_3[48]),
    .Y(net747));
 BUFx2_ASAP7_75t_R input748 (.A(io_ins_left_3[49]),
    .Y(net748));
 BUFx2_ASAP7_75t_R input749 (.A(io_ins_left_3[4]),
    .Y(net749));
 BUFx2_ASAP7_75t_R input750 (.A(io_ins_left_3[50]),
    .Y(net750));
 BUFx2_ASAP7_75t_R input751 (.A(io_ins_left_3[51]),
    .Y(net751));
 BUFx2_ASAP7_75t_R input752 (.A(io_ins_left_3[52]),
    .Y(net752));
 BUFx2_ASAP7_75t_R input753 (.A(io_ins_left_3[53]),
    .Y(net753));
 BUFx2_ASAP7_75t_R input754 (.A(io_ins_left_3[54]),
    .Y(net754));
 BUFx2_ASAP7_75t_R input755 (.A(io_ins_left_3[55]),
    .Y(net755));
 BUFx2_ASAP7_75t_R input756 (.A(io_ins_left_3[56]),
    .Y(net756));
 BUFx2_ASAP7_75t_R input757 (.A(io_ins_left_3[57]),
    .Y(net757));
 BUFx2_ASAP7_75t_R input758 (.A(io_ins_left_3[58]),
    .Y(net758));
 BUFx2_ASAP7_75t_R input759 (.A(io_ins_left_3[59]),
    .Y(net759));
 BUFx2_ASAP7_75t_R input760 (.A(io_ins_left_3[5]),
    .Y(net760));
 BUFx2_ASAP7_75t_R input761 (.A(io_ins_left_3[60]),
    .Y(net761));
 BUFx2_ASAP7_75t_R input762 (.A(io_ins_left_3[61]),
    .Y(net762));
 BUFx2_ASAP7_75t_R input763 (.A(io_ins_left_3[62]),
    .Y(net763));
 BUFx2_ASAP7_75t_R input764 (.A(io_ins_left_3[63]),
    .Y(net764));
 BUFx2_ASAP7_75t_R input765 (.A(io_ins_left_3[6]),
    .Y(net765));
 BUFx2_ASAP7_75t_R input766 (.A(io_ins_left_3[7]),
    .Y(net766));
 BUFx2_ASAP7_75t_R input767 (.A(io_ins_left_3[8]),
    .Y(net767));
 BUFx2_ASAP7_75t_R input768 (.A(io_ins_left_3[9]),
    .Y(net768));
 BUFx2_ASAP7_75t_R input769 (.A(io_ins_left_4[0]),
    .Y(net769));
 BUFx2_ASAP7_75t_R input770 (.A(io_ins_left_4[10]),
    .Y(net770));
 BUFx2_ASAP7_75t_R input771 (.A(io_ins_left_4[11]),
    .Y(net771));
 BUFx2_ASAP7_75t_R input772 (.A(io_ins_left_4[12]),
    .Y(net772));
 BUFx2_ASAP7_75t_R input773 (.A(io_ins_left_4[13]),
    .Y(net773));
 BUFx2_ASAP7_75t_R input774 (.A(io_ins_left_4[14]),
    .Y(net774));
 BUFx2_ASAP7_75t_R input775 (.A(io_ins_left_4[15]),
    .Y(net775));
 BUFx2_ASAP7_75t_R input776 (.A(io_ins_left_4[16]),
    .Y(net776));
 BUFx2_ASAP7_75t_R input777 (.A(io_ins_left_4[17]),
    .Y(net777));
 BUFx2_ASAP7_75t_R input778 (.A(io_ins_left_4[18]),
    .Y(net778));
 BUFx2_ASAP7_75t_R input779 (.A(io_ins_left_4[19]),
    .Y(net779));
 BUFx2_ASAP7_75t_R input780 (.A(io_ins_left_4[1]),
    .Y(net780));
 BUFx2_ASAP7_75t_R input781 (.A(io_ins_left_4[20]),
    .Y(net781));
 BUFx2_ASAP7_75t_R input782 (.A(io_ins_left_4[21]),
    .Y(net782));
 BUFx2_ASAP7_75t_R input783 (.A(io_ins_left_4[22]),
    .Y(net783));
 BUFx2_ASAP7_75t_R input784 (.A(io_ins_left_4[23]),
    .Y(net784));
 BUFx2_ASAP7_75t_R input785 (.A(io_ins_left_4[24]),
    .Y(net785));
 BUFx2_ASAP7_75t_R input786 (.A(io_ins_left_4[25]),
    .Y(net786));
 BUFx2_ASAP7_75t_R input787 (.A(io_ins_left_4[26]),
    .Y(net787));
 BUFx2_ASAP7_75t_R input788 (.A(io_ins_left_4[27]),
    .Y(net788));
 BUFx2_ASAP7_75t_R input789 (.A(io_ins_left_4[28]),
    .Y(net789));
 BUFx2_ASAP7_75t_R input790 (.A(io_ins_left_4[29]),
    .Y(net790));
 BUFx2_ASAP7_75t_R input791 (.A(io_ins_left_4[2]),
    .Y(net791));
 BUFx2_ASAP7_75t_R input792 (.A(io_ins_left_4[30]),
    .Y(net792));
 BUFx2_ASAP7_75t_R input793 (.A(io_ins_left_4[31]),
    .Y(net793));
 BUFx2_ASAP7_75t_R input794 (.A(io_ins_left_4[32]),
    .Y(net794));
 BUFx2_ASAP7_75t_R input795 (.A(io_ins_left_4[33]),
    .Y(net795));
 BUFx2_ASAP7_75t_R input796 (.A(io_ins_left_4[34]),
    .Y(net796));
 BUFx2_ASAP7_75t_R input797 (.A(io_ins_left_4[35]),
    .Y(net797));
 BUFx2_ASAP7_75t_R input798 (.A(io_ins_left_4[36]),
    .Y(net798));
 BUFx2_ASAP7_75t_R input799 (.A(io_ins_left_4[37]),
    .Y(net799));
 BUFx2_ASAP7_75t_R input800 (.A(io_ins_left_4[38]),
    .Y(net800));
 BUFx2_ASAP7_75t_R input801 (.A(io_ins_left_4[39]),
    .Y(net801));
 BUFx2_ASAP7_75t_R input802 (.A(io_ins_left_4[3]),
    .Y(net802));
 BUFx2_ASAP7_75t_R input803 (.A(io_ins_left_4[40]),
    .Y(net803));
 BUFx2_ASAP7_75t_R input804 (.A(io_ins_left_4[41]),
    .Y(net804));
 BUFx2_ASAP7_75t_R input805 (.A(io_ins_left_4[42]),
    .Y(net805));
 BUFx2_ASAP7_75t_R input806 (.A(io_ins_left_4[43]),
    .Y(net806));
 BUFx2_ASAP7_75t_R input807 (.A(io_ins_left_4[44]),
    .Y(net807));
 BUFx2_ASAP7_75t_R input808 (.A(io_ins_left_4[45]),
    .Y(net808));
 BUFx2_ASAP7_75t_R input809 (.A(io_ins_left_4[46]),
    .Y(net809));
 BUFx2_ASAP7_75t_R input810 (.A(io_ins_left_4[47]),
    .Y(net810));
 BUFx2_ASAP7_75t_R input811 (.A(io_ins_left_4[48]),
    .Y(net811));
 BUFx2_ASAP7_75t_R input812 (.A(io_ins_left_4[49]),
    .Y(net812));
 BUFx2_ASAP7_75t_R input813 (.A(io_ins_left_4[4]),
    .Y(net813));
 BUFx2_ASAP7_75t_R input814 (.A(io_ins_left_4[50]),
    .Y(net814));
 BUFx2_ASAP7_75t_R input815 (.A(io_ins_left_4[51]),
    .Y(net815));
 BUFx2_ASAP7_75t_R input816 (.A(io_ins_left_4[52]),
    .Y(net816));
 BUFx2_ASAP7_75t_R input817 (.A(io_ins_left_4[53]),
    .Y(net817));
 BUFx2_ASAP7_75t_R input818 (.A(io_ins_left_4[54]),
    .Y(net818));
 BUFx2_ASAP7_75t_R input819 (.A(io_ins_left_4[55]),
    .Y(net819));
 BUFx2_ASAP7_75t_R input820 (.A(io_ins_left_4[56]),
    .Y(net820));
 BUFx2_ASAP7_75t_R input821 (.A(io_ins_left_4[57]),
    .Y(net821));
 BUFx2_ASAP7_75t_R input822 (.A(io_ins_left_4[58]),
    .Y(net822));
 BUFx2_ASAP7_75t_R input823 (.A(io_ins_left_4[59]),
    .Y(net823));
 BUFx2_ASAP7_75t_R input824 (.A(io_ins_left_4[5]),
    .Y(net824));
 BUFx2_ASAP7_75t_R input825 (.A(io_ins_left_4[60]),
    .Y(net825));
 BUFx2_ASAP7_75t_R input826 (.A(io_ins_left_4[61]),
    .Y(net826));
 BUFx2_ASAP7_75t_R input827 (.A(io_ins_left_4[62]),
    .Y(net827));
 BUFx2_ASAP7_75t_R input828 (.A(io_ins_left_4[63]),
    .Y(net828));
 BUFx2_ASAP7_75t_R input829 (.A(io_ins_left_4[6]),
    .Y(net829));
 BUFx2_ASAP7_75t_R input830 (.A(io_ins_left_4[7]),
    .Y(net830));
 BUFx2_ASAP7_75t_R input831 (.A(io_ins_left_4[8]),
    .Y(net831));
 BUFx2_ASAP7_75t_R input832 (.A(io_ins_left_4[9]),
    .Y(net832));
 BUFx2_ASAP7_75t_R input833 (.A(io_ins_left_5[0]),
    .Y(net833));
 BUFx2_ASAP7_75t_R input834 (.A(io_ins_left_5[10]),
    .Y(net834));
 BUFx2_ASAP7_75t_R input835 (.A(io_ins_left_5[11]),
    .Y(net835));
 BUFx2_ASAP7_75t_R input836 (.A(io_ins_left_5[12]),
    .Y(net836));
 BUFx2_ASAP7_75t_R input837 (.A(io_ins_left_5[13]),
    .Y(net837));
 BUFx2_ASAP7_75t_R input838 (.A(io_ins_left_5[14]),
    .Y(net838));
 BUFx2_ASAP7_75t_R input839 (.A(io_ins_left_5[15]),
    .Y(net839));
 BUFx2_ASAP7_75t_R input840 (.A(io_ins_left_5[16]),
    .Y(net840));
 BUFx2_ASAP7_75t_R input841 (.A(io_ins_left_5[17]),
    .Y(net841));
 BUFx2_ASAP7_75t_R input842 (.A(io_ins_left_5[18]),
    .Y(net842));
 BUFx2_ASAP7_75t_R input843 (.A(io_ins_left_5[19]),
    .Y(net843));
 BUFx2_ASAP7_75t_R input844 (.A(io_ins_left_5[1]),
    .Y(net844));
 BUFx2_ASAP7_75t_R input845 (.A(io_ins_left_5[20]),
    .Y(net845));
 BUFx2_ASAP7_75t_R input846 (.A(io_ins_left_5[21]),
    .Y(net846));
 BUFx2_ASAP7_75t_R input847 (.A(io_ins_left_5[22]),
    .Y(net847));
 BUFx2_ASAP7_75t_R input848 (.A(io_ins_left_5[23]),
    .Y(net848));
 BUFx2_ASAP7_75t_R input849 (.A(io_ins_left_5[24]),
    .Y(net849));
 BUFx2_ASAP7_75t_R input850 (.A(io_ins_left_5[25]),
    .Y(net850));
 BUFx2_ASAP7_75t_R input851 (.A(io_ins_left_5[26]),
    .Y(net851));
 BUFx2_ASAP7_75t_R input852 (.A(io_ins_left_5[27]),
    .Y(net852));
 BUFx2_ASAP7_75t_R input853 (.A(io_ins_left_5[28]),
    .Y(net853));
 BUFx2_ASAP7_75t_R input854 (.A(io_ins_left_5[29]),
    .Y(net854));
 BUFx2_ASAP7_75t_R input855 (.A(io_ins_left_5[2]),
    .Y(net855));
 BUFx2_ASAP7_75t_R input856 (.A(io_ins_left_5[30]),
    .Y(net856));
 BUFx2_ASAP7_75t_R input857 (.A(io_ins_left_5[31]),
    .Y(net857));
 BUFx2_ASAP7_75t_R input858 (.A(io_ins_left_5[32]),
    .Y(net858));
 BUFx2_ASAP7_75t_R input859 (.A(io_ins_left_5[33]),
    .Y(net859));
 BUFx2_ASAP7_75t_R input860 (.A(io_ins_left_5[34]),
    .Y(net860));
 BUFx2_ASAP7_75t_R input861 (.A(io_ins_left_5[35]),
    .Y(net861));
 BUFx2_ASAP7_75t_R input862 (.A(io_ins_left_5[36]),
    .Y(net862));
 BUFx2_ASAP7_75t_R input863 (.A(io_ins_left_5[37]),
    .Y(net863));
 BUFx2_ASAP7_75t_R input864 (.A(io_ins_left_5[38]),
    .Y(net864));
 BUFx2_ASAP7_75t_R input865 (.A(io_ins_left_5[39]),
    .Y(net865));
 BUFx2_ASAP7_75t_R input866 (.A(io_ins_left_5[3]),
    .Y(net866));
 BUFx2_ASAP7_75t_R input867 (.A(io_ins_left_5[40]),
    .Y(net867));
 BUFx2_ASAP7_75t_R input868 (.A(io_ins_left_5[41]),
    .Y(net868));
 BUFx2_ASAP7_75t_R input869 (.A(io_ins_left_5[42]),
    .Y(net869));
 BUFx2_ASAP7_75t_R input870 (.A(io_ins_left_5[43]),
    .Y(net870));
 BUFx2_ASAP7_75t_R input871 (.A(io_ins_left_5[44]),
    .Y(net871));
 BUFx2_ASAP7_75t_R input872 (.A(io_ins_left_5[45]),
    .Y(net872));
 BUFx2_ASAP7_75t_R input873 (.A(io_ins_left_5[46]),
    .Y(net873));
 BUFx2_ASAP7_75t_R input874 (.A(io_ins_left_5[47]),
    .Y(net874));
 BUFx2_ASAP7_75t_R input875 (.A(io_ins_left_5[48]),
    .Y(net875));
 BUFx2_ASAP7_75t_R input876 (.A(io_ins_left_5[49]),
    .Y(net876));
 BUFx2_ASAP7_75t_R input877 (.A(io_ins_left_5[4]),
    .Y(net877));
 BUFx2_ASAP7_75t_R input878 (.A(io_ins_left_5[50]),
    .Y(net878));
 BUFx2_ASAP7_75t_R input879 (.A(io_ins_left_5[51]),
    .Y(net879));
 BUFx2_ASAP7_75t_R input880 (.A(io_ins_left_5[52]),
    .Y(net880));
 BUFx2_ASAP7_75t_R input881 (.A(io_ins_left_5[53]),
    .Y(net881));
 BUFx2_ASAP7_75t_R input882 (.A(io_ins_left_5[54]),
    .Y(net882));
 BUFx2_ASAP7_75t_R input883 (.A(io_ins_left_5[55]),
    .Y(net883));
 BUFx2_ASAP7_75t_R input884 (.A(io_ins_left_5[56]),
    .Y(net884));
 BUFx2_ASAP7_75t_R input885 (.A(io_ins_left_5[57]),
    .Y(net885));
 BUFx2_ASAP7_75t_R input886 (.A(io_ins_left_5[58]),
    .Y(net886));
 BUFx2_ASAP7_75t_R input887 (.A(io_ins_left_5[59]),
    .Y(net887));
 BUFx2_ASAP7_75t_R input888 (.A(io_ins_left_5[5]),
    .Y(net888));
 BUFx2_ASAP7_75t_R input889 (.A(io_ins_left_5[60]),
    .Y(net889));
 BUFx2_ASAP7_75t_R input890 (.A(io_ins_left_5[61]),
    .Y(net890));
 BUFx2_ASAP7_75t_R input891 (.A(io_ins_left_5[62]),
    .Y(net891));
 BUFx2_ASAP7_75t_R input892 (.A(io_ins_left_5[63]),
    .Y(net892));
 BUFx2_ASAP7_75t_R input893 (.A(io_ins_left_5[6]),
    .Y(net893));
 BUFx2_ASAP7_75t_R input894 (.A(io_ins_left_5[7]),
    .Y(net894));
 BUFx2_ASAP7_75t_R input895 (.A(io_ins_left_5[8]),
    .Y(net895));
 BUFx2_ASAP7_75t_R input896 (.A(io_ins_left_5[9]),
    .Y(net896));
 BUFx2_ASAP7_75t_R input897 (.A(io_ins_left_6[0]),
    .Y(net897));
 BUFx2_ASAP7_75t_R input898 (.A(io_ins_left_6[10]),
    .Y(net898));
 BUFx2_ASAP7_75t_R input899 (.A(io_ins_left_6[11]),
    .Y(net899));
 BUFx2_ASAP7_75t_R input900 (.A(io_ins_left_6[12]),
    .Y(net900));
 BUFx2_ASAP7_75t_R input901 (.A(io_ins_left_6[13]),
    .Y(net901));
 BUFx2_ASAP7_75t_R input902 (.A(io_ins_left_6[14]),
    .Y(net902));
 BUFx2_ASAP7_75t_R input903 (.A(io_ins_left_6[15]),
    .Y(net903));
 BUFx2_ASAP7_75t_R input904 (.A(io_ins_left_6[16]),
    .Y(net904));
 BUFx2_ASAP7_75t_R input905 (.A(io_ins_left_6[17]),
    .Y(net905));
 BUFx2_ASAP7_75t_R input906 (.A(io_ins_left_6[18]),
    .Y(net906));
 BUFx2_ASAP7_75t_R input907 (.A(io_ins_left_6[19]),
    .Y(net907));
 BUFx2_ASAP7_75t_R input908 (.A(io_ins_left_6[1]),
    .Y(net908));
 BUFx2_ASAP7_75t_R input909 (.A(io_ins_left_6[20]),
    .Y(net909));
 BUFx2_ASAP7_75t_R input910 (.A(io_ins_left_6[21]),
    .Y(net910));
 BUFx2_ASAP7_75t_R input911 (.A(io_ins_left_6[22]),
    .Y(net911));
 BUFx2_ASAP7_75t_R input912 (.A(io_ins_left_6[23]),
    .Y(net912));
 BUFx2_ASAP7_75t_R input913 (.A(io_ins_left_6[24]),
    .Y(net913));
 BUFx2_ASAP7_75t_R input914 (.A(io_ins_left_6[25]),
    .Y(net914));
 BUFx2_ASAP7_75t_R input915 (.A(io_ins_left_6[26]),
    .Y(net915));
 BUFx2_ASAP7_75t_R input916 (.A(io_ins_left_6[27]),
    .Y(net916));
 BUFx2_ASAP7_75t_R input917 (.A(io_ins_left_6[28]),
    .Y(net917));
 BUFx2_ASAP7_75t_R input918 (.A(io_ins_left_6[29]),
    .Y(net918));
 BUFx2_ASAP7_75t_R input919 (.A(io_ins_left_6[2]),
    .Y(net919));
 BUFx2_ASAP7_75t_R input920 (.A(io_ins_left_6[30]),
    .Y(net920));
 BUFx2_ASAP7_75t_R input921 (.A(io_ins_left_6[31]),
    .Y(net921));
 BUFx2_ASAP7_75t_R input922 (.A(io_ins_left_6[32]),
    .Y(net922));
 BUFx2_ASAP7_75t_R input923 (.A(io_ins_left_6[33]),
    .Y(net923));
 BUFx2_ASAP7_75t_R input924 (.A(io_ins_left_6[34]),
    .Y(net924));
 BUFx2_ASAP7_75t_R input925 (.A(io_ins_left_6[35]),
    .Y(net925));
 BUFx2_ASAP7_75t_R input926 (.A(io_ins_left_6[36]),
    .Y(net926));
 BUFx2_ASAP7_75t_R input927 (.A(io_ins_left_6[37]),
    .Y(net927));
 BUFx2_ASAP7_75t_R input928 (.A(io_ins_left_6[38]),
    .Y(net928));
 BUFx2_ASAP7_75t_R input929 (.A(io_ins_left_6[39]),
    .Y(net929));
 BUFx2_ASAP7_75t_R input930 (.A(io_ins_left_6[3]),
    .Y(net930));
 BUFx2_ASAP7_75t_R input931 (.A(io_ins_left_6[40]),
    .Y(net931));
 BUFx2_ASAP7_75t_R input932 (.A(io_ins_left_6[41]),
    .Y(net932));
 BUFx2_ASAP7_75t_R input933 (.A(io_ins_left_6[42]),
    .Y(net933));
 BUFx2_ASAP7_75t_R input934 (.A(io_ins_left_6[43]),
    .Y(net934));
 BUFx2_ASAP7_75t_R input935 (.A(io_ins_left_6[44]),
    .Y(net935));
 BUFx2_ASAP7_75t_R input936 (.A(io_ins_left_6[45]),
    .Y(net936));
 BUFx2_ASAP7_75t_R input937 (.A(io_ins_left_6[46]),
    .Y(net937));
 BUFx2_ASAP7_75t_R input938 (.A(io_ins_left_6[47]),
    .Y(net938));
 BUFx2_ASAP7_75t_R input939 (.A(io_ins_left_6[48]),
    .Y(net939));
 BUFx2_ASAP7_75t_R input940 (.A(io_ins_left_6[49]),
    .Y(net940));
 BUFx2_ASAP7_75t_R input941 (.A(io_ins_left_6[4]),
    .Y(net941));
 BUFx2_ASAP7_75t_R input942 (.A(io_ins_left_6[50]),
    .Y(net942));
 BUFx2_ASAP7_75t_R input943 (.A(io_ins_left_6[51]),
    .Y(net943));
 BUFx2_ASAP7_75t_R input944 (.A(io_ins_left_6[52]),
    .Y(net944));
 BUFx2_ASAP7_75t_R input945 (.A(io_ins_left_6[53]),
    .Y(net945));
 BUFx2_ASAP7_75t_R input946 (.A(io_ins_left_6[54]),
    .Y(net946));
 BUFx2_ASAP7_75t_R input947 (.A(io_ins_left_6[55]),
    .Y(net947));
 BUFx2_ASAP7_75t_R input948 (.A(io_ins_left_6[56]),
    .Y(net948));
 BUFx2_ASAP7_75t_R input949 (.A(io_ins_left_6[57]),
    .Y(net949));
 BUFx2_ASAP7_75t_R input950 (.A(io_ins_left_6[58]),
    .Y(net950));
 BUFx2_ASAP7_75t_R input951 (.A(io_ins_left_6[59]),
    .Y(net951));
 BUFx2_ASAP7_75t_R input952 (.A(io_ins_left_6[5]),
    .Y(net952));
 BUFx2_ASAP7_75t_R input953 (.A(io_ins_left_6[60]),
    .Y(net953));
 BUFx2_ASAP7_75t_R input954 (.A(io_ins_left_6[61]),
    .Y(net954));
 BUFx2_ASAP7_75t_R input955 (.A(io_ins_left_6[62]),
    .Y(net955));
 BUFx2_ASAP7_75t_R input956 (.A(io_ins_left_6[63]),
    .Y(net956));
 BUFx2_ASAP7_75t_R input957 (.A(io_ins_left_6[6]),
    .Y(net957));
 BUFx2_ASAP7_75t_R input958 (.A(io_ins_left_6[7]),
    .Y(net958));
 BUFx2_ASAP7_75t_R input959 (.A(io_ins_left_6[8]),
    .Y(net959));
 BUFx2_ASAP7_75t_R input960 (.A(io_ins_left_6[9]),
    .Y(net960));
 BUFx2_ASAP7_75t_R input961 (.A(io_ins_left_7[0]),
    .Y(net961));
 BUFx2_ASAP7_75t_R input962 (.A(io_ins_left_7[10]),
    .Y(net962));
 BUFx2_ASAP7_75t_R input963 (.A(io_ins_left_7[11]),
    .Y(net963));
 BUFx2_ASAP7_75t_R input964 (.A(io_ins_left_7[12]),
    .Y(net964));
 BUFx2_ASAP7_75t_R input965 (.A(io_ins_left_7[13]),
    .Y(net965));
 BUFx2_ASAP7_75t_R input966 (.A(io_ins_left_7[14]),
    .Y(net966));
 BUFx2_ASAP7_75t_R input967 (.A(io_ins_left_7[15]),
    .Y(net967));
 BUFx2_ASAP7_75t_R input968 (.A(io_ins_left_7[16]),
    .Y(net968));
 BUFx2_ASAP7_75t_R input969 (.A(io_ins_left_7[17]),
    .Y(net969));
 BUFx2_ASAP7_75t_R input970 (.A(io_ins_left_7[18]),
    .Y(net970));
 BUFx2_ASAP7_75t_R input971 (.A(io_ins_left_7[19]),
    .Y(net971));
 BUFx2_ASAP7_75t_R input972 (.A(io_ins_left_7[1]),
    .Y(net972));
 BUFx2_ASAP7_75t_R input973 (.A(io_ins_left_7[20]),
    .Y(net973));
 BUFx2_ASAP7_75t_R input974 (.A(io_ins_left_7[21]),
    .Y(net974));
 BUFx2_ASAP7_75t_R input975 (.A(io_ins_left_7[22]),
    .Y(net975));
 BUFx2_ASAP7_75t_R input976 (.A(io_ins_left_7[23]),
    .Y(net976));
 BUFx2_ASAP7_75t_R input977 (.A(io_ins_left_7[24]),
    .Y(net977));
 BUFx2_ASAP7_75t_R input978 (.A(io_ins_left_7[25]),
    .Y(net978));
 BUFx2_ASAP7_75t_R input979 (.A(io_ins_left_7[26]),
    .Y(net979));
 BUFx2_ASAP7_75t_R input980 (.A(io_ins_left_7[27]),
    .Y(net980));
 BUFx2_ASAP7_75t_R input981 (.A(io_ins_left_7[28]),
    .Y(net981));
 BUFx2_ASAP7_75t_R input982 (.A(io_ins_left_7[29]),
    .Y(net982));
 BUFx2_ASAP7_75t_R input983 (.A(io_ins_left_7[2]),
    .Y(net983));
 BUFx2_ASAP7_75t_R input984 (.A(io_ins_left_7[30]),
    .Y(net984));
 BUFx2_ASAP7_75t_R input985 (.A(io_ins_left_7[31]),
    .Y(net985));
 BUFx2_ASAP7_75t_R input986 (.A(io_ins_left_7[32]),
    .Y(net986));
 BUFx2_ASAP7_75t_R input987 (.A(io_ins_left_7[33]),
    .Y(net987));
 BUFx2_ASAP7_75t_R input988 (.A(io_ins_left_7[34]),
    .Y(net988));
 BUFx2_ASAP7_75t_R input989 (.A(io_ins_left_7[35]),
    .Y(net989));
 BUFx2_ASAP7_75t_R input990 (.A(io_ins_left_7[36]),
    .Y(net990));
 BUFx2_ASAP7_75t_R input991 (.A(io_ins_left_7[37]),
    .Y(net991));
 BUFx2_ASAP7_75t_R input992 (.A(io_ins_left_7[38]),
    .Y(net992));
 BUFx2_ASAP7_75t_R input993 (.A(io_ins_left_7[39]),
    .Y(net993));
 BUFx2_ASAP7_75t_R input994 (.A(io_ins_left_7[3]),
    .Y(net994));
 BUFx2_ASAP7_75t_R input995 (.A(io_ins_left_7[40]),
    .Y(net995));
 BUFx2_ASAP7_75t_R input996 (.A(io_ins_left_7[41]),
    .Y(net996));
 BUFx2_ASAP7_75t_R input997 (.A(io_ins_left_7[42]),
    .Y(net997));
 BUFx2_ASAP7_75t_R input998 (.A(io_ins_left_7[43]),
    .Y(net998));
 BUFx2_ASAP7_75t_R input999 (.A(io_ins_left_7[44]),
    .Y(net999));
 BUFx2_ASAP7_75t_R input1000 (.A(io_ins_left_7[45]),
    .Y(net1000));
 BUFx2_ASAP7_75t_R input1001 (.A(io_ins_left_7[46]),
    .Y(net1001));
 BUFx2_ASAP7_75t_R input1002 (.A(io_ins_left_7[47]),
    .Y(net1002));
 BUFx2_ASAP7_75t_R input1003 (.A(io_ins_left_7[48]),
    .Y(net1003));
 BUFx2_ASAP7_75t_R input1004 (.A(io_ins_left_7[49]),
    .Y(net1004));
 BUFx2_ASAP7_75t_R input1005 (.A(io_ins_left_7[4]),
    .Y(net1005));
 BUFx2_ASAP7_75t_R input1006 (.A(io_ins_left_7[50]),
    .Y(net1006));
 BUFx2_ASAP7_75t_R input1007 (.A(io_ins_left_7[51]),
    .Y(net1007));
 BUFx2_ASAP7_75t_R input1008 (.A(io_ins_left_7[52]),
    .Y(net1008));
 BUFx2_ASAP7_75t_R input1009 (.A(io_ins_left_7[53]),
    .Y(net1009));
 BUFx2_ASAP7_75t_R input1010 (.A(io_ins_left_7[54]),
    .Y(net1010));
 BUFx2_ASAP7_75t_R input1011 (.A(io_ins_left_7[55]),
    .Y(net1011));
 BUFx2_ASAP7_75t_R input1012 (.A(io_ins_left_7[56]),
    .Y(net1012));
 BUFx2_ASAP7_75t_R input1013 (.A(io_ins_left_7[57]),
    .Y(net1013));
 BUFx2_ASAP7_75t_R input1014 (.A(io_ins_left_7[58]),
    .Y(net1014));
 BUFx2_ASAP7_75t_R input1015 (.A(io_ins_left_7[59]),
    .Y(net1015));
 BUFx2_ASAP7_75t_R input1016 (.A(io_ins_left_7[5]),
    .Y(net1016));
 BUFx2_ASAP7_75t_R input1017 (.A(io_ins_left_7[60]),
    .Y(net1017));
 BUFx2_ASAP7_75t_R input1018 (.A(io_ins_left_7[61]),
    .Y(net1018));
 BUFx2_ASAP7_75t_R input1019 (.A(io_ins_left_7[62]),
    .Y(net1019));
 BUFx2_ASAP7_75t_R input1020 (.A(io_ins_left_7[63]),
    .Y(net1020));
 BUFx2_ASAP7_75t_R input1021 (.A(io_ins_left_7[6]),
    .Y(net1021));
 BUFx2_ASAP7_75t_R input1022 (.A(io_ins_left_7[7]),
    .Y(net1022));
 BUFx2_ASAP7_75t_R input1023 (.A(io_ins_left_7[8]),
    .Y(net1023));
 BUFx2_ASAP7_75t_R input1024 (.A(io_ins_left_7[9]),
    .Y(net1024));
 BUFx2_ASAP7_75t_R input1025 (.A(io_ins_right_0[0]),
    .Y(net1025));
 BUFx2_ASAP7_75t_R input1026 (.A(io_ins_right_0[10]),
    .Y(net1026));
 BUFx2_ASAP7_75t_R input1027 (.A(io_ins_right_0[11]),
    .Y(net1027));
 BUFx2_ASAP7_75t_R input1028 (.A(io_ins_right_0[12]),
    .Y(net1028));
 BUFx2_ASAP7_75t_R input1029 (.A(io_ins_right_0[13]),
    .Y(net1029));
 BUFx2_ASAP7_75t_R input1030 (.A(io_ins_right_0[14]),
    .Y(net1030));
 BUFx2_ASAP7_75t_R input1031 (.A(io_ins_right_0[15]),
    .Y(net1031));
 BUFx2_ASAP7_75t_R input1032 (.A(io_ins_right_0[16]),
    .Y(net1032));
 BUFx2_ASAP7_75t_R input1033 (.A(io_ins_right_0[17]),
    .Y(net1033));
 BUFx2_ASAP7_75t_R input1034 (.A(io_ins_right_0[18]),
    .Y(net1034));
 BUFx2_ASAP7_75t_R input1035 (.A(io_ins_right_0[19]),
    .Y(net1035));
 BUFx2_ASAP7_75t_R input1036 (.A(io_ins_right_0[1]),
    .Y(net1036));
 BUFx2_ASAP7_75t_R input1037 (.A(io_ins_right_0[20]),
    .Y(net1037));
 BUFx2_ASAP7_75t_R input1038 (.A(io_ins_right_0[21]),
    .Y(net1038));
 BUFx2_ASAP7_75t_R input1039 (.A(io_ins_right_0[22]),
    .Y(net1039));
 BUFx2_ASAP7_75t_R input1040 (.A(io_ins_right_0[23]),
    .Y(net1040));
 BUFx2_ASAP7_75t_R input1041 (.A(io_ins_right_0[24]),
    .Y(net1041));
 BUFx2_ASAP7_75t_R input1042 (.A(io_ins_right_0[25]),
    .Y(net1042));
 BUFx2_ASAP7_75t_R input1043 (.A(io_ins_right_0[26]),
    .Y(net1043));
 BUFx2_ASAP7_75t_R input1044 (.A(io_ins_right_0[27]),
    .Y(net1044));
 BUFx2_ASAP7_75t_R input1045 (.A(io_ins_right_0[28]),
    .Y(net1045));
 BUFx2_ASAP7_75t_R input1046 (.A(io_ins_right_0[29]),
    .Y(net1046));
 BUFx2_ASAP7_75t_R input1047 (.A(io_ins_right_0[2]),
    .Y(net1047));
 BUFx2_ASAP7_75t_R input1048 (.A(io_ins_right_0[30]),
    .Y(net1048));
 BUFx2_ASAP7_75t_R input1049 (.A(io_ins_right_0[31]),
    .Y(net1049));
 BUFx2_ASAP7_75t_R input1050 (.A(io_ins_right_0[32]),
    .Y(net1050));
 BUFx2_ASAP7_75t_R input1051 (.A(io_ins_right_0[33]),
    .Y(net1051));
 BUFx2_ASAP7_75t_R input1052 (.A(io_ins_right_0[34]),
    .Y(net1052));
 BUFx2_ASAP7_75t_R input1053 (.A(io_ins_right_0[35]),
    .Y(net1053));
 BUFx2_ASAP7_75t_R input1054 (.A(io_ins_right_0[36]),
    .Y(net1054));
 BUFx2_ASAP7_75t_R input1055 (.A(io_ins_right_0[37]),
    .Y(net1055));
 BUFx2_ASAP7_75t_R input1056 (.A(io_ins_right_0[38]),
    .Y(net1056));
 BUFx2_ASAP7_75t_R input1057 (.A(io_ins_right_0[39]),
    .Y(net1057));
 BUFx2_ASAP7_75t_R input1058 (.A(io_ins_right_0[3]),
    .Y(net1058));
 BUFx2_ASAP7_75t_R input1059 (.A(io_ins_right_0[40]),
    .Y(net1059));
 BUFx2_ASAP7_75t_R input1060 (.A(io_ins_right_0[41]),
    .Y(net1060));
 BUFx2_ASAP7_75t_R input1061 (.A(io_ins_right_0[42]),
    .Y(net1061));
 BUFx2_ASAP7_75t_R input1062 (.A(io_ins_right_0[43]),
    .Y(net1062));
 BUFx2_ASAP7_75t_R input1063 (.A(io_ins_right_0[44]),
    .Y(net1063));
 BUFx2_ASAP7_75t_R input1064 (.A(io_ins_right_0[45]),
    .Y(net1064));
 BUFx2_ASAP7_75t_R input1065 (.A(io_ins_right_0[46]),
    .Y(net1065));
 BUFx2_ASAP7_75t_R input1066 (.A(io_ins_right_0[47]),
    .Y(net1066));
 BUFx2_ASAP7_75t_R input1067 (.A(io_ins_right_0[48]),
    .Y(net1067));
 BUFx2_ASAP7_75t_R input1068 (.A(io_ins_right_0[49]),
    .Y(net1068));
 BUFx2_ASAP7_75t_R input1069 (.A(io_ins_right_0[4]),
    .Y(net1069));
 BUFx2_ASAP7_75t_R input1070 (.A(io_ins_right_0[50]),
    .Y(net1070));
 BUFx2_ASAP7_75t_R input1071 (.A(io_ins_right_0[51]),
    .Y(net1071));
 BUFx2_ASAP7_75t_R input1072 (.A(io_ins_right_0[52]),
    .Y(net1072));
 BUFx2_ASAP7_75t_R input1073 (.A(io_ins_right_0[53]),
    .Y(net1073));
 BUFx2_ASAP7_75t_R input1074 (.A(io_ins_right_0[54]),
    .Y(net1074));
 BUFx2_ASAP7_75t_R input1075 (.A(io_ins_right_0[55]),
    .Y(net1075));
 BUFx2_ASAP7_75t_R input1076 (.A(io_ins_right_0[56]),
    .Y(net1076));
 BUFx2_ASAP7_75t_R input1077 (.A(io_ins_right_0[57]),
    .Y(net1077));
 BUFx2_ASAP7_75t_R input1078 (.A(io_ins_right_0[58]),
    .Y(net1078));
 BUFx2_ASAP7_75t_R input1079 (.A(io_ins_right_0[59]),
    .Y(net1079));
 BUFx2_ASAP7_75t_R input1080 (.A(io_ins_right_0[5]),
    .Y(net1080));
 BUFx2_ASAP7_75t_R input1081 (.A(io_ins_right_0[60]),
    .Y(net1081));
 BUFx2_ASAP7_75t_R input1082 (.A(io_ins_right_0[61]),
    .Y(net1082));
 BUFx2_ASAP7_75t_R input1083 (.A(io_ins_right_0[62]),
    .Y(net1083));
 BUFx2_ASAP7_75t_R input1084 (.A(io_ins_right_0[63]),
    .Y(net1084));
 BUFx2_ASAP7_75t_R input1085 (.A(io_ins_right_0[6]),
    .Y(net1085));
 BUFx2_ASAP7_75t_R input1086 (.A(io_ins_right_0[7]),
    .Y(net1086));
 BUFx2_ASAP7_75t_R input1087 (.A(io_ins_right_0[8]),
    .Y(net1087));
 BUFx2_ASAP7_75t_R input1088 (.A(io_ins_right_0[9]),
    .Y(net1088));
 BUFx2_ASAP7_75t_R input1089 (.A(io_ins_right_1[0]),
    .Y(net1089));
 BUFx2_ASAP7_75t_R input1090 (.A(io_ins_right_1[10]),
    .Y(net1090));
 BUFx2_ASAP7_75t_R input1091 (.A(io_ins_right_1[11]),
    .Y(net1091));
 BUFx2_ASAP7_75t_R input1092 (.A(io_ins_right_1[12]),
    .Y(net1092));
 BUFx2_ASAP7_75t_R input1093 (.A(io_ins_right_1[13]),
    .Y(net1093));
 BUFx2_ASAP7_75t_R input1094 (.A(io_ins_right_1[14]),
    .Y(net1094));
 BUFx2_ASAP7_75t_R input1095 (.A(io_ins_right_1[15]),
    .Y(net1095));
 BUFx2_ASAP7_75t_R input1096 (.A(io_ins_right_1[16]),
    .Y(net1096));
 BUFx2_ASAP7_75t_R input1097 (.A(io_ins_right_1[17]),
    .Y(net1097));
 BUFx2_ASAP7_75t_R input1098 (.A(io_ins_right_1[18]),
    .Y(net1098));
 BUFx2_ASAP7_75t_R input1099 (.A(io_ins_right_1[19]),
    .Y(net1099));
 BUFx2_ASAP7_75t_R input1100 (.A(io_ins_right_1[1]),
    .Y(net1100));
 BUFx2_ASAP7_75t_R input1101 (.A(io_ins_right_1[20]),
    .Y(net1101));
 BUFx2_ASAP7_75t_R input1102 (.A(io_ins_right_1[21]),
    .Y(net1102));
 BUFx2_ASAP7_75t_R input1103 (.A(io_ins_right_1[22]),
    .Y(net1103));
 BUFx2_ASAP7_75t_R input1104 (.A(io_ins_right_1[23]),
    .Y(net1104));
 BUFx2_ASAP7_75t_R input1105 (.A(io_ins_right_1[24]),
    .Y(net1105));
 BUFx2_ASAP7_75t_R input1106 (.A(io_ins_right_1[25]),
    .Y(net1106));
 BUFx2_ASAP7_75t_R input1107 (.A(io_ins_right_1[26]),
    .Y(net1107));
 BUFx2_ASAP7_75t_R input1108 (.A(io_ins_right_1[27]),
    .Y(net1108));
 BUFx2_ASAP7_75t_R input1109 (.A(io_ins_right_1[28]),
    .Y(net1109));
 BUFx2_ASAP7_75t_R input1110 (.A(io_ins_right_1[29]),
    .Y(net1110));
 BUFx2_ASAP7_75t_R input1111 (.A(io_ins_right_1[2]),
    .Y(net1111));
 BUFx2_ASAP7_75t_R input1112 (.A(io_ins_right_1[30]),
    .Y(net1112));
 BUFx2_ASAP7_75t_R input1113 (.A(io_ins_right_1[31]),
    .Y(net1113));
 BUFx2_ASAP7_75t_R input1114 (.A(io_ins_right_1[32]),
    .Y(net1114));
 BUFx2_ASAP7_75t_R input1115 (.A(io_ins_right_1[33]),
    .Y(net1115));
 BUFx2_ASAP7_75t_R input1116 (.A(io_ins_right_1[34]),
    .Y(net1116));
 BUFx2_ASAP7_75t_R input1117 (.A(io_ins_right_1[35]),
    .Y(net1117));
 BUFx2_ASAP7_75t_R input1118 (.A(io_ins_right_1[36]),
    .Y(net1118));
 BUFx2_ASAP7_75t_R input1119 (.A(io_ins_right_1[37]),
    .Y(net1119));
 BUFx2_ASAP7_75t_R input1120 (.A(io_ins_right_1[38]),
    .Y(net1120));
 BUFx2_ASAP7_75t_R input1121 (.A(io_ins_right_1[39]),
    .Y(net1121));
 BUFx2_ASAP7_75t_R input1122 (.A(io_ins_right_1[3]),
    .Y(net1122));
 BUFx2_ASAP7_75t_R input1123 (.A(io_ins_right_1[40]),
    .Y(net1123));
 BUFx2_ASAP7_75t_R input1124 (.A(io_ins_right_1[41]),
    .Y(net1124));
 BUFx2_ASAP7_75t_R input1125 (.A(io_ins_right_1[42]),
    .Y(net1125));
 BUFx2_ASAP7_75t_R input1126 (.A(io_ins_right_1[43]),
    .Y(net1126));
 BUFx2_ASAP7_75t_R input1127 (.A(io_ins_right_1[44]),
    .Y(net1127));
 BUFx2_ASAP7_75t_R input1128 (.A(io_ins_right_1[45]),
    .Y(net1128));
 BUFx2_ASAP7_75t_R input1129 (.A(io_ins_right_1[46]),
    .Y(net1129));
 BUFx2_ASAP7_75t_R input1130 (.A(io_ins_right_1[47]),
    .Y(net1130));
 BUFx2_ASAP7_75t_R input1131 (.A(io_ins_right_1[48]),
    .Y(net1131));
 BUFx2_ASAP7_75t_R input1132 (.A(io_ins_right_1[49]),
    .Y(net1132));
 BUFx2_ASAP7_75t_R input1133 (.A(io_ins_right_1[4]),
    .Y(net1133));
 BUFx2_ASAP7_75t_R input1134 (.A(io_ins_right_1[50]),
    .Y(net1134));
 BUFx2_ASAP7_75t_R input1135 (.A(io_ins_right_1[51]),
    .Y(net1135));
 BUFx2_ASAP7_75t_R input1136 (.A(io_ins_right_1[52]),
    .Y(net1136));
 BUFx2_ASAP7_75t_R input1137 (.A(io_ins_right_1[53]),
    .Y(net1137));
 BUFx2_ASAP7_75t_R input1138 (.A(io_ins_right_1[54]),
    .Y(net1138));
 BUFx2_ASAP7_75t_R input1139 (.A(io_ins_right_1[55]),
    .Y(net1139));
 BUFx2_ASAP7_75t_R input1140 (.A(io_ins_right_1[56]),
    .Y(net1140));
 BUFx2_ASAP7_75t_R input1141 (.A(io_ins_right_1[57]),
    .Y(net1141));
 BUFx2_ASAP7_75t_R input1142 (.A(io_ins_right_1[58]),
    .Y(net1142));
 BUFx2_ASAP7_75t_R input1143 (.A(io_ins_right_1[59]),
    .Y(net1143));
 BUFx2_ASAP7_75t_R input1144 (.A(io_ins_right_1[5]),
    .Y(net1144));
 BUFx2_ASAP7_75t_R input1145 (.A(io_ins_right_1[60]),
    .Y(net1145));
 BUFx2_ASAP7_75t_R input1146 (.A(io_ins_right_1[61]),
    .Y(net1146));
 BUFx2_ASAP7_75t_R input1147 (.A(io_ins_right_1[62]),
    .Y(net1147));
 BUFx2_ASAP7_75t_R input1148 (.A(io_ins_right_1[63]),
    .Y(net1148));
 BUFx2_ASAP7_75t_R input1149 (.A(io_ins_right_1[6]),
    .Y(net1149));
 BUFx2_ASAP7_75t_R input1150 (.A(io_ins_right_1[7]),
    .Y(net1150));
 BUFx2_ASAP7_75t_R input1151 (.A(io_ins_right_1[8]),
    .Y(net1151));
 BUFx2_ASAP7_75t_R input1152 (.A(io_ins_right_1[9]),
    .Y(net1152));
 BUFx2_ASAP7_75t_R input1153 (.A(io_ins_right_2[0]),
    .Y(net1153));
 BUFx2_ASAP7_75t_R input1154 (.A(io_ins_right_2[10]),
    .Y(net1154));
 BUFx2_ASAP7_75t_R input1155 (.A(io_ins_right_2[11]),
    .Y(net1155));
 BUFx2_ASAP7_75t_R input1156 (.A(io_ins_right_2[12]),
    .Y(net1156));
 BUFx2_ASAP7_75t_R input1157 (.A(io_ins_right_2[13]),
    .Y(net1157));
 BUFx2_ASAP7_75t_R input1158 (.A(io_ins_right_2[14]),
    .Y(net1158));
 BUFx2_ASAP7_75t_R input1159 (.A(io_ins_right_2[15]),
    .Y(net1159));
 BUFx2_ASAP7_75t_R input1160 (.A(io_ins_right_2[16]),
    .Y(net1160));
 BUFx2_ASAP7_75t_R input1161 (.A(io_ins_right_2[17]),
    .Y(net1161));
 BUFx2_ASAP7_75t_R input1162 (.A(io_ins_right_2[18]),
    .Y(net1162));
 BUFx2_ASAP7_75t_R input1163 (.A(io_ins_right_2[19]),
    .Y(net1163));
 BUFx2_ASAP7_75t_R input1164 (.A(io_ins_right_2[1]),
    .Y(net1164));
 BUFx2_ASAP7_75t_R input1165 (.A(io_ins_right_2[20]),
    .Y(net1165));
 BUFx2_ASAP7_75t_R input1166 (.A(io_ins_right_2[21]),
    .Y(net1166));
 BUFx2_ASAP7_75t_R input1167 (.A(io_ins_right_2[22]),
    .Y(net1167));
 BUFx2_ASAP7_75t_R input1168 (.A(io_ins_right_2[23]),
    .Y(net1168));
 BUFx2_ASAP7_75t_R input1169 (.A(io_ins_right_2[24]),
    .Y(net1169));
 BUFx2_ASAP7_75t_R input1170 (.A(io_ins_right_2[25]),
    .Y(net1170));
 BUFx2_ASAP7_75t_R input1171 (.A(io_ins_right_2[26]),
    .Y(net1171));
 BUFx2_ASAP7_75t_R input1172 (.A(io_ins_right_2[27]),
    .Y(net1172));
 BUFx2_ASAP7_75t_R input1173 (.A(io_ins_right_2[28]),
    .Y(net1173));
 BUFx2_ASAP7_75t_R input1174 (.A(io_ins_right_2[29]),
    .Y(net1174));
 BUFx2_ASAP7_75t_R input1175 (.A(io_ins_right_2[2]),
    .Y(net1175));
 BUFx2_ASAP7_75t_R input1176 (.A(io_ins_right_2[30]),
    .Y(net1176));
 BUFx2_ASAP7_75t_R input1177 (.A(io_ins_right_2[31]),
    .Y(net1177));
 BUFx2_ASAP7_75t_R input1178 (.A(io_ins_right_2[32]),
    .Y(net1178));
 BUFx2_ASAP7_75t_R input1179 (.A(io_ins_right_2[33]),
    .Y(net1179));
 BUFx2_ASAP7_75t_R input1180 (.A(io_ins_right_2[34]),
    .Y(net1180));
 BUFx2_ASAP7_75t_R input1181 (.A(io_ins_right_2[35]),
    .Y(net1181));
 BUFx2_ASAP7_75t_R input1182 (.A(io_ins_right_2[36]),
    .Y(net1182));
 BUFx2_ASAP7_75t_R input1183 (.A(io_ins_right_2[37]),
    .Y(net1183));
 BUFx2_ASAP7_75t_R input1184 (.A(io_ins_right_2[38]),
    .Y(net1184));
 BUFx2_ASAP7_75t_R input1185 (.A(io_ins_right_2[39]),
    .Y(net1185));
 BUFx2_ASAP7_75t_R input1186 (.A(io_ins_right_2[3]),
    .Y(net1186));
 BUFx2_ASAP7_75t_R input1187 (.A(io_ins_right_2[40]),
    .Y(net1187));
 BUFx2_ASAP7_75t_R input1188 (.A(io_ins_right_2[41]),
    .Y(net1188));
 BUFx2_ASAP7_75t_R input1189 (.A(io_ins_right_2[42]),
    .Y(net1189));
 BUFx2_ASAP7_75t_R input1190 (.A(io_ins_right_2[43]),
    .Y(net1190));
 BUFx2_ASAP7_75t_R input1191 (.A(io_ins_right_2[44]),
    .Y(net1191));
 BUFx2_ASAP7_75t_R input1192 (.A(io_ins_right_2[45]),
    .Y(net1192));
 BUFx2_ASAP7_75t_R input1193 (.A(io_ins_right_2[46]),
    .Y(net1193));
 BUFx2_ASAP7_75t_R input1194 (.A(io_ins_right_2[47]),
    .Y(net1194));
 BUFx2_ASAP7_75t_R input1195 (.A(io_ins_right_2[48]),
    .Y(net1195));
 BUFx2_ASAP7_75t_R input1196 (.A(io_ins_right_2[49]),
    .Y(net1196));
 BUFx2_ASAP7_75t_R input1197 (.A(io_ins_right_2[4]),
    .Y(net1197));
 BUFx2_ASAP7_75t_R input1198 (.A(io_ins_right_2[50]),
    .Y(net1198));
 BUFx2_ASAP7_75t_R input1199 (.A(io_ins_right_2[51]),
    .Y(net1199));
 BUFx2_ASAP7_75t_R input1200 (.A(io_ins_right_2[52]),
    .Y(net1200));
 BUFx2_ASAP7_75t_R input1201 (.A(io_ins_right_2[53]),
    .Y(net1201));
 BUFx2_ASAP7_75t_R input1202 (.A(io_ins_right_2[54]),
    .Y(net1202));
 BUFx2_ASAP7_75t_R input1203 (.A(io_ins_right_2[55]),
    .Y(net1203));
 BUFx2_ASAP7_75t_R input1204 (.A(io_ins_right_2[56]),
    .Y(net1204));
 BUFx2_ASAP7_75t_R input1205 (.A(io_ins_right_2[57]),
    .Y(net1205));
 BUFx2_ASAP7_75t_R input1206 (.A(io_ins_right_2[58]),
    .Y(net1206));
 BUFx2_ASAP7_75t_R input1207 (.A(io_ins_right_2[59]),
    .Y(net1207));
 BUFx2_ASAP7_75t_R input1208 (.A(io_ins_right_2[5]),
    .Y(net1208));
 BUFx2_ASAP7_75t_R input1209 (.A(io_ins_right_2[60]),
    .Y(net1209));
 BUFx2_ASAP7_75t_R input1210 (.A(io_ins_right_2[61]),
    .Y(net1210));
 BUFx2_ASAP7_75t_R input1211 (.A(io_ins_right_2[62]),
    .Y(net1211));
 BUFx2_ASAP7_75t_R input1212 (.A(io_ins_right_2[63]),
    .Y(net1212));
 BUFx2_ASAP7_75t_R input1213 (.A(io_ins_right_2[6]),
    .Y(net1213));
 BUFx2_ASAP7_75t_R input1214 (.A(io_ins_right_2[7]),
    .Y(net1214));
 BUFx2_ASAP7_75t_R input1215 (.A(io_ins_right_2[8]),
    .Y(net1215));
 BUFx2_ASAP7_75t_R input1216 (.A(io_ins_right_2[9]),
    .Y(net1216));
 BUFx2_ASAP7_75t_R input1217 (.A(io_ins_right_3[0]),
    .Y(net1217));
 BUFx2_ASAP7_75t_R input1218 (.A(io_ins_right_3[10]),
    .Y(net1218));
 BUFx2_ASAP7_75t_R input1219 (.A(io_ins_right_3[11]),
    .Y(net1219));
 BUFx2_ASAP7_75t_R input1220 (.A(io_ins_right_3[12]),
    .Y(net1220));
 BUFx2_ASAP7_75t_R input1221 (.A(io_ins_right_3[13]),
    .Y(net1221));
 BUFx2_ASAP7_75t_R input1222 (.A(io_ins_right_3[14]),
    .Y(net1222));
 BUFx2_ASAP7_75t_R input1223 (.A(io_ins_right_3[15]),
    .Y(net1223));
 BUFx2_ASAP7_75t_R input1224 (.A(io_ins_right_3[16]),
    .Y(net1224));
 BUFx2_ASAP7_75t_R input1225 (.A(io_ins_right_3[17]),
    .Y(net1225));
 BUFx2_ASAP7_75t_R input1226 (.A(io_ins_right_3[18]),
    .Y(net1226));
 BUFx2_ASAP7_75t_R input1227 (.A(io_ins_right_3[19]),
    .Y(net1227));
 BUFx2_ASAP7_75t_R input1228 (.A(io_ins_right_3[1]),
    .Y(net1228));
 BUFx2_ASAP7_75t_R input1229 (.A(io_ins_right_3[20]),
    .Y(net1229));
 BUFx2_ASAP7_75t_R input1230 (.A(io_ins_right_3[21]),
    .Y(net1230));
 BUFx2_ASAP7_75t_R input1231 (.A(io_ins_right_3[22]),
    .Y(net1231));
 BUFx2_ASAP7_75t_R input1232 (.A(io_ins_right_3[23]),
    .Y(net1232));
 BUFx2_ASAP7_75t_R input1233 (.A(io_ins_right_3[24]),
    .Y(net1233));
 BUFx2_ASAP7_75t_R input1234 (.A(io_ins_right_3[25]),
    .Y(net1234));
 BUFx2_ASAP7_75t_R input1235 (.A(io_ins_right_3[26]),
    .Y(net1235));
 BUFx2_ASAP7_75t_R input1236 (.A(io_ins_right_3[27]),
    .Y(net1236));
 BUFx2_ASAP7_75t_R input1237 (.A(io_ins_right_3[28]),
    .Y(net1237));
 BUFx2_ASAP7_75t_R input1238 (.A(io_ins_right_3[29]),
    .Y(net1238));
 BUFx2_ASAP7_75t_R input1239 (.A(io_ins_right_3[2]),
    .Y(net1239));
 BUFx2_ASAP7_75t_R input1240 (.A(io_ins_right_3[30]),
    .Y(net1240));
 BUFx2_ASAP7_75t_R input1241 (.A(io_ins_right_3[31]),
    .Y(net1241));
 BUFx2_ASAP7_75t_R input1242 (.A(io_ins_right_3[32]),
    .Y(net1242));
 BUFx2_ASAP7_75t_R input1243 (.A(io_ins_right_3[33]),
    .Y(net1243));
 BUFx2_ASAP7_75t_R input1244 (.A(io_ins_right_3[34]),
    .Y(net1244));
 BUFx2_ASAP7_75t_R input1245 (.A(io_ins_right_3[35]),
    .Y(net1245));
 BUFx2_ASAP7_75t_R input1246 (.A(io_ins_right_3[36]),
    .Y(net1246));
 BUFx2_ASAP7_75t_R input1247 (.A(io_ins_right_3[37]),
    .Y(net1247));
 BUFx2_ASAP7_75t_R input1248 (.A(io_ins_right_3[38]),
    .Y(net1248));
 BUFx2_ASAP7_75t_R input1249 (.A(io_ins_right_3[39]),
    .Y(net1249));
 BUFx2_ASAP7_75t_R input1250 (.A(io_ins_right_3[3]),
    .Y(net1250));
 BUFx2_ASAP7_75t_R input1251 (.A(io_ins_right_3[40]),
    .Y(net1251));
 BUFx2_ASAP7_75t_R input1252 (.A(io_ins_right_3[41]),
    .Y(net1252));
 BUFx2_ASAP7_75t_R input1253 (.A(io_ins_right_3[42]),
    .Y(net1253));
 BUFx2_ASAP7_75t_R input1254 (.A(io_ins_right_3[43]),
    .Y(net1254));
 BUFx2_ASAP7_75t_R input1255 (.A(io_ins_right_3[44]),
    .Y(net1255));
 BUFx2_ASAP7_75t_R input1256 (.A(io_ins_right_3[45]),
    .Y(net1256));
 BUFx2_ASAP7_75t_R input1257 (.A(io_ins_right_3[46]),
    .Y(net1257));
 BUFx2_ASAP7_75t_R input1258 (.A(io_ins_right_3[47]),
    .Y(net1258));
 BUFx2_ASAP7_75t_R input1259 (.A(io_ins_right_3[48]),
    .Y(net1259));
 BUFx2_ASAP7_75t_R input1260 (.A(io_ins_right_3[49]),
    .Y(net1260));
 BUFx2_ASAP7_75t_R input1261 (.A(io_ins_right_3[4]),
    .Y(net1261));
 BUFx2_ASAP7_75t_R input1262 (.A(io_ins_right_3[50]),
    .Y(net1262));
 BUFx2_ASAP7_75t_R input1263 (.A(io_ins_right_3[51]),
    .Y(net1263));
 BUFx2_ASAP7_75t_R input1264 (.A(io_ins_right_3[52]),
    .Y(net1264));
 BUFx2_ASAP7_75t_R input1265 (.A(io_ins_right_3[53]),
    .Y(net1265));
 BUFx2_ASAP7_75t_R input1266 (.A(io_ins_right_3[54]),
    .Y(net1266));
 BUFx2_ASAP7_75t_R input1267 (.A(io_ins_right_3[55]),
    .Y(net1267));
 BUFx2_ASAP7_75t_R input1268 (.A(io_ins_right_3[56]),
    .Y(net1268));
 BUFx2_ASAP7_75t_R input1269 (.A(io_ins_right_3[57]),
    .Y(net1269));
 BUFx2_ASAP7_75t_R input1270 (.A(io_ins_right_3[58]),
    .Y(net1270));
 BUFx2_ASAP7_75t_R input1271 (.A(io_ins_right_3[59]),
    .Y(net1271));
 BUFx2_ASAP7_75t_R input1272 (.A(io_ins_right_3[5]),
    .Y(net1272));
 BUFx2_ASAP7_75t_R input1273 (.A(io_ins_right_3[60]),
    .Y(net1273));
 BUFx2_ASAP7_75t_R input1274 (.A(io_ins_right_3[61]),
    .Y(net1274));
 BUFx2_ASAP7_75t_R input1275 (.A(io_ins_right_3[62]),
    .Y(net1275));
 BUFx2_ASAP7_75t_R input1276 (.A(io_ins_right_3[63]),
    .Y(net1276));
 BUFx2_ASAP7_75t_R input1277 (.A(io_ins_right_3[6]),
    .Y(net1277));
 BUFx2_ASAP7_75t_R input1278 (.A(io_ins_right_3[7]),
    .Y(net1278));
 BUFx2_ASAP7_75t_R input1279 (.A(io_ins_right_3[8]),
    .Y(net1279));
 BUFx2_ASAP7_75t_R input1280 (.A(io_ins_right_3[9]),
    .Y(net1280));
 BUFx2_ASAP7_75t_R input1281 (.A(io_ins_right_4[0]),
    .Y(net1281));
 BUFx2_ASAP7_75t_R input1282 (.A(io_ins_right_4[10]),
    .Y(net1282));
 BUFx2_ASAP7_75t_R input1283 (.A(io_ins_right_4[11]),
    .Y(net1283));
 BUFx2_ASAP7_75t_R input1284 (.A(io_ins_right_4[12]),
    .Y(net1284));
 BUFx2_ASAP7_75t_R input1285 (.A(io_ins_right_4[13]),
    .Y(net1285));
 BUFx2_ASAP7_75t_R input1286 (.A(io_ins_right_4[14]),
    .Y(net1286));
 BUFx2_ASAP7_75t_R input1287 (.A(io_ins_right_4[15]),
    .Y(net1287));
 BUFx2_ASAP7_75t_R input1288 (.A(io_ins_right_4[16]),
    .Y(net1288));
 BUFx2_ASAP7_75t_R input1289 (.A(io_ins_right_4[17]),
    .Y(net1289));
 BUFx2_ASAP7_75t_R input1290 (.A(io_ins_right_4[18]),
    .Y(net1290));
 BUFx2_ASAP7_75t_R input1291 (.A(io_ins_right_4[19]),
    .Y(net1291));
 BUFx2_ASAP7_75t_R input1292 (.A(io_ins_right_4[1]),
    .Y(net1292));
 BUFx2_ASAP7_75t_R input1293 (.A(io_ins_right_4[20]),
    .Y(net1293));
 BUFx2_ASAP7_75t_R input1294 (.A(io_ins_right_4[21]),
    .Y(net1294));
 BUFx2_ASAP7_75t_R input1295 (.A(io_ins_right_4[22]),
    .Y(net1295));
 BUFx2_ASAP7_75t_R input1296 (.A(io_ins_right_4[23]),
    .Y(net1296));
 BUFx2_ASAP7_75t_R input1297 (.A(io_ins_right_4[24]),
    .Y(net1297));
 BUFx2_ASAP7_75t_R input1298 (.A(io_ins_right_4[25]),
    .Y(net1298));
 BUFx2_ASAP7_75t_R input1299 (.A(io_ins_right_4[26]),
    .Y(net1299));
 BUFx2_ASAP7_75t_R input1300 (.A(io_ins_right_4[27]),
    .Y(net1300));
 BUFx2_ASAP7_75t_R input1301 (.A(io_ins_right_4[28]),
    .Y(net1301));
 BUFx2_ASAP7_75t_R input1302 (.A(io_ins_right_4[29]),
    .Y(net1302));
 BUFx2_ASAP7_75t_R input1303 (.A(io_ins_right_4[2]),
    .Y(net1303));
 BUFx2_ASAP7_75t_R input1304 (.A(io_ins_right_4[30]),
    .Y(net1304));
 BUFx2_ASAP7_75t_R input1305 (.A(io_ins_right_4[31]),
    .Y(net1305));
 BUFx2_ASAP7_75t_R input1306 (.A(io_ins_right_4[32]),
    .Y(net1306));
 BUFx2_ASAP7_75t_R input1307 (.A(io_ins_right_4[33]),
    .Y(net1307));
 BUFx2_ASAP7_75t_R input1308 (.A(io_ins_right_4[34]),
    .Y(net1308));
 BUFx2_ASAP7_75t_R input1309 (.A(io_ins_right_4[35]),
    .Y(net1309));
 BUFx2_ASAP7_75t_R input1310 (.A(io_ins_right_4[36]),
    .Y(net1310));
 BUFx2_ASAP7_75t_R input1311 (.A(io_ins_right_4[37]),
    .Y(net1311));
 BUFx2_ASAP7_75t_R input1312 (.A(io_ins_right_4[38]),
    .Y(net1312));
 BUFx2_ASAP7_75t_R input1313 (.A(io_ins_right_4[39]),
    .Y(net1313));
 BUFx2_ASAP7_75t_R input1314 (.A(io_ins_right_4[3]),
    .Y(net1314));
 BUFx2_ASAP7_75t_R input1315 (.A(io_ins_right_4[40]),
    .Y(net1315));
 BUFx2_ASAP7_75t_R input1316 (.A(io_ins_right_4[41]),
    .Y(net1316));
 BUFx2_ASAP7_75t_R input1317 (.A(io_ins_right_4[42]),
    .Y(net1317));
 BUFx2_ASAP7_75t_R input1318 (.A(io_ins_right_4[43]),
    .Y(net1318));
 BUFx2_ASAP7_75t_R input1319 (.A(io_ins_right_4[44]),
    .Y(net1319));
 BUFx2_ASAP7_75t_R input1320 (.A(io_ins_right_4[45]),
    .Y(net1320));
 BUFx2_ASAP7_75t_R input1321 (.A(io_ins_right_4[46]),
    .Y(net1321));
 BUFx2_ASAP7_75t_R input1322 (.A(io_ins_right_4[47]),
    .Y(net1322));
 BUFx2_ASAP7_75t_R input1323 (.A(io_ins_right_4[48]),
    .Y(net1323));
 BUFx2_ASAP7_75t_R input1324 (.A(io_ins_right_4[49]),
    .Y(net1324));
 BUFx2_ASAP7_75t_R input1325 (.A(io_ins_right_4[4]),
    .Y(net1325));
 BUFx2_ASAP7_75t_R input1326 (.A(io_ins_right_4[50]),
    .Y(net1326));
 BUFx2_ASAP7_75t_R input1327 (.A(io_ins_right_4[51]),
    .Y(net1327));
 BUFx2_ASAP7_75t_R input1328 (.A(io_ins_right_4[52]),
    .Y(net1328));
 BUFx2_ASAP7_75t_R input1329 (.A(io_ins_right_4[53]),
    .Y(net1329));
 BUFx2_ASAP7_75t_R input1330 (.A(io_ins_right_4[54]),
    .Y(net1330));
 BUFx2_ASAP7_75t_R input1331 (.A(io_ins_right_4[55]),
    .Y(net1331));
 BUFx2_ASAP7_75t_R input1332 (.A(io_ins_right_4[56]),
    .Y(net1332));
 BUFx2_ASAP7_75t_R input1333 (.A(io_ins_right_4[57]),
    .Y(net1333));
 BUFx2_ASAP7_75t_R input1334 (.A(io_ins_right_4[58]),
    .Y(net1334));
 BUFx2_ASAP7_75t_R input1335 (.A(io_ins_right_4[59]),
    .Y(net1335));
 BUFx2_ASAP7_75t_R input1336 (.A(io_ins_right_4[5]),
    .Y(net1336));
 BUFx2_ASAP7_75t_R input1337 (.A(io_ins_right_4[60]),
    .Y(net1337));
 BUFx2_ASAP7_75t_R input1338 (.A(io_ins_right_4[61]),
    .Y(net1338));
 BUFx2_ASAP7_75t_R input1339 (.A(io_ins_right_4[62]),
    .Y(net1339));
 BUFx2_ASAP7_75t_R input1340 (.A(io_ins_right_4[63]),
    .Y(net1340));
 BUFx2_ASAP7_75t_R input1341 (.A(io_ins_right_4[6]),
    .Y(net1341));
 BUFx2_ASAP7_75t_R input1342 (.A(io_ins_right_4[7]),
    .Y(net1342));
 BUFx2_ASAP7_75t_R input1343 (.A(io_ins_right_4[8]),
    .Y(net1343));
 BUFx2_ASAP7_75t_R input1344 (.A(io_ins_right_4[9]),
    .Y(net1344));
 BUFx2_ASAP7_75t_R input1345 (.A(io_ins_right_5[0]),
    .Y(net1345));
 BUFx2_ASAP7_75t_R input1346 (.A(io_ins_right_5[10]),
    .Y(net1346));
 BUFx2_ASAP7_75t_R input1347 (.A(io_ins_right_5[11]),
    .Y(net1347));
 BUFx2_ASAP7_75t_R input1348 (.A(io_ins_right_5[12]),
    .Y(net1348));
 BUFx2_ASAP7_75t_R input1349 (.A(io_ins_right_5[13]),
    .Y(net1349));
 BUFx2_ASAP7_75t_R input1350 (.A(io_ins_right_5[14]),
    .Y(net1350));
 BUFx2_ASAP7_75t_R input1351 (.A(io_ins_right_5[15]),
    .Y(net1351));
 BUFx2_ASAP7_75t_R input1352 (.A(io_ins_right_5[16]),
    .Y(net1352));
 BUFx2_ASAP7_75t_R input1353 (.A(io_ins_right_5[17]),
    .Y(net1353));
 BUFx2_ASAP7_75t_R input1354 (.A(io_ins_right_5[18]),
    .Y(net1354));
 BUFx2_ASAP7_75t_R input1355 (.A(io_ins_right_5[19]),
    .Y(net1355));
 BUFx2_ASAP7_75t_R input1356 (.A(io_ins_right_5[1]),
    .Y(net1356));
 BUFx2_ASAP7_75t_R input1357 (.A(io_ins_right_5[20]),
    .Y(net1357));
 BUFx2_ASAP7_75t_R input1358 (.A(io_ins_right_5[21]),
    .Y(net1358));
 BUFx2_ASAP7_75t_R input1359 (.A(io_ins_right_5[22]),
    .Y(net1359));
 BUFx2_ASAP7_75t_R input1360 (.A(io_ins_right_5[23]),
    .Y(net1360));
 BUFx2_ASAP7_75t_R input1361 (.A(io_ins_right_5[24]),
    .Y(net1361));
 BUFx2_ASAP7_75t_R input1362 (.A(io_ins_right_5[25]),
    .Y(net1362));
 BUFx2_ASAP7_75t_R input1363 (.A(io_ins_right_5[26]),
    .Y(net1363));
 BUFx2_ASAP7_75t_R input1364 (.A(io_ins_right_5[27]),
    .Y(net1364));
 BUFx2_ASAP7_75t_R input1365 (.A(io_ins_right_5[28]),
    .Y(net1365));
 BUFx2_ASAP7_75t_R input1366 (.A(io_ins_right_5[29]),
    .Y(net1366));
 BUFx2_ASAP7_75t_R input1367 (.A(io_ins_right_5[2]),
    .Y(net1367));
 BUFx2_ASAP7_75t_R input1368 (.A(io_ins_right_5[30]),
    .Y(net1368));
 BUFx2_ASAP7_75t_R input1369 (.A(io_ins_right_5[31]),
    .Y(net1369));
 BUFx2_ASAP7_75t_R input1370 (.A(io_ins_right_5[32]),
    .Y(net1370));
 BUFx2_ASAP7_75t_R input1371 (.A(io_ins_right_5[33]),
    .Y(net1371));
 BUFx2_ASAP7_75t_R input1372 (.A(io_ins_right_5[34]),
    .Y(net1372));
 BUFx2_ASAP7_75t_R input1373 (.A(io_ins_right_5[35]),
    .Y(net1373));
 BUFx2_ASAP7_75t_R input1374 (.A(io_ins_right_5[36]),
    .Y(net1374));
 BUFx2_ASAP7_75t_R input1375 (.A(io_ins_right_5[37]),
    .Y(net1375));
 BUFx2_ASAP7_75t_R input1376 (.A(io_ins_right_5[38]),
    .Y(net1376));
 BUFx2_ASAP7_75t_R input1377 (.A(io_ins_right_5[39]),
    .Y(net1377));
 BUFx2_ASAP7_75t_R input1378 (.A(io_ins_right_5[3]),
    .Y(net1378));
 BUFx2_ASAP7_75t_R input1379 (.A(io_ins_right_5[40]),
    .Y(net1379));
 BUFx2_ASAP7_75t_R input1380 (.A(io_ins_right_5[41]),
    .Y(net1380));
 BUFx2_ASAP7_75t_R input1381 (.A(io_ins_right_5[42]),
    .Y(net1381));
 BUFx2_ASAP7_75t_R input1382 (.A(io_ins_right_5[43]),
    .Y(net1382));
 BUFx2_ASAP7_75t_R input1383 (.A(io_ins_right_5[44]),
    .Y(net1383));
 BUFx2_ASAP7_75t_R input1384 (.A(io_ins_right_5[45]),
    .Y(net1384));
 BUFx2_ASAP7_75t_R input1385 (.A(io_ins_right_5[46]),
    .Y(net1385));
 BUFx2_ASAP7_75t_R input1386 (.A(io_ins_right_5[47]),
    .Y(net1386));
 BUFx2_ASAP7_75t_R input1387 (.A(io_ins_right_5[48]),
    .Y(net1387));
 BUFx2_ASAP7_75t_R input1388 (.A(io_ins_right_5[49]),
    .Y(net1388));
 BUFx2_ASAP7_75t_R input1389 (.A(io_ins_right_5[4]),
    .Y(net1389));
 BUFx2_ASAP7_75t_R input1390 (.A(io_ins_right_5[50]),
    .Y(net1390));
 BUFx2_ASAP7_75t_R input1391 (.A(io_ins_right_5[51]),
    .Y(net1391));
 BUFx2_ASAP7_75t_R input1392 (.A(io_ins_right_5[52]),
    .Y(net1392));
 BUFx2_ASAP7_75t_R input1393 (.A(io_ins_right_5[53]),
    .Y(net1393));
 BUFx2_ASAP7_75t_R input1394 (.A(io_ins_right_5[54]),
    .Y(net1394));
 BUFx2_ASAP7_75t_R input1395 (.A(io_ins_right_5[55]),
    .Y(net1395));
 BUFx2_ASAP7_75t_R input1396 (.A(io_ins_right_5[56]),
    .Y(net1396));
 BUFx2_ASAP7_75t_R input1397 (.A(io_ins_right_5[57]),
    .Y(net1397));
 BUFx2_ASAP7_75t_R input1398 (.A(io_ins_right_5[58]),
    .Y(net1398));
 BUFx2_ASAP7_75t_R input1399 (.A(io_ins_right_5[59]),
    .Y(net1399));
 BUFx2_ASAP7_75t_R input1400 (.A(io_ins_right_5[5]),
    .Y(net1400));
 BUFx2_ASAP7_75t_R input1401 (.A(io_ins_right_5[60]),
    .Y(net1401));
 BUFx2_ASAP7_75t_R input1402 (.A(io_ins_right_5[61]),
    .Y(net1402));
 BUFx2_ASAP7_75t_R input1403 (.A(io_ins_right_5[62]),
    .Y(net1403));
 BUFx2_ASAP7_75t_R input1404 (.A(io_ins_right_5[63]),
    .Y(net1404));
 BUFx2_ASAP7_75t_R input1405 (.A(io_ins_right_5[6]),
    .Y(net1405));
 BUFx2_ASAP7_75t_R input1406 (.A(io_ins_right_5[7]),
    .Y(net1406));
 BUFx2_ASAP7_75t_R input1407 (.A(io_ins_right_5[8]),
    .Y(net1407));
 BUFx2_ASAP7_75t_R input1408 (.A(io_ins_right_5[9]),
    .Y(net1408));
 BUFx2_ASAP7_75t_R input1409 (.A(io_ins_right_6[0]),
    .Y(net1409));
 BUFx2_ASAP7_75t_R input1410 (.A(io_ins_right_6[10]),
    .Y(net1410));
 BUFx2_ASAP7_75t_R input1411 (.A(io_ins_right_6[11]),
    .Y(net1411));
 BUFx2_ASAP7_75t_R input1412 (.A(io_ins_right_6[12]),
    .Y(net1412));
 BUFx2_ASAP7_75t_R input1413 (.A(io_ins_right_6[13]),
    .Y(net1413));
 BUFx2_ASAP7_75t_R input1414 (.A(io_ins_right_6[14]),
    .Y(net1414));
 BUFx2_ASAP7_75t_R input1415 (.A(io_ins_right_6[15]),
    .Y(net1415));
 BUFx2_ASAP7_75t_R input1416 (.A(io_ins_right_6[16]),
    .Y(net1416));
 BUFx2_ASAP7_75t_R input1417 (.A(io_ins_right_6[17]),
    .Y(net1417));
 BUFx2_ASAP7_75t_R input1418 (.A(io_ins_right_6[18]),
    .Y(net1418));
 BUFx2_ASAP7_75t_R input1419 (.A(io_ins_right_6[19]),
    .Y(net1419));
 BUFx2_ASAP7_75t_R input1420 (.A(io_ins_right_6[1]),
    .Y(net1420));
 BUFx2_ASAP7_75t_R input1421 (.A(io_ins_right_6[20]),
    .Y(net1421));
 BUFx2_ASAP7_75t_R input1422 (.A(io_ins_right_6[21]),
    .Y(net1422));
 BUFx2_ASAP7_75t_R input1423 (.A(io_ins_right_6[22]),
    .Y(net1423));
 BUFx2_ASAP7_75t_R input1424 (.A(io_ins_right_6[23]),
    .Y(net1424));
 BUFx2_ASAP7_75t_R input1425 (.A(io_ins_right_6[24]),
    .Y(net1425));
 BUFx2_ASAP7_75t_R input1426 (.A(io_ins_right_6[25]),
    .Y(net1426));
 BUFx2_ASAP7_75t_R input1427 (.A(io_ins_right_6[26]),
    .Y(net1427));
 BUFx2_ASAP7_75t_R input1428 (.A(io_ins_right_6[27]),
    .Y(net1428));
 BUFx2_ASAP7_75t_R input1429 (.A(io_ins_right_6[28]),
    .Y(net1429));
 BUFx2_ASAP7_75t_R input1430 (.A(io_ins_right_6[29]),
    .Y(net1430));
 BUFx2_ASAP7_75t_R input1431 (.A(io_ins_right_6[2]),
    .Y(net1431));
 BUFx2_ASAP7_75t_R input1432 (.A(io_ins_right_6[30]),
    .Y(net1432));
 BUFx2_ASAP7_75t_R input1433 (.A(io_ins_right_6[31]),
    .Y(net1433));
 BUFx2_ASAP7_75t_R input1434 (.A(io_ins_right_6[32]),
    .Y(net1434));
 BUFx2_ASAP7_75t_R input1435 (.A(io_ins_right_6[33]),
    .Y(net1435));
 BUFx2_ASAP7_75t_R input1436 (.A(io_ins_right_6[34]),
    .Y(net1436));
 BUFx2_ASAP7_75t_R input1437 (.A(io_ins_right_6[35]),
    .Y(net1437));
 BUFx2_ASAP7_75t_R input1438 (.A(io_ins_right_6[36]),
    .Y(net1438));
 BUFx2_ASAP7_75t_R input1439 (.A(io_ins_right_6[37]),
    .Y(net1439));
 BUFx2_ASAP7_75t_R input1440 (.A(io_ins_right_6[38]),
    .Y(net1440));
 BUFx2_ASAP7_75t_R input1441 (.A(io_ins_right_6[39]),
    .Y(net1441));
 BUFx2_ASAP7_75t_R input1442 (.A(io_ins_right_6[3]),
    .Y(net1442));
 BUFx2_ASAP7_75t_R input1443 (.A(io_ins_right_6[40]),
    .Y(net1443));
 BUFx2_ASAP7_75t_R input1444 (.A(io_ins_right_6[41]),
    .Y(net1444));
 BUFx2_ASAP7_75t_R input1445 (.A(io_ins_right_6[42]),
    .Y(net1445));
 BUFx2_ASAP7_75t_R input1446 (.A(io_ins_right_6[43]),
    .Y(net1446));
 BUFx2_ASAP7_75t_R input1447 (.A(io_ins_right_6[44]),
    .Y(net1447));
 BUFx2_ASAP7_75t_R input1448 (.A(io_ins_right_6[45]),
    .Y(net1448));
 BUFx2_ASAP7_75t_R input1449 (.A(io_ins_right_6[46]),
    .Y(net1449));
 BUFx2_ASAP7_75t_R input1450 (.A(io_ins_right_6[47]),
    .Y(net1450));
 BUFx2_ASAP7_75t_R input1451 (.A(io_ins_right_6[48]),
    .Y(net1451));
 BUFx2_ASAP7_75t_R input1452 (.A(io_ins_right_6[49]),
    .Y(net1452));
 BUFx2_ASAP7_75t_R input1453 (.A(io_ins_right_6[4]),
    .Y(net1453));
 BUFx2_ASAP7_75t_R input1454 (.A(io_ins_right_6[50]),
    .Y(net1454));
 BUFx2_ASAP7_75t_R input1455 (.A(io_ins_right_6[51]),
    .Y(net1455));
 BUFx2_ASAP7_75t_R input1456 (.A(io_ins_right_6[52]),
    .Y(net1456));
 BUFx2_ASAP7_75t_R input1457 (.A(io_ins_right_6[53]),
    .Y(net1457));
 BUFx2_ASAP7_75t_R input1458 (.A(io_ins_right_6[54]),
    .Y(net1458));
 BUFx2_ASAP7_75t_R input1459 (.A(io_ins_right_6[55]),
    .Y(net1459));
 BUFx2_ASAP7_75t_R input1460 (.A(io_ins_right_6[56]),
    .Y(net1460));
 BUFx2_ASAP7_75t_R input1461 (.A(io_ins_right_6[57]),
    .Y(net1461));
 BUFx2_ASAP7_75t_R input1462 (.A(io_ins_right_6[58]),
    .Y(net1462));
 BUFx2_ASAP7_75t_R input1463 (.A(io_ins_right_6[59]),
    .Y(net1463));
 BUFx2_ASAP7_75t_R input1464 (.A(io_ins_right_6[5]),
    .Y(net1464));
 BUFx2_ASAP7_75t_R input1465 (.A(io_ins_right_6[60]),
    .Y(net1465));
 BUFx2_ASAP7_75t_R input1466 (.A(io_ins_right_6[61]),
    .Y(net1466));
 BUFx2_ASAP7_75t_R input1467 (.A(io_ins_right_6[62]),
    .Y(net1467));
 BUFx2_ASAP7_75t_R input1468 (.A(io_ins_right_6[63]),
    .Y(net1468));
 BUFx2_ASAP7_75t_R input1469 (.A(io_ins_right_6[6]),
    .Y(net1469));
 BUFx2_ASAP7_75t_R input1470 (.A(io_ins_right_6[7]),
    .Y(net1470));
 BUFx2_ASAP7_75t_R input1471 (.A(io_ins_right_6[8]),
    .Y(net1471));
 BUFx2_ASAP7_75t_R input1472 (.A(io_ins_right_6[9]),
    .Y(net1472));
 BUFx2_ASAP7_75t_R input1473 (.A(io_ins_right_7[0]),
    .Y(net1473));
 BUFx2_ASAP7_75t_R input1474 (.A(io_ins_right_7[10]),
    .Y(net1474));
 BUFx2_ASAP7_75t_R input1475 (.A(io_ins_right_7[11]),
    .Y(net1475));
 BUFx2_ASAP7_75t_R input1476 (.A(io_ins_right_7[12]),
    .Y(net1476));
 BUFx2_ASAP7_75t_R input1477 (.A(io_ins_right_7[13]),
    .Y(net1477));
 BUFx2_ASAP7_75t_R input1478 (.A(io_ins_right_7[14]),
    .Y(net1478));
 BUFx2_ASAP7_75t_R input1479 (.A(io_ins_right_7[15]),
    .Y(net1479));
 BUFx2_ASAP7_75t_R input1480 (.A(io_ins_right_7[16]),
    .Y(net1480));
 BUFx2_ASAP7_75t_R input1481 (.A(io_ins_right_7[17]),
    .Y(net1481));
 BUFx2_ASAP7_75t_R input1482 (.A(io_ins_right_7[18]),
    .Y(net1482));
 BUFx2_ASAP7_75t_R input1483 (.A(io_ins_right_7[19]),
    .Y(net1483));
 BUFx2_ASAP7_75t_R input1484 (.A(io_ins_right_7[1]),
    .Y(net1484));
 BUFx2_ASAP7_75t_R input1485 (.A(io_ins_right_7[20]),
    .Y(net1485));
 BUFx2_ASAP7_75t_R input1486 (.A(io_ins_right_7[21]),
    .Y(net1486));
 BUFx2_ASAP7_75t_R input1487 (.A(io_ins_right_7[22]),
    .Y(net1487));
 BUFx2_ASAP7_75t_R input1488 (.A(io_ins_right_7[23]),
    .Y(net1488));
 BUFx2_ASAP7_75t_R input1489 (.A(io_ins_right_7[24]),
    .Y(net1489));
 BUFx2_ASAP7_75t_R input1490 (.A(io_ins_right_7[25]),
    .Y(net1490));
 BUFx2_ASAP7_75t_R input1491 (.A(io_ins_right_7[26]),
    .Y(net1491));
 BUFx2_ASAP7_75t_R input1492 (.A(io_ins_right_7[27]),
    .Y(net1492));
 BUFx2_ASAP7_75t_R input1493 (.A(io_ins_right_7[28]),
    .Y(net1493));
 BUFx2_ASAP7_75t_R input1494 (.A(io_ins_right_7[29]),
    .Y(net1494));
 BUFx2_ASAP7_75t_R input1495 (.A(io_ins_right_7[2]),
    .Y(net1495));
 BUFx2_ASAP7_75t_R input1496 (.A(io_ins_right_7[30]),
    .Y(net1496));
 BUFx2_ASAP7_75t_R input1497 (.A(io_ins_right_7[31]),
    .Y(net1497));
 BUFx2_ASAP7_75t_R input1498 (.A(io_ins_right_7[32]),
    .Y(net1498));
 BUFx2_ASAP7_75t_R input1499 (.A(io_ins_right_7[33]),
    .Y(net1499));
 BUFx2_ASAP7_75t_R input1500 (.A(io_ins_right_7[34]),
    .Y(net1500));
 BUFx2_ASAP7_75t_R input1501 (.A(io_ins_right_7[35]),
    .Y(net1501));
 BUFx2_ASAP7_75t_R input1502 (.A(io_ins_right_7[36]),
    .Y(net1502));
 BUFx2_ASAP7_75t_R input1503 (.A(io_ins_right_7[37]),
    .Y(net1503));
 BUFx2_ASAP7_75t_R input1504 (.A(io_ins_right_7[38]),
    .Y(net1504));
 BUFx2_ASAP7_75t_R input1505 (.A(io_ins_right_7[39]),
    .Y(net1505));
 BUFx2_ASAP7_75t_R input1506 (.A(io_ins_right_7[3]),
    .Y(net1506));
 BUFx2_ASAP7_75t_R input1507 (.A(io_ins_right_7[40]),
    .Y(net1507));
 BUFx2_ASAP7_75t_R input1508 (.A(io_ins_right_7[41]),
    .Y(net1508));
 BUFx2_ASAP7_75t_R input1509 (.A(io_ins_right_7[42]),
    .Y(net1509));
 BUFx2_ASAP7_75t_R input1510 (.A(io_ins_right_7[43]),
    .Y(net1510));
 BUFx2_ASAP7_75t_R input1511 (.A(io_ins_right_7[44]),
    .Y(net1511));
 BUFx2_ASAP7_75t_R input1512 (.A(io_ins_right_7[45]),
    .Y(net1512));
 BUFx2_ASAP7_75t_R input1513 (.A(io_ins_right_7[46]),
    .Y(net1513));
 BUFx2_ASAP7_75t_R input1514 (.A(io_ins_right_7[47]),
    .Y(net1514));
 BUFx2_ASAP7_75t_R input1515 (.A(io_ins_right_7[48]),
    .Y(net1515));
 BUFx2_ASAP7_75t_R input1516 (.A(io_ins_right_7[49]),
    .Y(net1516));
 BUFx2_ASAP7_75t_R input1517 (.A(io_ins_right_7[4]),
    .Y(net1517));
 BUFx2_ASAP7_75t_R input1518 (.A(io_ins_right_7[50]),
    .Y(net1518));
 BUFx2_ASAP7_75t_R input1519 (.A(io_ins_right_7[51]),
    .Y(net1519));
 BUFx2_ASAP7_75t_R input1520 (.A(io_ins_right_7[52]),
    .Y(net1520));
 BUFx2_ASAP7_75t_R input1521 (.A(io_ins_right_7[53]),
    .Y(net1521));
 BUFx2_ASAP7_75t_R input1522 (.A(io_ins_right_7[54]),
    .Y(net1522));
 BUFx2_ASAP7_75t_R input1523 (.A(io_ins_right_7[55]),
    .Y(net1523));
 BUFx2_ASAP7_75t_R input1524 (.A(io_ins_right_7[56]),
    .Y(net1524));
 BUFx2_ASAP7_75t_R input1525 (.A(io_ins_right_7[57]),
    .Y(net1525));
 BUFx2_ASAP7_75t_R input1526 (.A(io_ins_right_7[58]),
    .Y(net1526));
 BUFx2_ASAP7_75t_R input1527 (.A(io_ins_right_7[59]),
    .Y(net1527));
 BUFx2_ASAP7_75t_R input1528 (.A(io_ins_right_7[5]),
    .Y(net1528));
 BUFx2_ASAP7_75t_R input1529 (.A(io_ins_right_7[60]),
    .Y(net1529));
 BUFx2_ASAP7_75t_R input1530 (.A(io_ins_right_7[61]),
    .Y(net1530));
 BUFx2_ASAP7_75t_R input1531 (.A(io_ins_right_7[62]),
    .Y(net1531));
 BUFx2_ASAP7_75t_R input1532 (.A(io_ins_right_7[63]),
    .Y(net1532));
 BUFx2_ASAP7_75t_R input1533 (.A(io_ins_right_7[6]),
    .Y(net1533));
 BUFx2_ASAP7_75t_R input1534 (.A(io_ins_right_7[7]),
    .Y(net1534));
 BUFx2_ASAP7_75t_R input1535 (.A(io_ins_right_7[8]),
    .Y(net1535));
 BUFx2_ASAP7_75t_R input1536 (.A(io_ins_right_7[9]),
    .Y(net1536));
 BUFx2_ASAP7_75t_R input1537 (.A(io_ins_up_0[0]),
    .Y(net1537));
 BUFx2_ASAP7_75t_R input1538 (.A(io_ins_up_0[10]),
    .Y(net1538));
 BUFx2_ASAP7_75t_R input1539 (.A(io_ins_up_0[11]),
    .Y(net1539));
 BUFx2_ASAP7_75t_R input1540 (.A(io_ins_up_0[12]),
    .Y(net1540));
 BUFx2_ASAP7_75t_R input1541 (.A(io_ins_up_0[13]),
    .Y(net1541));
 BUFx2_ASAP7_75t_R input1542 (.A(io_ins_up_0[14]),
    .Y(net1542));
 BUFx2_ASAP7_75t_R input1543 (.A(io_ins_up_0[15]),
    .Y(net1543));
 BUFx2_ASAP7_75t_R input1544 (.A(io_ins_up_0[16]),
    .Y(net1544));
 BUFx2_ASAP7_75t_R input1545 (.A(io_ins_up_0[17]),
    .Y(net1545));
 BUFx2_ASAP7_75t_R input1546 (.A(io_ins_up_0[18]),
    .Y(net1546));
 BUFx2_ASAP7_75t_R input1547 (.A(io_ins_up_0[19]),
    .Y(net1547));
 BUFx2_ASAP7_75t_R input1548 (.A(io_ins_up_0[1]),
    .Y(net1548));
 BUFx2_ASAP7_75t_R input1549 (.A(io_ins_up_0[20]),
    .Y(net1549));
 BUFx2_ASAP7_75t_R input1550 (.A(io_ins_up_0[21]),
    .Y(net1550));
 BUFx2_ASAP7_75t_R input1551 (.A(io_ins_up_0[22]),
    .Y(net1551));
 BUFx2_ASAP7_75t_R input1552 (.A(io_ins_up_0[23]),
    .Y(net1552));
 BUFx2_ASAP7_75t_R input1553 (.A(io_ins_up_0[24]),
    .Y(net1553));
 BUFx2_ASAP7_75t_R input1554 (.A(io_ins_up_0[25]),
    .Y(net1554));
 BUFx2_ASAP7_75t_R input1555 (.A(io_ins_up_0[26]),
    .Y(net1555));
 BUFx2_ASAP7_75t_R input1556 (.A(io_ins_up_0[27]),
    .Y(net1556));
 BUFx2_ASAP7_75t_R input1557 (.A(io_ins_up_0[28]),
    .Y(net1557));
 BUFx2_ASAP7_75t_R input1558 (.A(io_ins_up_0[29]),
    .Y(net1558));
 BUFx2_ASAP7_75t_R input1559 (.A(io_ins_up_0[2]),
    .Y(net1559));
 BUFx2_ASAP7_75t_R input1560 (.A(io_ins_up_0[30]),
    .Y(net1560));
 BUFx2_ASAP7_75t_R input1561 (.A(io_ins_up_0[31]),
    .Y(net1561));
 BUFx2_ASAP7_75t_R input1562 (.A(io_ins_up_0[32]),
    .Y(net1562));
 BUFx2_ASAP7_75t_R input1563 (.A(io_ins_up_0[33]),
    .Y(net1563));
 BUFx2_ASAP7_75t_R input1564 (.A(io_ins_up_0[34]),
    .Y(net1564));
 BUFx2_ASAP7_75t_R input1565 (.A(io_ins_up_0[35]),
    .Y(net1565));
 BUFx2_ASAP7_75t_R input1566 (.A(io_ins_up_0[36]),
    .Y(net1566));
 BUFx2_ASAP7_75t_R input1567 (.A(io_ins_up_0[37]),
    .Y(net1567));
 BUFx2_ASAP7_75t_R input1568 (.A(io_ins_up_0[38]),
    .Y(net1568));
 BUFx2_ASAP7_75t_R input1569 (.A(io_ins_up_0[39]),
    .Y(net1569));
 BUFx2_ASAP7_75t_R input1570 (.A(io_ins_up_0[3]),
    .Y(net1570));
 BUFx2_ASAP7_75t_R input1571 (.A(io_ins_up_0[40]),
    .Y(net1571));
 BUFx2_ASAP7_75t_R input1572 (.A(io_ins_up_0[41]),
    .Y(net1572));
 BUFx2_ASAP7_75t_R input1573 (.A(io_ins_up_0[42]),
    .Y(net1573));
 BUFx2_ASAP7_75t_R input1574 (.A(io_ins_up_0[43]),
    .Y(net1574));
 BUFx2_ASAP7_75t_R input1575 (.A(io_ins_up_0[44]),
    .Y(net1575));
 BUFx2_ASAP7_75t_R input1576 (.A(io_ins_up_0[45]),
    .Y(net1576));
 BUFx2_ASAP7_75t_R input1577 (.A(io_ins_up_0[46]),
    .Y(net1577));
 BUFx2_ASAP7_75t_R input1578 (.A(io_ins_up_0[47]),
    .Y(net1578));
 BUFx2_ASAP7_75t_R input1579 (.A(io_ins_up_0[48]),
    .Y(net1579));
 BUFx2_ASAP7_75t_R input1580 (.A(io_ins_up_0[49]),
    .Y(net1580));
 BUFx2_ASAP7_75t_R input1581 (.A(io_ins_up_0[4]),
    .Y(net1581));
 BUFx2_ASAP7_75t_R input1582 (.A(io_ins_up_0[50]),
    .Y(net1582));
 BUFx2_ASAP7_75t_R input1583 (.A(io_ins_up_0[51]),
    .Y(net1583));
 BUFx2_ASAP7_75t_R input1584 (.A(io_ins_up_0[52]),
    .Y(net1584));
 BUFx2_ASAP7_75t_R input1585 (.A(io_ins_up_0[53]),
    .Y(net1585));
 BUFx2_ASAP7_75t_R input1586 (.A(io_ins_up_0[54]),
    .Y(net1586));
 BUFx2_ASAP7_75t_R input1587 (.A(io_ins_up_0[55]),
    .Y(net1587));
 BUFx2_ASAP7_75t_R input1588 (.A(io_ins_up_0[56]),
    .Y(net1588));
 BUFx2_ASAP7_75t_R input1589 (.A(io_ins_up_0[57]),
    .Y(net1589));
 BUFx2_ASAP7_75t_R input1590 (.A(io_ins_up_0[58]),
    .Y(net1590));
 BUFx2_ASAP7_75t_R input1591 (.A(io_ins_up_0[59]),
    .Y(net1591));
 BUFx2_ASAP7_75t_R input1592 (.A(io_ins_up_0[5]),
    .Y(net1592));
 BUFx2_ASAP7_75t_R input1593 (.A(io_ins_up_0[60]),
    .Y(net1593));
 BUFx2_ASAP7_75t_R input1594 (.A(io_ins_up_0[61]),
    .Y(net1594));
 BUFx2_ASAP7_75t_R input1595 (.A(io_ins_up_0[62]),
    .Y(net1595));
 BUFx2_ASAP7_75t_R input1596 (.A(io_ins_up_0[63]),
    .Y(net1596));
 BUFx2_ASAP7_75t_R input1597 (.A(io_ins_up_0[6]),
    .Y(net1597));
 BUFx2_ASAP7_75t_R input1598 (.A(io_ins_up_0[7]),
    .Y(net1598));
 BUFx2_ASAP7_75t_R input1599 (.A(io_ins_up_0[8]),
    .Y(net1599));
 BUFx2_ASAP7_75t_R input1600 (.A(io_ins_up_0[9]),
    .Y(net1600));
 BUFx2_ASAP7_75t_R input1601 (.A(io_ins_up_1[0]),
    .Y(net1601));
 BUFx2_ASAP7_75t_R input1602 (.A(io_ins_up_1[10]),
    .Y(net1602));
 BUFx2_ASAP7_75t_R input1603 (.A(io_ins_up_1[11]),
    .Y(net1603));
 BUFx2_ASAP7_75t_R input1604 (.A(io_ins_up_1[12]),
    .Y(net1604));
 BUFx2_ASAP7_75t_R input1605 (.A(io_ins_up_1[13]),
    .Y(net1605));
 BUFx2_ASAP7_75t_R input1606 (.A(io_ins_up_1[14]),
    .Y(net1606));
 BUFx2_ASAP7_75t_R input1607 (.A(io_ins_up_1[15]),
    .Y(net1607));
 BUFx2_ASAP7_75t_R input1608 (.A(io_ins_up_1[16]),
    .Y(net1608));
 BUFx2_ASAP7_75t_R input1609 (.A(io_ins_up_1[17]),
    .Y(net1609));
 BUFx2_ASAP7_75t_R input1610 (.A(io_ins_up_1[18]),
    .Y(net1610));
 BUFx2_ASAP7_75t_R input1611 (.A(io_ins_up_1[19]),
    .Y(net1611));
 BUFx2_ASAP7_75t_R input1612 (.A(io_ins_up_1[1]),
    .Y(net1612));
 BUFx2_ASAP7_75t_R input1613 (.A(io_ins_up_1[20]),
    .Y(net1613));
 BUFx2_ASAP7_75t_R input1614 (.A(io_ins_up_1[21]),
    .Y(net1614));
 BUFx2_ASAP7_75t_R input1615 (.A(io_ins_up_1[22]),
    .Y(net1615));
 BUFx2_ASAP7_75t_R input1616 (.A(io_ins_up_1[23]),
    .Y(net1616));
 BUFx2_ASAP7_75t_R input1617 (.A(io_ins_up_1[24]),
    .Y(net1617));
 BUFx2_ASAP7_75t_R input1618 (.A(io_ins_up_1[25]),
    .Y(net1618));
 BUFx2_ASAP7_75t_R input1619 (.A(io_ins_up_1[26]),
    .Y(net1619));
 BUFx2_ASAP7_75t_R input1620 (.A(io_ins_up_1[27]),
    .Y(net1620));
 BUFx2_ASAP7_75t_R input1621 (.A(io_ins_up_1[28]),
    .Y(net1621));
 BUFx2_ASAP7_75t_R input1622 (.A(io_ins_up_1[29]),
    .Y(net1622));
 BUFx2_ASAP7_75t_R input1623 (.A(io_ins_up_1[2]),
    .Y(net1623));
 BUFx2_ASAP7_75t_R input1624 (.A(io_ins_up_1[30]),
    .Y(net1624));
 BUFx2_ASAP7_75t_R input1625 (.A(io_ins_up_1[31]),
    .Y(net1625));
 BUFx2_ASAP7_75t_R input1626 (.A(io_ins_up_1[32]),
    .Y(net1626));
 BUFx2_ASAP7_75t_R input1627 (.A(io_ins_up_1[33]),
    .Y(net1627));
 BUFx2_ASAP7_75t_R input1628 (.A(io_ins_up_1[34]),
    .Y(net1628));
 BUFx2_ASAP7_75t_R input1629 (.A(io_ins_up_1[35]),
    .Y(net1629));
 BUFx2_ASAP7_75t_R input1630 (.A(io_ins_up_1[36]),
    .Y(net1630));
 BUFx2_ASAP7_75t_R input1631 (.A(io_ins_up_1[37]),
    .Y(net1631));
 BUFx2_ASAP7_75t_R input1632 (.A(io_ins_up_1[38]),
    .Y(net1632));
 BUFx2_ASAP7_75t_R input1633 (.A(io_ins_up_1[39]),
    .Y(net1633));
 BUFx2_ASAP7_75t_R input1634 (.A(io_ins_up_1[3]),
    .Y(net1634));
 BUFx2_ASAP7_75t_R input1635 (.A(io_ins_up_1[40]),
    .Y(net1635));
 BUFx2_ASAP7_75t_R input1636 (.A(io_ins_up_1[41]),
    .Y(net1636));
 BUFx2_ASAP7_75t_R input1637 (.A(io_ins_up_1[42]),
    .Y(net1637));
 BUFx2_ASAP7_75t_R input1638 (.A(io_ins_up_1[43]),
    .Y(net1638));
 BUFx2_ASAP7_75t_R input1639 (.A(io_ins_up_1[44]),
    .Y(net1639));
 BUFx2_ASAP7_75t_R input1640 (.A(io_ins_up_1[45]),
    .Y(net1640));
 BUFx2_ASAP7_75t_R input1641 (.A(io_ins_up_1[46]),
    .Y(net1641));
 BUFx2_ASAP7_75t_R input1642 (.A(io_ins_up_1[47]),
    .Y(net1642));
 BUFx2_ASAP7_75t_R input1643 (.A(io_ins_up_1[48]),
    .Y(net1643));
 BUFx2_ASAP7_75t_R input1644 (.A(io_ins_up_1[49]),
    .Y(net1644));
 BUFx2_ASAP7_75t_R input1645 (.A(io_ins_up_1[4]),
    .Y(net1645));
 BUFx2_ASAP7_75t_R input1646 (.A(io_ins_up_1[50]),
    .Y(net1646));
 BUFx2_ASAP7_75t_R input1647 (.A(io_ins_up_1[51]),
    .Y(net1647));
 BUFx2_ASAP7_75t_R input1648 (.A(io_ins_up_1[52]),
    .Y(net1648));
 BUFx2_ASAP7_75t_R input1649 (.A(io_ins_up_1[53]),
    .Y(net1649));
 BUFx2_ASAP7_75t_R input1650 (.A(io_ins_up_1[54]),
    .Y(net1650));
 BUFx2_ASAP7_75t_R input1651 (.A(io_ins_up_1[55]),
    .Y(net1651));
 BUFx2_ASAP7_75t_R input1652 (.A(io_ins_up_1[56]),
    .Y(net1652));
 BUFx2_ASAP7_75t_R input1653 (.A(io_ins_up_1[57]),
    .Y(net1653));
 BUFx2_ASAP7_75t_R input1654 (.A(io_ins_up_1[58]),
    .Y(net1654));
 BUFx2_ASAP7_75t_R input1655 (.A(io_ins_up_1[59]),
    .Y(net1655));
 BUFx2_ASAP7_75t_R input1656 (.A(io_ins_up_1[5]),
    .Y(net1656));
 BUFx2_ASAP7_75t_R input1657 (.A(io_ins_up_1[60]),
    .Y(net1657));
 BUFx2_ASAP7_75t_R input1658 (.A(io_ins_up_1[61]),
    .Y(net1658));
 BUFx2_ASAP7_75t_R input1659 (.A(io_ins_up_1[62]),
    .Y(net1659));
 BUFx2_ASAP7_75t_R input1660 (.A(io_ins_up_1[63]),
    .Y(net1660));
 BUFx2_ASAP7_75t_R input1661 (.A(io_ins_up_1[6]),
    .Y(net1661));
 BUFx2_ASAP7_75t_R input1662 (.A(io_ins_up_1[7]),
    .Y(net1662));
 BUFx2_ASAP7_75t_R input1663 (.A(io_ins_up_1[8]),
    .Y(net1663));
 BUFx2_ASAP7_75t_R input1664 (.A(io_ins_up_1[9]),
    .Y(net1664));
 BUFx2_ASAP7_75t_R input1665 (.A(io_ins_up_2[0]),
    .Y(net1665));
 BUFx2_ASAP7_75t_R input1666 (.A(io_ins_up_2[10]),
    .Y(net1666));
 BUFx2_ASAP7_75t_R input1667 (.A(io_ins_up_2[11]),
    .Y(net1667));
 BUFx2_ASAP7_75t_R input1668 (.A(io_ins_up_2[12]),
    .Y(net1668));
 BUFx2_ASAP7_75t_R input1669 (.A(io_ins_up_2[13]),
    .Y(net1669));
 BUFx2_ASAP7_75t_R input1670 (.A(io_ins_up_2[14]),
    .Y(net1670));
 BUFx2_ASAP7_75t_R input1671 (.A(io_ins_up_2[15]),
    .Y(net1671));
 BUFx2_ASAP7_75t_R input1672 (.A(io_ins_up_2[16]),
    .Y(net1672));
 BUFx2_ASAP7_75t_R input1673 (.A(io_ins_up_2[17]),
    .Y(net1673));
 BUFx2_ASAP7_75t_R input1674 (.A(io_ins_up_2[18]),
    .Y(net1674));
 BUFx2_ASAP7_75t_R input1675 (.A(io_ins_up_2[19]),
    .Y(net1675));
 BUFx2_ASAP7_75t_R input1676 (.A(io_ins_up_2[1]),
    .Y(net1676));
 BUFx2_ASAP7_75t_R input1677 (.A(io_ins_up_2[20]),
    .Y(net1677));
 BUFx2_ASAP7_75t_R input1678 (.A(io_ins_up_2[21]),
    .Y(net1678));
 BUFx2_ASAP7_75t_R input1679 (.A(io_ins_up_2[22]),
    .Y(net1679));
 BUFx2_ASAP7_75t_R input1680 (.A(io_ins_up_2[23]),
    .Y(net1680));
 BUFx2_ASAP7_75t_R input1681 (.A(io_ins_up_2[24]),
    .Y(net1681));
 BUFx2_ASAP7_75t_R input1682 (.A(io_ins_up_2[25]),
    .Y(net1682));
 BUFx2_ASAP7_75t_R input1683 (.A(io_ins_up_2[26]),
    .Y(net1683));
 BUFx2_ASAP7_75t_R input1684 (.A(io_ins_up_2[27]),
    .Y(net1684));
 BUFx2_ASAP7_75t_R input1685 (.A(io_ins_up_2[28]),
    .Y(net1685));
 BUFx2_ASAP7_75t_R input1686 (.A(io_ins_up_2[29]),
    .Y(net1686));
 BUFx2_ASAP7_75t_R input1687 (.A(io_ins_up_2[2]),
    .Y(net1687));
 BUFx2_ASAP7_75t_R input1688 (.A(io_ins_up_2[30]),
    .Y(net1688));
 BUFx2_ASAP7_75t_R input1689 (.A(io_ins_up_2[31]),
    .Y(net1689));
 BUFx2_ASAP7_75t_R input1690 (.A(io_ins_up_2[32]),
    .Y(net1690));
 BUFx2_ASAP7_75t_R input1691 (.A(io_ins_up_2[33]),
    .Y(net1691));
 BUFx2_ASAP7_75t_R input1692 (.A(io_ins_up_2[34]),
    .Y(net1692));
 BUFx2_ASAP7_75t_R input1693 (.A(io_ins_up_2[35]),
    .Y(net1693));
 BUFx2_ASAP7_75t_R input1694 (.A(io_ins_up_2[36]),
    .Y(net1694));
 BUFx2_ASAP7_75t_R input1695 (.A(io_ins_up_2[37]),
    .Y(net1695));
 BUFx2_ASAP7_75t_R input1696 (.A(io_ins_up_2[38]),
    .Y(net1696));
 BUFx2_ASAP7_75t_R input1697 (.A(io_ins_up_2[39]),
    .Y(net1697));
 BUFx2_ASAP7_75t_R input1698 (.A(io_ins_up_2[3]),
    .Y(net1698));
 BUFx2_ASAP7_75t_R input1699 (.A(io_ins_up_2[40]),
    .Y(net1699));
 BUFx2_ASAP7_75t_R input1700 (.A(io_ins_up_2[41]),
    .Y(net1700));
 BUFx2_ASAP7_75t_R input1701 (.A(io_ins_up_2[42]),
    .Y(net1701));
 BUFx2_ASAP7_75t_R input1702 (.A(io_ins_up_2[43]),
    .Y(net1702));
 BUFx2_ASAP7_75t_R input1703 (.A(io_ins_up_2[44]),
    .Y(net1703));
 BUFx2_ASAP7_75t_R input1704 (.A(io_ins_up_2[45]),
    .Y(net1704));
 BUFx2_ASAP7_75t_R input1705 (.A(io_ins_up_2[46]),
    .Y(net1705));
 BUFx2_ASAP7_75t_R input1706 (.A(io_ins_up_2[47]),
    .Y(net1706));
 BUFx2_ASAP7_75t_R input1707 (.A(io_ins_up_2[48]),
    .Y(net1707));
 BUFx2_ASAP7_75t_R input1708 (.A(io_ins_up_2[49]),
    .Y(net1708));
 BUFx2_ASAP7_75t_R input1709 (.A(io_ins_up_2[4]),
    .Y(net1709));
 BUFx2_ASAP7_75t_R input1710 (.A(io_ins_up_2[50]),
    .Y(net1710));
 BUFx2_ASAP7_75t_R input1711 (.A(io_ins_up_2[51]),
    .Y(net1711));
 BUFx2_ASAP7_75t_R input1712 (.A(io_ins_up_2[52]),
    .Y(net1712));
 BUFx2_ASAP7_75t_R input1713 (.A(io_ins_up_2[53]),
    .Y(net1713));
 BUFx2_ASAP7_75t_R input1714 (.A(io_ins_up_2[54]),
    .Y(net1714));
 BUFx2_ASAP7_75t_R input1715 (.A(io_ins_up_2[55]),
    .Y(net1715));
 BUFx2_ASAP7_75t_R input1716 (.A(io_ins_up_2[56]),
    .Y(net1716));
 BUFx2_ASAP7_75t_R input1717 (.A(io_ins_up_2[57]),
    .Y(net1717));
 BUFx2_ASAP7_75t_R input1718 (.A(io_ins_up_2[58]),
    .Y(net1718));
 BUFx2_ASAP7_75t_R input1719 (.A(io_ins_up_2[59]),
    .Y(net1719));
 BUFx2_ASAP7_75t_R input1720 (.A(io_ins_up_2[5]),
    .Y(net1720));
 BUFx2_ASAP7_75t_R input1721 (.A(io_ins_up_2[60]),
    .Y(net1721));
 BUFx2_ASAP7_75t_R input1722 (.A(io_ins_up_2[61]),
    .Y(net1722));
 BUFx2_ASAP7_75t_R input1723 (.A(io_ins_up_2[62]),
    .Y(net1723));
 BUFx2_ASAP7_75t_R input1724 (.A(io_ins_up_2[63]),
    .Y(net1724));
 BUFx2_ASAP7_75t_R input1725 (.A(io_ins_up_2[6]),
    .Y(net1725));
 BUFx2_ASAP7_75t_R input1726 (.A(io_ins_up_2[7]),
    .Y(net1726));
 BUFx2_ASAP7_75t_R input1727 (.A(io_ins_up_2[8]),
    .Y(net1727));
 BUFx2_ASAP7_75t_R input1728 (.A(io_ins_up_2[9]),
    .Y(net1728));
 BUFx2_ASAP7_75t_R input1729 (.A(io_ins_up_3[0]),
    .Y(net1729));
 BUFx2_ASAP7_75t_R input1730 (.A(io_ins_up_3[10]),
    .Y(net1730));
 BUFx2_ASAP7_75t_R input1731 (.A(io_ins_up_3[11]),
    .Y(net1731));
 BUFx2_ASAP7_75t_R input1732 (.A(io_ins_up_3[12]),
    .Y(net1732));
 BUFx2_ASAP7_75t_R input1733 (.A(io_ins_up_3[13]),
    .Y(net1733));
 BUFx2_ASAP7_75t_R input1734 (.A(io_ins_up_3[14]),
    .Y(net1734));
 BUFx2_ASAP7_75t_R input1735 (.A(io_ins_up_3[15]),
    .Y(net1735));
 BUFx2_ASAP7_75t_R input1736 (.A(io_ins_up_3[16]),
    .Y(net1736));
 BUFx2_ASAP7_75t_R input1737 (.A(io_ins_up_3[17]),
    .Y(net1737));
 BUFx2_ASAP7_75t_R input1738 (.A(io_ins_up_3[18]),
    .Y(net1738));
 BUFx2_ASAP7_75t_R input1739 (.A(io_ins_up_3[19]),
    .Y(net1739));
 BUFx2_ASAP7_75t_R input1740 (.A(io_ins_up_3[1]),
    .Y(net1740));
 BUFx2_ASAP7_75t_R input1741 (.A(io_ins_up_3[20]),
    .Y(net1741));
 BUFx2_ASAP7_75t_R input1742 (.A(io_ins_up_3[21]),
    .Y(net1742));
 BUFx2_ASAP7_75t_R input1743 (.A(io_ins_up_3[22]),
    .Y(net1743));
 BUFx2_ASAP7_75t_R input1744 (.A(io_ins_up_3[23]),
    .Y(net1744));
 BUFx2_ASAP7_75t_R input1745 (.A(io_ins_up_3[24]),
    .Y(net1745));
 BUFx2_ASAP7_75t_R input1746 (.A(io_ins_up_3[25]),
    .Y(net1746));
 BUFx2_ASAP7_75t_R input1747 (.A(io_ins_up_3[26]),
    .Y(net1747));
 BUFx2_ASAP7_75t_R input1748 (.A(io_ins_up_3[27]),
    .Y(net1748));
 BUFx2_ASAP7_75t_R input1749 (.A(io_ins_up_3[28]),
    .Y(net1749));
 BUFx2_ASAP7_75t_R input1750 (.A(io_ins_up_3[29]),
    .Y(net1750));
 BUFx2_ASAP7_75t_R input1751 (.A(io_ins_up_3[2]),
    .Y(net1751));
 BUFx2_ASAP7_75t_R input1752 (.A(io_ins_up_3[30]),
    .Y(net1752));
 BUFx2_ASAP7_75t_R input1753 (.A(io_ins_up_3[31]),
    .Y(net1753));
 BUFx2_ASAP7_75t_R input1754 (.A(io_ins_up_3[32]),
    .Y(net1754));
 BUFx2_ASAP7_75t_R input1755 (.A(io_ins_up_3[33]),
    .Y(net1755));
 BUFx2_ASAP7_75t_R input1756 (.A(io_ins_up_3[34]),
    .Y(net1756));
 BUFx2_ASAP7_75t_R input1757 (.A(io_ins_up_3[35]),
    .Y(net1757));
 BUFx2_ASAP7_75t_R input1758 (.A(io_ins_up_3[36]),
    .Y(net1758));
 BUFx2_ASAP7_75t_R input1759 (.A(io_ins_up_3[37]),
    .Y(net1759));
 BUFx2_ASAP7_75t_R input1760 (.A(io_ins_up_3[38]),
    .Y(net1760));
 BUFx2_ASAP7_75t_R input1761 (.A(io_ins_up_3[39]),
    .Y(net1761));
 BUFx2_ASAP7_75t_R input1762 (.A(io_ins_up_3[3]),
    .Y(net1762));
 BUFx2_ASAP7_75t_R input1763 (.A(io_ins_up_3[40]),
    .Y(net1763));
 BUFx2_ASAP7_75t_R input1764 (.A(io_ins_up_3[41]),
    .Y(net1764));
 BUFx2_ASAP7_75t_R input1765 (.A(io_ins_up_3[42]),
    .Y(net1765));
 BUFx2_ASAP7_75t_R input1766 (.A(io_ins_up_3[43]),
    .Y(net1766));
 BUFx2_ASAP7_75t_R input1767 (.A(io_ins_up_3[44]),
    .Y(net1767));
 BUFx2_ASAP7_75t_R input1768 (.A(io_ins_up_3[45]),
    .Y(net1768));
 BUFx2_ASAP7_75t_R input1769 (.A(io_ins_up_3[46]),
    .Y(net1769));
 BUFx2_ASAP7_75t_R input1770 (.A(io_ins_up_3[47]),
    .Y(net1770));
 BUFx2_ASAP7_75t_R input1771 (.A(io_ins_up_3[48]),
    .Y(net1771));
 BUFx2_ASAP7_75t_R input1772 (.A(io_ins_up_3[49]),
    .Y(net1772));
 BUFx2_ASAP7_75t_R input1773 (.A(io_ins_up_3[4]),
    .Y(net1773));
 BUFx2_ASAP7_75t_R input1774 (.A(io_ins_up_3[50]),
    .Y(net1774));
 BUFx2_ASAP7_75t_R input1775 (.A(io_ins_up_3[51]),
    .Y(net1775));
 BUFx2_ASAP7_75t_R input1776 (.A(io_ins_up_3[52]),
    .Y(net1776));
 BUFx2_ASAP7_75t_R input1777 (.A(io_ins_up_3[53]),
    .Y(net1777));
 BUFx2_ASAP7_75t_R input1778 (.A(io_ins_up_3[54]),
    .Y(net1778));
 BUFx2_ASAP7_75t_R input1779 (.A(io_ins_up_3[55]),
    .Y(net1779));
 BUFx2_ASAP7_75t_R input1780 (.A(io_ins_up_3[56]),
    .Y(net1780));
 BUFx2_ASAP7_75t_R input1781 (.A(io_ins_up_3[57]),
    .Y(net1781));
 BUFx2_ASAP7_75t_R input1782 (.A(io_ins_up_3[58]),
    .Y(net1782));
 BUFx2_ASAP7_75t_R input1783 (.A(io_ins_up_3[59]),
    .Y(net1783));
 BUFx2_ASAP7_75t_R input1784 (.A(io_ins_up_3[5]),
    .Y(net1784));
 BUFx2_ASAP7_75t_R input1785 (.A(io_ins_up_3[60]),
    .Y(net1785));
 BUFx2_ASAP7_75t_R input1786 (.A(io_ins_up_3[61]),
    .Y(net1786));
 BUFx2_ASAP7_75t_R input1787 (.A(io_ins_up_3[62]),
    .Y(net1787));
 BUFx2_ASAP7_75t_R input1788 (.A(io_ins_up_3[63]),
    .Y(net1788));
 BUFx2_ASAP7_75t_R input1789 (.A(io_ins_up_3[6]),
    .Y(net1789));
 BUFx2_ASAP7_75t_R input1790 (.A(io_ins_up_3[7]),
    .Y(net1790));
 BUFx2_ASAP7_75t_R input1791 (.A(io_ins_up_3[8]),
    .Y(net1791));
 BUFx2_ASAP7_75t_R input1792 (.A(io_ins_up_3[9]),
    .Y(net1792));
 BUFx2_ASAP7_75t_R input1793 (.A(io_ins_up_4[0]),
    .Y(net1793));
 BUFx2_ASAP7_75t_R input1794 (.A(io_ins_up_4[10]),
    .Y(net1794));
 BUFx2_ASAP7_75t_R input1795 (.A(io_ins_up_4[11]),
    .Y(net1795));
 BUFx2_ASAP7_75t_R input1796 (.A(io_ins_up_4[12]),
    .Y(net1796));
 BUFx2_ASAP7_75t_R input1797 (.A(io_ins_up_4[13]),
    .Y(net1797));
 BUFx2_ASAP7_75t_R input1798 (.A(io_ins_up_4[14]),
    .Y(net1798));
 BUFx2_ASAP7_75t_R input1799 (.A(io_ins_up_4[15]),
    .Y(net1799));
 BUFx2_ASAP7_75t_R input1800 (.A(io_ins_up_4[16]),
    .Y(net1800));
 BUFx2_ASAP7_75t_R input1801 (.A(io_ins_up_4[17]),
    .Y(net1801));
 BUFx2_ASAP7_75t_R input1802 (.A(io_ins_up_4[18]),
    .Y(net1802));
 BUFx2_ASAP7_75t_R input1803 (.A(io_ins_up_4[19]),
    .Y(net1803));
 BUFx2_ASAP7_75t_R input1804 (.A(io_ins_up_4[1]),
    .Y(net1804));
 BUFx2_ASAP7_75t_R input1805 (.A(io_ins_up_4[20]),
    .Y(net1805));
 BUFx2_ASAP7_75t_R input1806 (.A(io_ins_up_4[21]),
    .Y(net1806));
 BUFx2_ASAP7_75t_R input1807 (.A(io_ins_up_4[22]),
    .Y(net1807));
 BUFx2_ASAP7_75t_R input1808 (.A(io_ins_up_4[23]),
    .Y(net1808));
 BUFx2_ASAP7_75t_R input1809 (.A(io_ins_up_4[24]),
    .Y(net1809));
 BUFx2_ASAP7_75t_R input1810 (.A(io_ins_up_4[25]),
    .Y(net1810));
 BUFx2_ASAP7_75t_R input1811 (.A(io_ins_up_4[26]),
    .Y(net1811));
 BUFx2_ASAP7_75t_R input1812 (.A(io_ins_up_4[27]),
    .Y(net1812));
 BUFx2_ASAP7_75t_R input1813 (.A(io_ins_up_4[28]),
    .Y(net1813));
 BUFx2_ASAP7_75t_R input1814 (.A(io_ins_up_4[29]),
    .Y(net1814));
 BUFx2_ASAP7_75t_R input1815 (.A(io_ins_up_4[2]),
    .Y(net1815));
 BUFx2_ASAP7_75t_R input1816 (.A(io_ins_up_4[30]),
    .Y(net1816));
 BUFx2_ASAP7_75t_R input1817 (.A(io_ins_up_4[31]),
    .Y(net1817));
 BUFx2_ASAP7_75t_R input1818 (.A(io_ins_up_4[32]),
    .Y(net1818));
 BUFx2_ASAP7_75t_R input1819 (.A(io_ins_up_4[33]),
    .Y(net1819));
 BUFx2_ASAP7_75t_R input1820 (.A(io_ins_up_4[34]),
    .Y(net1820));
 BUFx2_ASAP7_75t_R input1821 (.A(io_ins_up_4[35]),
    .Y(net1821));
 BUFx2_ASAP7_75t_R input1822 (.A(io_ins_up_4[36]),
    .Y(net1822));
 BUFx2_ASAP7_75t_R input1823 (.A(io_ins_up_4[37]),
    .Y(net1823));
 BUFx2_ASAP7_75t_R input1824 (.A(io_ins_up_4[38]),
    .Y(net1824));
 BUFx2_ASAP7_75t_R input1825 (.A(io_ins_up_4[39]),
    .Y(net1825));
 BUFx2_ASAP7_75t_R input1826 (.A(io_ins_up_4[3]),
    .Y(net1826));
 BUFx2_ASAP7_75t_R input1827 (.A(io_ins_up_4[40]),
    .Y(net1827));
 BUFx2_ASAP7_75t_R input1828 (.A(io_ins_up_4[41]),
    .Y(net1828));
 BUFx2_ASAP7_75t_R input1829 (.A(io_ins_up_4[42]),
    .Y(net1829));
 BUFx2_ASAP7_75t_R input1830 (.A(io_ins_up_4[43]),
    .Y(net1830));
 BUFx2_ASAP7_75t_R input1831 (.A(io_ins_up_4[44]),
    .Y(net1831));
 BUFx2_ASAP7_75t_R input1832 (.A(io_ins_up_4[45]),
    .Y(net1832));
 BUFx2_ASAP7_75t_R input1833 (.A(io_ins_up_4[46]),
    .Y(net1833));
 BUFx2_ASAP7_75t_R input1834 (.A(io_ins_up_4[47]),
    .Y(net1834));
 BUFx2_ASAP7_75t_R input1835 (.A(io_ins_up_4[48]),
    .Y(net1835));
 BUFx2_ASAP7_75t_R input1836 (.A(io_ins_up_4[49]),
    .Y(net1836));
 BUFx2_ASAP7_75t_R input1837 (.A(io_ins_up_4[4]),
    .Y(net1837));
 BUFx2_ASAP7_75t_R input1838 (.A(io_ins_up_4[50]),
    .Y(net1838));
 BUFx2_ASAP7_75t_R input1839 (.A(io_ins_up_4[51]),
    .Y(net1839));
 BUFx2_ASAP7_75t_R input1840 (.A(io_ins_up_4[52]),
    .Y(net1840));
 BUFx2_ASAP7_75t_R input1841 (.A(io_ins_up_4[53]),
    .Y(net1841));
 BUFx2_ASAP7_75t_R input1842 (.A(io_ins_up_4[54]),
    .Y(net1842));
 BUFx2_ASAP7_75t_R input1843 (.A(io_ins_up_4[55]),
    .Y(net1843));
 BUFx2_ASAP7_75t_R input1844 (.A(io_ins_up_4[56]),
    .Y(net1844));
 BUFx2_ASAP7_75t_R input1845 (.A(io_ins_up_4[57]),
    .Y(net1845));
 BUFx2_ASAP7_75t_R input1846 (.A(io_ins_up_4[58]),
    .Y(net1846));
 BUFx2_ASAP7_75t_R input1847 (.A(io_ins_up_4[59]),
    .Y(net1847));
 BUFx2_ASAP7_75t_R input1848 (.A(io_ins_up_4[5]),
    .Y(net1848));
 BUFx2_ASAP7_75t_R input1849 (.A(io_ins_up_4[60]),
    .Y(net1849));
 BUFx2_ASAP7_75t_R input1850 (.A(io_ins_up_4[61]),
    .Y(net1850));
 BUFx2_ASAP7_75t_R input1851 (.A(io_ins_up_4[62]),
    .Y(net1851));
 BUFx2_ASAP7_75t_R input1852 (.A(io_ins_up_4[63]),
    .Y(net1852));
 BUFx2_ASAP7_75t_R input1853 (.A(io_ins_up_4[6]),
    .Y(net1853));
 BUFx2_ASAP7_75t_R input1854 (.A(io_ins_up_4[7]),
    .Y(net1854));
 BUFx2_ASAP7_75t_R input1855 (.A(io_ins_up_4[8]),
    .Y(net1855));
 BUFx2_ASAP7_75t_R input1856 (.A(io_ins_up_4[9]),
    .Y(net1856));
 BUFx2_ASAP7_75t_R input1857 (.A(io_ins_up_5[0]),
    .Y(net1857));
 BUFx2_ASAP7_75t_R input1858 (.A(io_ins_up_5[10]),
    .Y(net1858));
 BUFx2_ASAP7_75t_R input1859 (.A(io_ins_up_5[11]),
    .Y(net1859));
 BUFx2_ASAP7_75t_R input1860 (.A(io_ins_up_5[12]),
    .Y(net1860));
 BUFx2_ASAP7_75t_R input1861 (.A(io_ins_up_5[13]),
    .Y(net1861));
 BUFx2_ASAP7_75t_R input1862 (.A(io_ins_up_5[14]),
    .Y(net1862));
 BUFx2_ASAP7_75t_R input1863 (.A(io_ins_up_5[15]),
    .Y(net1863));
 BUFx2_ASAP7_75t_R input1864 (.A(io_ins_up_5[16]),
    .Y(net1864));
 BUFx2_ASAP7_75t_R input1865 (.A(io_ins_up_5[17]),
    .Y(net1865));
 BUFx2_ASAP7_75t_R input1866 (.A(io_ins_up_5[18]),
    .Y(net1866));
 BUFx2_ASAP7_75t_R input1867 (.A(io_ins_up_5[19]),
    .Y(net1867));
 BUFx2_ASAP7_75t_R input1868 (.A(io_ins_up_5[1]),
    .Y(net1868));
 BUFx2_ASAP7_75t_R input1869 (.A(io_ins_up_5[20]),
    .Y(net1869));
 BUFx2_ASAP7_75t_R input1870 (.A(io_ins_up_5[21]),
    .Y(net1870));
 BUFx2_ASAP7_75t_R input1871 (.A(io_ins_up_5[22]),
    .Y(net1871));
 BUFx2_ASAP7_75t_R input1872 (.A(io_ins_up_5[23]),
    .Y(net1872));
 BUFx2_ASAP7_75t_R input1873 (.A(io_ins_up_5[24]),
    .Y(net1873));
 BUFx2_ASAP7_75t_R input1874 (.A(io_ins_up_5[25]),
    .Y(net1874));
 BUFx2_ASAP7_75t_R input1875 (.A(io_ins_up_5[26]),
    .Y(net1875));
 BUFx2_ASAP7_75t_R input1876 (.A(io_ins_up_5[27]),
    .Y(net1876));
 BUFx2_ASAP7_75t_R input1877 (.A(io_ins_up_5[28]),
    .Y(net1877));
 BUFx2_ASAP7_75t_R input1878 (.A(io_ins_up_5[29]),
    .Y(net1878));
 BUFx2_ASAP7_75t_R input1879 (.A(io_ins_up_5[2]),
    .Y(net1879));
 BUFx2_ASAP7_75t_R input1880 (.A(io_ins_up_5[30]),
    .Y(net1880));
 BUFx2_ASAP7_75t_R input1881 (.A(io_ins_up_5[31]),
    .Y(net1881));
 BUFx2_ASAP7_75t_R input1882 (.A(io_ins_up_5[32]),
    .Y(net1882));
 BUFx2_ASAP7_75t_R input1883 (.A(io_ins_up_5[33]),
    .Y(net1883));
 BUFx2_ASAP7_75t_R input1884 (.A(io_ins_up_5[34]),
    .Y(net1884));
 BUFx2_ASAP7_75t_R input1885 (.A(io_ins_up_5[35]),
    .Y(net1885));
 BUFx2_ASAP7_75t_R input1886 (.A(io_ins_up_5[36]),
    .Y(net1886));
 BUFx2_ASAP7_75t_R input1887 (.A(io_ins_up_5[37]),
    .Y(net1887));
 BUFx2_ASAP7_75t_R input1888 (.A(io_ins_up_5[38]),
    .Y(net1888));
 BUFx2_ASAP7_75t_R input1889 (.A(io_ins_up_5[39]),
    .Y(net1889));
 BUFx2_ASAP7_75t_R input1890 (.A(io_ins_up_5[3]),
    .Y(net1890));
 BUFx2_ASAP7_75t_R input1891 (.A(io_ins_up_5[40]),
    .Y(net1891));
 BUFx2_ASAP7_75t_R input1892 (.A(io_ins_up_5[41]),
    .Y(net1892));
 BUFx2_ASAP7_75t_R input1893 (.A(io_ins_up_5[42]),
    .Y(net1893));
 BUFx2_ASAP7_75t_R input1894 (.A(io_ins_up_5[43]),
    .Y(net1894));
 BUFx2_ASAP7_75t_R input1895 (.A(io_ins_up_5[44]),
    .Y(net1895));
 BUFx2_ASAP7_75t_R input1896 (.A(io_ins_up_5[45]),
    .Y(net1896));
 BUFx2_ASAP7_75t_R input1897 (.A(io_ins_up_5[46]),
    .Y(net1897));
 BUFx2_ASAP7_75t_R input1898 (.A(io_ins_up_5[47]),
    .Y(net1898));
 BUFx2_ASAP7_75t_R input1899 (.A(io_ins_up_5[48]),
    .Y(net1899));
 BUFx2_ASAP7_75t_R input1900 (.A(io_ins_up_5[49]),
    .Y(net1900));
 BUFx2_ASAP7_75t_R input1901 (.A(io_ins_up_5[4]),
    .Y(net1901));
 BUFx2_ASAP7_75t_R input1902 (.A(io_ins_up_5[50]),
    .Y(net1902));
 BUFx2_ASAP7_75t_R input1903 (.A(io_ins_up_5[51]),
    .Y(net1903));
 BUFx2_ASAP7_75t_R input1904 (.A(io_ins_up_5[52]),
    .Y(net1904));
 BUFx2_ASAP7_75t_R input1905 (.A(io_ins_up_5[53]),
    .Y(net1905));
 BUFx2_ASAP7_75t_R input1906 (.A(io_ins_up_5[54]),
    .Y(net1906));
 BUFx2_ASAP7_75t_R input1907 (.A(io_ins_up_5[55]),
    .Y(net1907));
 BUFx2_ASAP7_75t_R input1908 (.A(io_ins_up_5[56]),
    .Y(net1908));
 BUFx2_ASAP7_75t_R input1909 (.A(io_ins_up_5[57]),
    .Y(net1909));
 BUFx2_ASAP7_75t_R input1910 (.A(io_ins_up_5[58]),
    .Y(net1910));
 BUFx2_ASAP7_75t_R input1911 (.A(io_ins_up_5[59]),
    .Y(net1911));
 BUFx2_ASAP7_75t_R input1912 (.A(io_ins_up_5[5]),
    .Y(net1912));
 BUFx2_ASAP7_75t_R input1913 (.A(io_ins_up_5[60]),
    .Y(net1913));
 BUFx2_ASAP7_75t_R input1914 (.A(io_ins_up_5[61]),
    .Y(net1914));
 BUFx2_ASAP7_75t_R input1915 (.A(io_ins_up_5[62]),
    .Y(net1915));
 BUFx2_ASAP7_75t_R input1916 (.A(io_ins_up_5[63]),
    .Y(net1916));
 BUFx2_ASAP7_75t_R input1917 (.A(io_ins_up_5[6]),
    .Y(net1917));
 BUFx2_ASAP7_75t_R input1918 (.A(io_ins_up_5[7]),
    .Y(net1918));
 BUFx2_ASAP7_75t_R input1919 (.A(io_ins_up_5[8]),
    .Y(net1919));
 BUFx2_ASAP7_75t_R input1920 (.A(io_ins_up_5[9]),
    .Y(net1920));
 BUFx2_ASAP7_75t_R input1921 (.A(io_ins_up_6[0]),
    .Y(net1921));
 BUFx2_ASAP7_75t_R input1922 (.A(io_ins_up_6[10]),
    .Y(net1922));
 BUFx2_ASAP7_75t_R input1923 (.A(io_ins_up_6[11]),
    .Y(net1923));
 BUFx2_ASAP7_75t_R input1924 (.A(io_ins_up_6[12]),
    .Y(net1924));
 BUFx2_ASAP7_75t_R input1925 (.A(io_ins_up_6[13]),
    .Y(net1925));
 BUFx2_ASAP7_75t_R input1926 (.A(io_ins_up_6[14]),
    .Y(net1926));
 BUFx2_ASAP7_75t_R input1927 (.A(io_ins_up_6[15]),
    .Y(net1927));
 BUFx2_ASAP7_75t_R input1928 (.A(io_ins_up_6[16]),
    .Y(net1928));
 BUFx2_ASAP7_75t_R input1929 (.A(io_ins_up_6[17]),
    .Y(net1929));
 BUFx2_ASAP7_75t_R input1930 (.A(io_ins_up_6[18]),
    .Y(net1930));
 BUFx2_ASAP7_75t_R input1931 (.A(io_ins_up_6[19]),
    .Y(net1931));
 BUFx2_ASAP7_75t_R input1932 (.A(io_ins_up_6[1]),
    .Y(net1932));
 BUFx2_ASAP7_75t_R input1933 (.A(io_ins_up_6[20]),
    .Y(net1933));
 BUFx2_ASAP7_75t_R input1934 (.A(io_ins_up_6[21]),
    .Y(net1934));
 BUFx2_ASAP7_75t_R input1935 (.A(io_ins_up_6[22]),
    .Y(net1935));
 BUFx2_ASAP7_75t_R input1936 (.A(io_ins_up_6[23]),
    .Y(net1936));
 BUFx2_ASAP7_75t_R input1937 (.A(io_ins_up_6[24]),
    .Y(net1937));
 BUFx2_ASAP7_75t_R input1938 (.A(io_ins_up_6[25]),
    .Y(net1938));
 BUFx2_ASAP7_75t_R input1939 (.A(io_ins_up_6[26]),
    .Y(net1939));
 BUFx2_ASAP7_75t_R input1940 (.A(io_ins_up_6[27]),
    .Y(net1940));
 BUFx2_ASAP7_75t_R input1941 (.A(io_ins_up_6[28]),
    .Y(net1941));
 BUFx2_ASAP7_75t_R input1942 (.A(io_ins_up_6[29]),
    .Y(net1942));
 BUFx2_ASAP7_75t_R input1943 (.A(io_ins_up_6[2]),
    .Y(net1943));
 BUFx2_ASAP7_75t_R input1944 (.A(io_ins_up_6[30]),
    .Y(net1944));
 BUFx2_ASAP7_75t_R input1945 (.A(io_ins_up_6[31]),
    .Y(net1945));
 BUFx2_ASAP7_75t_R input1946 (.A(io_ins_up_6[32]),
    .Y(net1946));
 BUFx2_ASAP7_75t_R input1947 (.A(io_ins_up_6[33]),
    .Y(net1947));
 BUFx2_ASAP7_75t_R input1948 (.A(io_ins_up_6[34]),
    .Y(net1948));
 BUFx2_ASAP7_75t_R input1949 (.A(io_ins_up_6[35]),
    .Y(net1949));
 BUFx2_ASAP7_75t_R input1950 (.A(io_ins_up_6[36]),
    .Y(net1950));
 BUFx2_ASAP7_75t_R input1951 (.A(io_ins_up_6[37]),
    .Y(net1951));
 BUFx2_ASAP7_75t_R input1952 (.A(io_ins_up_6[38]),
    .Y(net1952));
 BUFx2_ASAP7_75t_R input1953 (.A(io_ins_up_6[39]),
    .Y(net1953));
 BUFx2_ASAP7_75t_R input1954 (.A(io_ins_up_6[3]),
    .Y(net1954));
 BUFx2_ASAP7_75t_R input1955 (.A(io_ins_up_6[40]),
    .Y(net1955));
 BUFx2_ASAP7_75t_R input1956 (.A(io_ins_up_6[41]),
    .Y(net1956));
 BUFx2_ASAP7_75t_R input1957 (.A(io_ins_up_6[42]),
    .Y(net1957));
 BUFx2_ASAP7_75t_R input1958 (.A(io_ins_up_6[43]),
    .Y(net1958));
 BUFx2_ASAP7_75t_R input1959 (.A(io_ins_up_6[44]),
    .Y(net1959));
 BUFx2_ASAP7_75t_R input1960 (.A(io_ins_up_6[45]),
    .Y(net1960));
 BUFx2_ASAP7_75t_R input1961 (.A(io_ins_up_6[46]),
    .Y(net1961));
 BUFx2_ASAP7_75t_R input1962 (.A(io_ins_up_6[47]),
    .Y(net1962));
 BUFx2_ASAP7_75t_R input1963 (.A(io_ins_up_6[48]),
    .Y(net1963));
 BUFx2_ASAP7_75t_R input1964 (.A(io_ins_up_6[49]),
    .Y(net1964));
 BUFx2_ASAP7_75t_R input1965 (.A(io_ins_up_6[4]),
    .Y(net1965));
 BUFx2_ASAP7_75t_R input1966 (.A(io_ins_up_6[50]),
    .Y(net1966));
 BUFx2_ASAP7_75t_R input1967 (.A(io_ins_up_6[51]),
    .Y(net1967));
 BUFx2_ASAP7_75t_R input1968 (.A(io_ins_up_6[52]),
    .Y(net1968));
 BUFx2_ASAP7_75t_R input1969 (.A(io_ins_up_6[53]),
    .Y(net1969));
 BUFx2_ASAP7_75t_R input1970 (.A(io_ins_up_6[54]),
    .Y(net1970));
 BUFx2_ASAP7_75t_R input1971 (.A(io_ins_up_6[55]),
    .Y(net1971));
 BUFx2_ASAP7_75t_R input1972 (.A(io_ins_up_6[56]),
    .Y(net1972));
 BUFx2_ASAP7_75t_R input1973 (.A(io_ins_up_6[57]),
    .Y(net1973));
 BUFx2_ASAP7_75t_R input1974 (.A(io_ins_up_6[58]),
    .Y(net1974));
 BUFx2_ASAP7_75t_R input1975 (.A(io_ins_up_6[59]),
    .Y(net1975));
 BUFx2_ASAP7_75t_R input1976 (.A(io_ins_up_6[5]),
    .Y(net1976));
 BUFx2_ASAP7_75t_R input1977 (.A(io_ins_up_6[60]),
    .Y(net1977));
 BUFx2_ASAP7_75t_R input1978 (.A(io_ins_up_6[61]),
    .Y(net1978));
 BUFx2_ASAP7_75t_R input1979 (.A(io_ins_up_6[62]),
    .Y(net1979));
 BUFx2_ASAP7_75t_R input1980 (.A(io_ins_up_6[63]),
    .Y(net1980));
 BUFx2_ASAP7_75t_R input1981 (.A(io_ins_up_6[6]),
    .Y(net1981));
 BUFx2_ASAP7_75t_R input1982 (.A(io_ins_up_6[7]),
    .Y(net1982));
 BUFx2_ASAP7_75t_R input1983 (.A(io_ins_up_6[8]),
    .Y(net1983));
 BUFx2_ASAP7_75t_R input1984 (.A(io_ins_up_6[9]),
    .Y(net1984));
 BUFx2_ASAP7_75t_R input1985 (.A(io_ins_up_7[0]),
    .Y(net1985));
 BUFx2_ASAP7_75t_R input1986 (.A(io_ins_up_7[10]),
    .Y(net1986));
 BUFx2_ASAP7_75t_R input1987 (.A(io_ins_up_7[11]),
    .Y(net1987));
 BUFx2_ASAP7_75t_R input1988 (.A(io_ins_up_7[12]),
    .Y(net1988));
 BUFx2_ASAP7_75t_R input1989 (.A(io_ins_up_7[13]),
    .Y(net1989));
 BUFx2_ASAP7_75t_R input1990 (.A(io_ins_up_7[14]),
    .Y(net1990));
 BUFx2_ASAP7_75t_R input1991 (.A(io_ins_up_7[15]),
    .Y(net1991));
 BUFx2_ASAP7_75t_R input1992 (.A(io_ins_up_7[16]),
    .Y(net1992));
 BUFx2_ASAP7_75t_R input1993 (.A(io_ins_up_7[17]),
    .Y(net1993));
 BUFx2_ASAP7_75t_R input1994 (.A(io_ins_up_7[18]),
    .Y(net1994));
 BUFx2_ASAP7_75t_R input1995 (.A(io_ins_up_7[19]),
    .Y(net1995));
 BUFx2_ASAP7_75t_R input1996 (.A(io_ins_up_7[1]),
    .Y(net1996));
 BUFx2_ASAP7_75t_R input1997 (.A(io_ins_up_7[20]),
    .Y(net1997));
 BUFx2_ASAP7_75t_R input1998 (.A(io_ins_up_7[21]),
    .Y(net1998));
 BUFx2_ASAP7_75t_R input1999 (.A(io_ins_up_7[22]),
    .Y(net1999));
 BUFx2_ASAP7_75t_R input2000 (.A(io_ins_up_7[23]),
    .Y(net2000));
 BUFx2_ASAP7_75t_R input2001 (.A(io_ins_up_7[24]),
    .Y(net2001));
 BUFx2_ASAP7_75t_R input2002 (.A(io_ins_up_7[25]),
    .Y(net2002));
 BUFx2_ASAP7_75t_R input2003 (.A(io_ins_up_7[26]),
    .Y(net2003));
 BUFx2_ASAP7_75t_R input2004 (.A(io_ins_up_7[27]),
    .Y(net2004));
 BUFx2_ASAP7_75t_R input2005 (.A(io_ins_up_7[28]),
    .Y(net2005));
 BUFx2_ASAP7_75t_R input2006 (.A(io_ins_up_7[29]),
    .Y(net2006));
 BUFx2_ASAP7_75t_R input2007 (.A(io_ins_up_7[2]),
    .Y(net2007));
 BUFx2_ASAP7_75t_R input2008 (.A(io_ins_up_7[30]),
    .Y(net2008));
 BUFx2_ASAP7_75t_R input2009 (.A(io_ins_up_7[31]),
    .Y(net2009));
 BUFx2_ASAP7_75t_R input2010 (.A(io_ins_up_7[32]),
    .Y(net2010));
 BUFx2_ASAP7_75t_R input2011 (.A(io_ins_up_7[33]),
    .Y(net2011));
 BUFx2_ASAP7_75t_R input2012 (.A(io_ins_up_7[34]),
    .Y(net2012));
 BUFx2_ASAP7_75t_R input2013 (.A(io_ins_up_7[35]),
    .Y(net2013));
 BUFx2_ASAP7_75t_R input2014 (.A(io_ins_up_7[36]),
    .Y(net2014));
 BUFx2_ASAP7_75t_R input2015 (.A(io_ins_up_7[37]),
    .Y(net2015));
 BUFx2_ASAP7_75t_R input2016 (.A(io_ins_up_7[38]),
    .Y(net2016));
 BUFx2_ASAP7_75t_R input2017 (.A(io_ins_up_7[39]),
    .Y(net2017));
 BUFx2_ASAP7_75t_R input2018 (.A(io_ins_up_7[3]),
    .Y(net2018));
 BUFx2_ASAP7_75t_R input2019 (.A(io_ins_up_7[40]),
    .Y(net2019));
 BUFx2_ASAP7_75t_R input2020 (.A(io_ins_up_7[41]),
    .Y(net2020));
 BUFx2_ASAP7_75t_R input2021 (.A(io_ins_up_7[42]),
    .Y(net2021));
 BUFx2_ASAP7_75t_R input2022 (.A(io_ins_up_7[43]),
    .Y(net2022));
 BUFx2_ASAP7_75t_R input2023 (.A(io_ins_up_7[44]),
    .Y(net2023));
 BUFx2_ASAP7_75t_R input2024 (.A(io_ins_up_7[45]),
    .Y(net2024));
 BUFx2_ASAP7_75t_R input2025 (.A(io_ins_up_7[46]),
    .Y(net2025));
 BUFx2_ASAP7_75t_R input2026 (.A(io_ins_up_7[47]),
    .Y(net2026));
 BUFx2_ASAP7_75t_R input2027 (.A(io_ins_up_7[48]),
    .Y(net2027));
 BUFx2_ASAP7_75t_R input2028 (.A(io_ins_up_7[49]),
    .Y(net2028));
 BUFx2_ASAP7_75t_R input2029 (.A(io_ins_up_7[4]),
    .Y(net2029));
 BUFx2_ASAP7_75t_R input2030 (.A(io_ins_up_7[50]),
    .Y(net2030));
 BUFx2_ASAP7_75t_R input2031 (.A(io_ins_up_7[51]),
    .Y(net2031));
 BUFx2_ASAP7_75t_R input2032 (.A(io_ins_up_7[52]),
    .Y(net2032));
 BUFx2_ASAP7_75t_R input2033 (.A(io_ins_up_7[53]),
    .Y(net2033));
 BUFx2_ASAP7_75t_R input2034 (.A(io_ins_up_7[54]),
    .Y(net2034));
 BUFx2_ASAP7_75t_R input2035 (.A(io_ins_up_7[55]),
    .Y(net2035));
 BUFx2_ASAP7_75t_R input2036 (.A(io_ins_up_7[56]),
    .Y(net2036));
 BUFx2_ASAP7_75t_R input2037 (.A(io_ins_up_7[57]),
    .Y(net2037));
 BUFx2_ASAP7_75t_R input2038 (.A(io_ins_up_7[58]),
    .Y(net2038));
 BUFx2_ASAP7_75t_R input2039 (.A(io_ins_up_7[59]),
    .Y(net2039));
 BUFx2_ASAP7_75t_R input2040 (.A(io_ins_up_7[5]),
    .Y(net2040));
 BUFx2_ASAP7_75t_R input2041 (.A(io_ins_up_7[60]),
    .Y(net2041));
 BUFx2_ASAP7_75t_R input2042 (.A(io_ins_up_7[61]),
    .Y(net2042));
 BUFx2_ASAP7_75t_R input2043 (.A(io_ins_up_7[62]),
    .Y(net2043));
 BUFx2_ASAP7_75t_R input2044 (.A(io_ins_up_7[63]),
    .Y(net2044));
 BUFx2_ASAP7_75t_R input2045 (.A(io_ins_up_7[6]),
    .Y(net2045));
 BUFx2_ASAP7_75t_R input2046 (.A(io_ins_up_7[7]),
    .Y(net2046));
 BUFx2_ASAP7_75t_R input2047 (.A(io_ins_up_7[8]),
    .Y(net2047));
 BUFx2_ASAP7_75t_R input2048 (.A(io_ins_up_7[9]),
    .Y(net2048));
 BUFx2_ASAP7_75t_R output2049 (.A(net2049),
    .Y(io_lsbs_0));
 BUFx2_ASAP7_75t_R output2050 (.A(net2050),
    .Y(io_lsbs_1));
 BUFx2_ASAP7_75t_R output2051 (.A(net2051),
    .Y(io_lsbs_10));
 BUFx2_ASAP7_75t_R output2052 (.A(net2052),
    .Y(io_lsbs_11));
 BUFx2_ASAP7_75t_R output2053 (.A(net2053),
    .Y(io_lsbs_12));
 BUFx2_ASAP7_75t_R output2054 (.A(net2054),
    .Y(io_lsbs_13));
 BUFx2_ASAP7_75t_R output2055 (.A(net2055),
    .Y(io_lsbs_14));
 BUFx2_ASAP7_75t_R output2056 (.A(net2056),
    .Y(io_lsbs_15));
 BUFx2_ASAP7_75t_R output2057 (.A(net2057),
    .Y(io_lsbs_16));
 BUFx2_ASAP7_75t_R output2058 (.A(net2058),
    .Y(io_lsbs_17));
 BUFx2_ASAP7_75t_R output2059 (.A(net2059),
    .Y(io_lsbs_18));
 BUFx2_ASAP7_75t_R output2060 (.A(net2060),
    .Y(io_lsbs_19));
 BUFx2_ASAP7_75t_R output2061 (.A(net2061),
    .Y(io_lsbs_2));
 BUFx2_ASAP7_75t_R output2062 (.A(net2062),
    .Y(io_lsbs_20));
 BUFx2_ASAP7_75t_R output2063 (.A(net2063),
    .Y(io_lsbs_21));
 BUFx2_ASAP7_75t_R output2064 (.A(net2064),
    .Y(io_lsbs_22));
 BUFx2_ASAP7_75t_R output2065 (.A(net2065),
    .Y(io_lsbs_23));
 BUFx2_ASAP7_75t_R output2066 (.A(net2066),
    .Y(io_lsbs_24));
 BUFx2_ASAP7_75t_R output2067 (.A(net2067),
    .Y(io_lsbs_25));
 BUFx2_ASAP7_75t_R output2068 (.A(net2068),
    .Y(io_lsbs_26));
 BUFx2_ASAP7_75t_R output2069 (.A(net2069),
    .Y(io_lsbs_27));
 BUFx2_ASAP7_75t_R output2070 (.A(net2070),
    .Y(io_lsbs_28));
 BUFx2_ASAP7_75t_R output2071 (.A(net2071),
    .Y(io_lsbs_29));
 BUFx2_ASAP7_75t_R output2072 (.A(net2072),
    .Y(io_lsbs_3));
 BUFx2_ASAP7_75t_R output2073 (.A(net2073),
    .Y(io_lsbs_30));
 BUFx2_ASAP7_75t_R output2074 (.A(net2074),
    .Y(io_lsbs_31));
 BUFx2_ASAP7_75t_R output2075 (.A(net2075),
    .Y(io_lsbs_32));
 BUFx2_ASAP7_75t_R output2076 (.A(net2076),
    .Y(io_lsbs_33));
 BUFx2_ASAP7_75t_R output2077 (.A(net2077),
    .Y(io_lsbs_34));
 BUFx2_ASAP7_75t_R output2078 (.A(net2078),
    .Y(io_lsbs_35));
 BUFx2_ASAP7_75t_R output2079 (.A(net2079),
    .Y(io_lsbs_36));
 BUFx2_ASAP7_75t_R output2080 (.A(net2080),
    .Y(io_lsbs_37));
 BUFx2_ASAP7_75t_R output2081 (.A(net2081),
    .Y(io_lsbs_38));
 BUFx2_ASAP7_75t_R output2082 (.A(net2082),
    .Y(io_lsbs_39));
 BUFx2_ASAP7_75t_R output2083 (.A(net2083),
    .Y(io_lsbs_4));
 BUFx2_ASAP7_75t_R output2084 (.A(net2084),
    .Y(io_lsbs_40));
 BUFx2_ASAP7_75t_R output2085 (.A(net2085),
    .Y(io_lsbs_41));
 BUFx2_ASAP7_75t_R output2086 (.A(net2086),
    .Y(io_lsbs_42));
 BUFx2_ASAP7_75t_R output2087 (.A(net2087),
    .Y(io_lsbs_43));
 BUFx2_ASAP7_75t_R output2088 (.A(net2088),
    .Y(io_lsbs_44));
 BUFx2_ASAP7_75t_R output2089 (.A(net2089),
    .Y(io_lsbs_45));
 BUFx2_ASAP7_75t_R output2090 (.A(net2090),
    .Y(io_lsbs_46));
 BUFx2_ASAP7_75t_R output2091 (.A(net2091),
    .Y(io_lsbs_47));
 BUFx2_ASAP7_75t_R output2092 (.A(net2092),
    .Y(io_lsbs_48));
 BUFx2_ASAP7_75t_R output2093 (.A(net2093),
    .Y(io_lsbs_49));
 BUFx2_ASAP7_75t_R output2094 (.A(net2094),
    .Y(io_lsbs_5));
 BUFx2_ASAP7_75t_R output2095 (.A(net2095),
    .Y(io_lsbs_50));
 BUFx2_ASAP7_75t_R output2096 (.A(net2096),
    .Y(io_lsbs_51));
 BUFx2_ASAP7_75t_R output2097 (.A(net2097),
    .Y(io_lsbs_52));
 BUFx2_ASAP7_75t_R output2098 (.A(net2098),
    .Y(io_lsbs_53));
 BUFx2_ASAP7_75t_R output2099 (.A(net2099),
    .Y(io_lsbs_54));
 BUFx2_ASAP7_75t_R output2100 (.A(net2100),
    .Y(io_lsbs_55));
 BUFx2_ASAP7_75t_R output2101 (.A(net2101),
    .Y(io_lsbs_56));
 BUFx2_ASAP7_75t_R output2102 (.A(net2102),
    .Y(io_lsbs_57));
 BUFx2_ASAP7_75t_R output2103 (.A(net2103),
    .Y(io_lsbs_58));
 BUFx2_ASAP7_75t_R output2104 (.A(net2104),
    .Y(io_lsbs_59));
 BUFx2_ASAP7_75t_R output2105 (.A(net2105),
    .Y(io_lsbs_6));
 BUFx2_ASAP7_75t_R output2106 (.A(net2106),
    .Y(io_lsbs_60));
 BUFx2_ASAP7_75t_R output2107 (.A(net2107),
    .Y(io_lsbs_61));
 BUFx2_ASAP7_75t_R output2108 (.A(net2108),
    .Y(io_lsbs_62));
 BUFx2_ASAP7_75t_R output2109 (.A(net2109),
    .Y(io_lsbs_63));
 BUFx2_ASAP7_75t_R output2110 (.A(net2110),
    .Y(io_lsbs_7));
 BUFx2_ASAP7_75t_R output2111 (.A(net2111),
    .Y(io_lsbs_8));
 BUFx2_ASAP7_75t_R output2112 (.A(net2112),
    .Y(io_lsbs_9));
 BUFx2_ASAP7_75t_R output2113 (.A(net2113),
    .Y(io_outs_down_0[0]));
 BUFx2_ASAP7_75t_R output2114 (.A(net2114),
    .Y(io_outs_down_0[10]));
 BUFx2_ASAP7_75t_R output2115 (.A(net2115),
    .Y(io_outs_down_0[11]));
 BUFx2_ASAP7_75t_R output2116 (.A(net2116),
    .Y(io_outs_down_0[12]));
 BUFx2_ASAP7_75t_R output2117 (.A(net2117),
    .Y(io_outs_down_0[13]));
 BUFx2_ASAP7_75t_R output2118 (.A(net2118),
    .Y(io_outs_down_0[14]));
 BUFx2_ASAP7_75t_R output2119 (.A(net2119),
    .Y(io_outs_down_0[15]));
 BUFx2_ASAP7_75t_R output2120 (.A(net2120),
    .Y(io_outs_down_0[16]));
 BUFx2_ASAP7_75t_R output2121 (.A(net2121),
    .Y(io_outs_down_0[17]));
 BUFx2_ASAP7_75t_R output2122 (.A(net2122),
    .Y(io_outs_down_0[18]));
 BUFx2_ASAP7_75t_R output2123 (.A(net2123),
    .Y(io_outs_down_0[19]));
 BUFx2_ASAP7_75t_R output2124 (.A(net2124),
    .Y(io_outs_down_0[1]));
 BUFx2_ASAP7_75t_R output2125 (.A(net2125),
    .Y(io_outs_down_0[20]));
 BUFx2_ASAP7_75t_R output2126 (.A(net2126),
    .Y(io_outs_down_0[21]));
 BUFx2_ASAP7_75t_R output2127 (.A(net2127),
    .Y(io_outs_down_0[22]));
 BUFx2_ASAP7_75t_R output2128 (.A(net2128),
    .Y(io_outs_down_0[23]));
 BUFx2_ASAP7_75t_R output2129 (.A(net2129),
    .Y(io_outs_down_0[24]));
 BUFx2_ASAP7_75t_R output2130 (.A(net2130),
    .Y(io_outs_down_0[25]));
 BUFx2_ASAP7_75t_R output2131 (.A(net2131),
    .Y(io_outs_down_0[26]));
 BUFx2_ASAP7_75t_R output2132 (.A(net2132),
    .Y(io_outs_down_0[27]));
 BUFx2_ASAP7_75t_R output2133 (.A(net2133),
    .Y(io_outs_down_0[28]));
 BUFx2_ASAP7_75t_R output2134 (.A(net2134),
    .Y(io_outs_down_0[29]));
 BUFx2_ASAP7_75t_R output2135 (.A(net2135),
    .Y(io_outs_down_0[2]));
 BUFx2_ASAP7_75t_R output2136 (.A(net2136),
    .Y(io_outs_down_0[30]));
 BUFx2_ASAP7_75t_R output2137 (.A(net2137),
    .Y(io_outs_down_0[31]));
 BUFx2_ASAP7_75t_R output2138 (.A(net2138),
    .Y(io_outs_down_0[32]));
 BUFx2_ASAP7_75t_R output2139 (.A(net2139),
    .Y(io_outs_down_0[33]));
 BUFx2_ASAP7_75t_R output2140 (.A(net2140),
    .Y(io_outs_down_0[34]));
 BUFx2_ASAP7_75t_R output2141 (.A(net2141),
    .Y(io_outs_down_0[35]));
 BUFx2_ASAP7_75t_R output2142 (.A(net2142),
    .Y(io_outs_down_0[36]));
 BUFx2_ASAP7_75t_R output2143 (.A(net2143),
    .Y(io_outs_down_0[37]));
 BUFx2_ASAP7_75t_R output2144 (.A(net2144),
    .Y(io_outs_down_0[38]));
 BUFx2_ASAP7_75t_R output2145 (.A(net2145),
    .Y(io_outs_down_0[39]));
 BUFx2_ASAP7_75t_R output2146 (.A(net2146),
    .Y(io_outs_down_0[3]));
 BUFx2_ASAP7_75t_R output2147 (.A(net2147),
    .Y(io_outs_down_0[40]));
 BUFx2_ASAP7_75t_R output2148 (.A(net2148),
    .Y(io_outs_down_0[41]));
 BUFx2_ASAP7_75t_R output2149 (.A(net2149),
    .Y(io_outs_down_0[42]));
 BUFx2_ASAP7_75t_R output2150 (.A(net2150),
    .Y(io_outs_down_0[43]));
 BUFx2_ASAP7_75t_R output2151 (.A(net2151),
    .Y(io_outs_down_0[44]));
 BUFx2_ASAP7_75t_R output2152 (.A(net2152),
    .Y(io_outs_down_0[45]));
 BUFx2_ASAP7_75t_R output2153 (.A(net2153),
    .Y(io_outs_down_0[46]));
 BUFx2_ASAP7_75t_R output2154 (.A(net2154),
    .Y(io_outs_down_0[47]));
 BUFx2_ASAP7_75t_R output2155 (.A(net2155),
    .Y(io_outs_down_0[48]));
 BUFx2_ASAP7_75t_R output2156 (.A(net2156),
    .Y(io_outs_down_0[49]));
 BUFx2_ASAP7_75t_R output2157 (.A(net2157),
    .Y(io_outs_down_0[4]));
 BUFx2_ASAP7_75t_R output2158 (.A(net2158),
    .Y(io_outs_down_0[50]));
 BUFx2_ASAP7_75t_R output2159 (.A(net2159),
    .Y(io_outs_down_0[51]));
 BUFx2_ASAP7_75t_R output2160 (.A(net2160),
    .Y(io_outs_down_0[52]));
 BUFx2_ASAP7_75t_R output2161 (.A(net2161),
    .Y(io_outs_down_0[53]));
 BUFx2_ASAP7_75t_R output2162 (.A(net2162),
    .Y(io_outs_down_0[54]));
 BUFx2_ASAP7_75t_R output2163 (.A(net2163),
    .Y(io_outs_down_0[55]));
 BUFx2_ASAP7_75t_R output2164 (.A(net2164),
    .Y(io_outs_down_0[56]));
 BUFx2_ASAP7_75t_R output2165 (.A(net2165),
    .Y(io_outs_down_0[57]));
 BUFx2_ASAP7_75t_R output2166 (.A(net2166),
    .Y(io_outs_down_0[58]));
 BUFx2_ASAP7_75t_R output2167 (.A(net2167),
    .Y(io_outs_down_0[59]));
 BUFx2_ASAP7_75t_R output2168 (.A(net2168),
    .Y(io_outs_down_0[5]));
 BUFx2_ASAP7_75t_R output2169 (.A(net2169),
    .Y(io_outs_down_0[60]));
 BUFx2_ASAP7_75t_R output2170 (.A(net2170),
    .Y(io_outs_down_0[61]));
 BUFx2_ASAP7_75t_R output2171 (.A(net2171),
    .Y(io_outs_down_0[62]));
 BUFx2_ASAP7_75t_R output2172 (.A(net2172),
    .Y(io_outs_down_0[63]));
 BUFx2_ASAP7_75t_R output2173 (.A(net2173),
    .Y(io_outs_down_0[6]));
 BUFx2_ASAP7_75t_R output2174 (.A(net2174),
    .Y(io_outs_down_0[7]));
 BUFx2_ASAP7_75t_R output2175 (.A(net2175),
    .Y(io_outs_down_0[8]));
 BUFx2_ASAP7_75t_R output2176 (.A(net2176),
    .Y(io_outs_down_0[9]));
 BUFx2_ASAP7_75t_R output2177 (.A(net2177),
    .Y(io_outs_down_1[0]));
 BUFx2_ASAP7_75t_R output2178 (.A(net2178),
    .Y(io_outs_down_1[10]));
 BUFx2_ASAP7_75t_R output2179 (.A(net2179),
    .Y(io_outs_down_1[11]));
 BUFx2_ASAP7_75t_R output2180 (.A(net2180),
    .Y(io_outs_down_1[12]));
 BUFx2_ASAP7_75t_R output2181 (.A(net2181),
    .Y(io_outs_down_1[13]));
 BUFx2_ASAP7_75t_R output2182 (.A(net2182),
    .Y(io_outs_down_1[14]));
 BUFx2_ASAP7_75t_R output2183 (.A(net2183),
    .Y(io_outs_down_1[15]));
 BUFx2_ASAP7_75t_R output2184 (.A(net2184),
    .Y(io_outs_down_1[16]));
 BUFx2_ASAP7_75t_R output2185 (.A(net2185),
    .Y(io_outs_down_1[17]));
 BUFx2_ASAP7_75t_R output2186 (.A(net2186),
    .Y(io_outs_down_1[18]));
 BUFx2_ASAP7_75t_R output2187 (.A(net2187),
    .Y(io_outs_down_1[19]));
 BUFx2_ASAP7_75t_R output2188 (.A(net2188),
    .Y(io_outs_down_1[1]));
 BUFx2_ASAP7_75t_R output2189 (.A(net2189),
    .Y(io_outs_down_1[20]));
 BUFx2_ASAP7_75t_R output2190 (.A(net2190),
    .Y(io_outs_down_1[21]));
 BUFx2_ASAP7_75t_R output2191 (.A(net2191),
    .Y(io_outs_down_1[22]));
 BUFx2_ASAP7_75t_R output2192 (.A(net2192),
    .Y(io_outs_down_1[23]));
 BUFx2_ASAP7_75t_R output2193 (.A(net2193),
    .Y(io_outs_down_1[24]));
 BUFx2_ASAP7_75t_R output2194 (.A(net2194),
    .Y(io_outs_down_1[25]));
 BUFx2_ASAP7_75t_R output2195 (.A(net2195),
    .Y(io_outs_down_1[26]));
 BUFx2_ASAP7_75t_R output2196 (.A(net2196),
    .Y(io_outs_down_1[27]));
 BUFx2_ASAP7_75t_R output2197 (.A(net2197),
    .Y(io_outs_down_1[28]));
 BUFx2_ASAP7_75t_R output2198 (.A(net2198),
    .Y(io_outs_down_1[29]));
 BUFx2_ASAP7_75t_R output2199 (.A(net2199),
    .Y(io_outs_down_1[2]));
 BUFx2_ASAP7_75t_R output2200 (.A(net2200),
    .Y(io_outs_down_1[30]));
 BUFx2_ASAP7_75t_R output2201 (.A(net2201),
    .Y(io_outs_down_1[31]));
 BUFx2_ASAP7_75t_R output2202 (.A(net2202),
    .Y(io_outs_down_1[32]));
 BUFx2_ASAP7_75t_R output2203 (.A(net2203),
    .Y(io_outs_down_1[33]));
 BUFx2_ASAP7_75t_R output2204 (.A(net2204),
    .Y(io_outs_down_1[34]));
 BUFx2_ASAP7_75t_R output2205 (.A(net2205),
    .Y(io_outs_down_1[35]));
 BUFx2_ASAP7_75t_R output2206 (.A(net2206),
    .Y(io_outs_down_1[36]));
 BUFx2_ASAP7_75t_R output2207 (.A(net2207),
    .Y(io_outs_down_1[37]));
 BUFx2_ASAP7_75t_R output2208 (.A(net2208),
    .Y(io_outs_down_1[38]));
 BUFx2_ASAP7_75t_R output2209 (.A(net2209),
    .Y(io_outs_down_1[39]));
 BUFx2_ASAP7_75t_R output2210 (.A(net2210),
    .Y(io_outs_down_1[3]));
 BUFx2_ASAP7_75t_R output2211 (.A(net2211),
    .Y(io_outs_down_1[40]));
 BUFx2_ASAP7_75t_R output2212 (.A(net2212),
    .Y(io_outs_down_1[41]));
 BUFx2_ASAP7_75t_R output2213 (.A(net2213),
    .Y(io_outs_down_1[42]));
 BUFx2_ASAP7_75t_R output2214 (.A(net2214),
    .Y(io_outs_down_1[43]));
 BUFx2_ASAP7_75t_R output2215 (.A(net2215),
    .Y(io_outs_down_1[44]));
 BUFx2_ASAP7_75t_R output2216 (.A(net2216),
    .Y(io_outs_down_1[45]));
 BUFx2_ASAP7_75t_R output2217 (.A(net2217),
    .Y(io_outs_down_1[46]));
 BUFx2_ASAP7_75t_R output2218 (.A(net2218),
    .Y(io_outs_down_1[47]));
 BUFx2_ASAP7_75t_R output2219 (.A(net2219),
    .Y(io_outs_down_1[48]));
 BUFx2_ASAP7_75t_R output2220 (.A(net2220),
    .Y(io_outs_down_1[49]));
 BUFx2_ASAP7_75t_R output2221 (.A(net2221),
    .Y(io_outs_down_1[4]));
 BUFx2_ASAP7_75t_R output2222 (.A(net2222),
    .Y(io_outs_down_1[50]));
 BUFx2_ASAP7_75t_R output2223 (.A(net2223),
    .Y(io_outs_down_1[51]));
 BUFx2_ASAP7_75t_R output2224 (.A(net2224),
    .Y(io_outs_down_1[52]));
 BUFx2_ASAP7_75t_R output2225 (.A(net2225),
    .Y(io_outs_down_1[53]));
 BUFx2_ASAP7_75t_R output2226 (.A(net2226),
    .Y(io_outs_down_1[54]));
 BUFx2_ASAP7_75t_R output2227 (.A(net2227),
    .Y(io_outs_down_1[55]));
 BUFx2_ASAP7_75t_R output2228 (.A(net2228),
    .Y(io_outs_down_1[56]));
 BUFx2_ASAP7_75t_R output2229 (.A(net2229),
    .Y(io_outs_down_1[57]));
 BUFx2_ASAP7_75t_R output2230 (.A(net2230),
    .Y(io_outs_down_1[58]));
 BUFx2_ASAP7_75t_R output2231 (.A(net2231),
    .Y(io_outs_down_1[59]));
 BUFx2_ASAP7_75t_R output2232 (.A(net2232),
    .Y(io_outs_down_1[5]));
 BUFx2_ASAP7_75t_R output2233 (.A(net2233),
    .Y(io_outs_down_1[60]));
 BUFx2_ASAP7_75t_R output2234 (.A(net2234),
    .Y(io_outs_down_1[61]));
 BUFx2_ASAP7_75t_R output2235 (.A(net2235),
    .Y(io_outs_down_1[62]));
 BUFx2_ASAP7_75t_R output2236 (.A(net2236),
    .Y(io_outs_down_1[63]));
 BUFx2_ASAP7_75t_R output2237 (.A(net2237),
    .Y(io_outs_down_1[6]));
 BUFx2_ASAP7_75t_R output2238 (.A(net2238),
    .Y(io_outs_down_1[7]));
 BUFx2_ASAP7_75t_R output2239 (.A(net2239),
    .Y(io_outs_down_1[8]));
 BUFx2_ASAP7_75t_R output2240 (.A(net2240),
    .Y(io_outs_down_1[9]));
 BUFx2_ASAP7_75t_R output2241 (.A(net2241),
    .Y(io_outs_down_2[0]));
 BUFx2_ASAP7_75t_R output2242 (.A(net2242),
    .Y(io_outs_down_2[10]));
 BUFx2_ASAP7_75t_R output2243 (.A(net2243),
    .Y(io_outs_down_2[11]));
 BUFx2_ASAP7_75t_R output2244 (.A(net2244),
    .Y(io_outs_down_2[12]));
 BUFx2_ASAP7_75t_R output2245 (.A(net2245),
    .Y(io_outs_down_2[13]));
 BUFx2_ASAP7_75t_R output2246 (.A(net2246),
    .Y(io_outs_down_2[14]));
 BUFx2_ASAP7_75t_R output2247 (.A(net2247),
    .Y(io_outs_down_2[15]));
 BUFx2_ASAP7_75t_R output2248 (.A(net2248),
    .Y(io_outs_down_2[16]));
 BUFx2_ASAP7_75t_R output2249 (.A(net2249),
    .Y(io_outs_down_2[17]));
 BUFx2_ASAP7_75t_R output2250 (.A(net2250),
    .Y(io_outs_down_2[18]));
 BUFx2_ASAP7_75t_R output2251 (.A(net2251),
    .Y(io_outs_down_2[19]));
 BUFx2_ASAP7_75t_R output2252 (.A(net2252),
    .Y(io_outs_down_2[1]));
 BUFx2_ASAP7_75t_R output2253 (.A(net2253),
    .Y(io_outs_down_2[20]));
 BUFx2_ASAP7_75t_R output2254 (.A(net2254),
    .Y(io_outs_down_2[21]));
 BUFx2_ASAP7_75t_R output2255 (.A(net2255),
    .Y(io_outs_down_2[22]));
 BUFx2_ASAP7_75t_R output2256 (.A(net2256),
    .Y(io_outs_down_2[23]));
 BUFx2_ASAP7_75t_R output2257 (.A(net2257),
    .Y(io_outs_down_2[24]));
 BUFx2_ASAP7_75t_R output2258 (.A(net2258),
    .Y(io_outs_down_2[25]));
 BUFx2_ASAP7_75t_R output2259 (.A(net2259),
    .Y(io_outs_down_2[26]));
 BUFx2_ASAP7_75t_R output2260 (.A(net2260),
    .Y(io_outs_down_2[27]));
 BUFx2_ASAP7_75t_R output2261 (.A(net2261),
    .Y(io_outs_down_2[28]));
 BUFx2_ASAP7_75t_R output2262 (.A(net2262),
    .Y(io_outs_down_2[29]));
 BUFx2_ASAP7_75t_R output2263 (.A(net2263),
    .Y(io_outs_down_2[2]));
 BUFx2_ASAP7_75t_R output2264 (.A(net2264),
    .Y(io_outs_down_2[30]));
 BUFx2_ASAP7_75t_R output2265 (.A(net2265),
    .Y(io_outs_down_2[31]));
 BUFx2_ASAP7_75t_R output2266 (.A(net2266),
    .Y(io_outs_down_2[32]));
 BUFx2_ASAP7_75t_R output2267 (.A(net2267),
    .Y(io_outs_down_2[33]));
 BUFx2_ASAP7_75t_R output2268 (.A(net2268),
    .Y(io_outs_down_2[34]));
 BUFx2_ASAP7_75t_R output2269 (.A(net2269),
    .Y(io_outs_down_2[35]));
 BUFx2_ASAP7_75t_R output2270 (.A(net2270),
    .Y(io_outs_down_2[36]));
 BUFx2_ASAP7_75t_R output2271 (.A(net2271),
    .Y(io_outs_down_2[37]));
 BUFx2_ASAP7_75t_R output2272 (.A(net2272),
    .Y(io_outs_down_2[38]));
 BUFx2_ASAP7_75t_R output2273 (.A(net2273),
    .Y(io_outs_down_2[39]));
 BUFx2_ASAP7_75t_R output2274 (.A(net2274),
    .Y(io_outs_down_2[3]));
 BUFx2_ASAP7_75t_R output2275 (.A(net2275),
    .Y(io_outs_down_2[40]));
 BUFx2_ASAP7_75t_R output2276 (.A(net2276),
    .Y(io_outs_down_2[41]));
 BUFx2_ASAP7_75t_R output2277 (.A(net2277),
    .Y(io_outs_down_2[42]));
 BUFx2_ASAP7_75t_R output2278 (.A(net2278),
    .Y(io_outs_down_2[43]));
 BUFx2_ASAP7_75t_R output2279 (.A(net2279),
    .Y(io_outs_down_2[44]));
 BUFx2_ASAP7_75t_R output2280 (.A(net2280),
    .Y(io_outs_down_2[45]));
 BUFx2_ASAP7_75t_R output2281 (.A(net2281),
    .Y(io_outs_down_2[46]));
 BUFx2_ASAP7_75t_R output2282 (.A(net2282),
    .Y(io_outs_down_2[47]));
 BUFx2_ASAP7_75t_R output2283 (.A(net2283),
    .Y(io_outs_down_2[48]));
 BUFx2_ASAP7_75t_R output2284 (.A(net2284),
    .Y(io_outs_down_2[49]));
 BUFx2_ASAP7_75t_R output2285 (.A(net2285),
    .Y(io_outs_down_2[4]));
 BUFx2_ASAP7_75t_R output2286 (.A(net2286),
    .Y(io_outs_down_2[50]));
 BUFx2_ASAP7_75t_R output2287 (.A(net2287),
    .Y(io_outs_down_2[51]));
 BUFx2_ASAP7_75t_R output2288 (.A(net2288),
    .Y(io_outs_down_2[52]));
 BUFx2_ASAP7_75t_R output2289 (.A(net2289),
    .Y(io_outs_down_2[53]));
 BUFx2_ASAP7_75t_R output2290 (.A(net2290),
    .Y(io_outs_down_2[54]));
 BUFx2_ASAP7_75t_R output2291 (.A(net2291),
    .Y(io_outs_down_2[55]));
 BUFx2_ASAP7_75t_R output2292 (.A(net2292),
    .Y(io_outs_down_2[56]));
 BUFx2_ASAP7_75t_R output2293 (.A(net2293),
    .Y(io_outs_down_2[57]));
 BUFx2_ASAP7_75t_R output2294 (.A(net2294),
    .Y(io_outs_down_2[58]));
 BUFx2_ASAP7_75t_R output2295 (.A(net2295),
    .Y(io_outs_down_2[59]));
 BUFx2_ASAP7_75t_R output2296 (.A(net2296),
    .Y(io_outs_down_2[5]));
 BUFx2_ASAP7_75t_R output2297 (.A(net2297),
    .Y(io_outs_down_2[60]));
 BUFx2_ASAP7_75t_R output2298 (.A(net2298),
    .Y(io_outs_down_2[61]));
 BUFx2_ASAP7_75t_R output2299 (.A(net2299),
    .Y(io_outs_down_2[62]));
 BUFx2_ASAP7_75t_R output2300 (.A(net2300),
    .Y(io_outs_down_2[63]));
 BUFx2_ASAP7_75t_R output2301 (.A(net2301),
    .Y(io_outs_down_2[6]));
 BUFx2_ASAP7_75t_R output2302 (.A(net2302),
    .Y(io_outs_down_2[7]));
 BUFx2_ASAP7_75t_R output2303 (.A(net2303),
    .Y(io_outs_down_2[8]));
 BUFx2_ASAP7_75t_R output2304 (.A(net2304),
    .Y(io_outs_down_2[9]));
 BUFx2_ASAP7_75t_R output2305 (.A(net2305),
    .Y(io_outs_down_3[0]));
 BUFx2_ASAP7_75t_R output2306 (.A(net2306),
    .Y(io_outs_down_3[10]));
 BUFx2_ASAP7_75t_R output2307 (.A(net2307),
    .Y(io_outs_down_3[11]));
 BUFx2_ASAP7_75t_R output2308 (.A(net2308),
    .Y(io_outs_down_3[12]));
 BUFx2_ASAP7_75t_R output2309 (.A(net2309),
    .Y(io_outs_down_3[13]));
 BUFx2_ASAP7_75t_R output2310 (.A(net2310),
    .Y(io_outs_down_3[14]));
 BUFx2_ASAP7_75t_R output2311 (.A(net2311),
    .Y(io_outs_down_3[15]));
 BUFx2_ASAP7_75t_R output2312 (.A(net2312),
    .Y(io_outs_down_3[16]));
 BUFx2_ASAP7_75t_R output2313 (.A(net2313),
    .Y(io_outs_down_3[17]));
 BUFx2_ASAP7_75t_R output2314 (.A(net2314),
    .Y(io_outs_down_3[18]));
 BUFx2_ASAP7_75t_R output2315 (.A(net2315),
    .Y(io_outs_down_3[19]));
 BUFx2_ASAP7_75t_R output2316 (.A(net2316),
    .Y(io_outs_down_3[1]));
 BUFx2_ASAP7_75t_R output2317 (.A(net2317),
    .Y(io_outs_down_3[20]));
 BUFx2_ASAP7_75t_R output2318 (.A(net2318),
    .Y(io_outs_down_3[21]));
 BUFx2_ASAP7_75t_R output2319 (.A(net2319),
    .Y(io_outs_down_3[22]));
 BUFx2_ASAP7_75t_R output2320 (.A(net2320),
    .Y(io_outs_down_3[23]));
 BUFx2_ASAP7_75t_R output2321 (.A(net2321),
    .Y(io_outs_down_3[24]));
 BUFx2_ASAP7_75t_R output2322 (.A(net2322),
    .Y(io_outs_down_3[25]));
 BUFx2_ASAP7_75t_R output2323 (.A(net2323),
    .Y(io_outs_down_3[26]));
 BUFx2_ASAP7_75t_R output2324 (.A(net2324),
    .Y(io_outs_down_3[27]));
 BUFx2_ASAP7_75t_R output2325 (.A(net2325),
    .Y(io_outs_down_3[28]));
 BUFx2_ASAP7_75t_R output2326 (.A(net2326),
    .Y(io_outs_down_3[29]));
 BUFx2_ASAP7_75t_R output2327 (.A(net2327),
    .Y(io_outs_down_3[2]));
 BUFx2_ASAP7_75t_R output2328 (.A(net2328),
    .Y(io_outs_down_3[30]));
 BUFx2_ASAP7_75t_R output2329 (.A(net2329),
    .Y(io_outs_down_3[31]));
 BUFx2_ASAP7_75t_R output2330 (.A(net2330),
    .Y(io_outs_down_3[32]));
 BUFx2_ASAP7_75t_R output2331 (.A(net2331),
    .Y(io_outs_down_3[33]));
 BUFx2_ASAP7_75t_R output2332 (.A(net2332),
    .Y(io_outs_down_3[34]));
 BUFx2_ASAP7_75t_R output2333 (.A(net2333),
    .Y(io_outs_down_3[35]));
 BUFx2_ASAP7_75t_R output2334 (.A(net2334),
    .Y(io_outs_down_3[36]));
 BUFx2_ASAP7_75t_R output2335 (.A(net2335),
    .Y(io_outs_down_3[37]));
 BUFx2_ASAP7_75t_R output2336 (.A(net2336),
    .Y(io_outs_down_3[38]));
 BUFx2_ASAP7_75t_R output2337 (.A(net2337),
    .Y(io_outs_down_3[39]));
 BUFx2_ASAP7_75t_R output2338 (.A(net2338),
    .Y(io_outs_down_3[3]));
 BUFx2_ASAP7_75t_R output2339 (.A(net2339),
    .Y(io_outs_down_3[40]));
 BUFx2_ASAP7_75t_R output2340 (.A(net2340),
    .Y(io_outs_down_3[41]));
 BUFx2_ASAP7_75t_R output2341 (.A(net2341),
    .Y(io_outs_down_3[42]));
 BUFx2_ASAP7_75t_R output2342 (.A(net2342),
    .Y(io_outs_down_3[43]));
 BUFx2_ASAP7_75t_R output2343 (.A(net2343),
    .Y(io_outs_down_3[44]));
 BUFx2_ASAP7_75t_R output2344 (.A(net2344),
    .Y(io_outs_down_3[45]));
 BUFx2_ASAP7_75t_R output2345 (.A(net2345),
    .Y(io_outs_down_3[46]));
 BUFx2_ASAP7_75t_R output2346 (.A(net2346),
    .Y(io_outs_down_3[47]));
 BUFx2_ASAP7_75t_R output2347 (.A(net2347),
    .Y(io_outs_down_3[48]));
 BUFx2_ASAP7_75t_R output2348 (.A(net2348),
    .Y(io_outs_down_3[49]));
 BUFx2_ASAP7_75t_R output2349 (.A(net2349),
    .Y(io_outs_down_3[4]));
 BUFx2_ASAP7_75t_R output2350 (.A(net2350),
    .Y(io_outs_down_3[50]));
 BUFx2_ASAP7_75t_R output2351 (.A(net2351),
    .Y(io_outs_down_3[51]));
 BUFx2_ASAP7_75t_R output2352 (.A(net2352),
    .Y(io_outs_down_3[52]));
 BUFx2_ASAP7_75t_R output2353 (.A(net2353),
    .Y(io_outs_down_3[53]));
 BUFx2_ASAP7_75t_R output2354 (.A(net2354),
    .Y(io_outs_down_3[54]));
 BUFx2_ASAP7_75t_R output2355 (.A(net2355),
    .Y(io_outs_down_3[55]));
 BUFx2_ASAP7_75t_R output2356 (.A(net2356),
    .Y(io_outs_down_3[56]));
 BUFx2_ASAP7_75t_R output2357 (.A(net2357),
    .Y(io_outs_down_3[57]));
 BUFx2_ASAP7_75t_R output2358 (.A(net2358),
    .Y(io_outs_down_3[58]));
 BUFx2_ASAP7_75t_R output2359 (.A(net2359),
    .Y(io_outs_down_3[59]));
 BUFx2_ASAP7_75t_R output2360 (.A(net2360),
    .Y(io_outs_down_3[5]));
 BUFx2_ASAP7_75t_R output2361 (.A(net2361),
    .Y(io_outs_down_3[60]));
 BUFx2_ASAP7_75t_R output2362 (.A(net2362),
    .Y(io_outs_down_3[61]));
 BUFx2_ASAP7_75t_R output2363 (.A(net2363),
    .Y(io_outs_down_3[62]));
 BUFx2_ASAP7_75t_R output2364 (.A(net2364),
    .Y(io_outs_down_3[63]));
 BUFx2_ASAP7_75t_R output2365 (.A(net2365),
    .Y(io_outs_down_3[6]));
 BUFx2_ASAP7_75t_R output2366 (.A(net2366),
    .Y(io_outs_down_3[7]));
 BUFx2_ASAP7_75t_R output2367 (.A(net2367),
    .Y(io_outs_down_3[8]));
 BUFx2_ASAP7_75t_R output2368 (.A(net2368),
    .Y(io_outs_down_3[9]));
 BUFx2_ASAP7_75t_R output2369 (.A(net2369),
    .Y(io_outs_down_4[0]));
 BUFx2_ASAP7_75t_R output2370 (.A(net2370),
    .Y(io_outs_down_4[10]));
 BUFx2_ASAP7_75t_R output2371 (.A(net2371),
    .Y(io_outs_down_4[11]));
 BUFx2_ASAP7_75t_R output2372 (.A(net2372),
    .Y(io_outs_down_4[12]));
 BUFx2_ASAP7_75t_R output2373 (.A(net2373),
    .Y(io_outs_down_4[13]));
 BUFx2_ASAP7_75t_R output2374 (.A(net2374),
    .Y(io_outs_down_4[14]));
 BUFx2_ASAP7_75t_R output2375 (.A(net2375),
    .Y(io_outs_down_4[15]));
 BUFx2_ASAP7_75t_R output2376 (.A(net2376),
    .Y(io_outs_down_4[16]));
 BUFx2_ASAP7_75t_R output2377 (.A(net2377),
    .Y(io_outs_down_4[17]));
 BUFx2_ASAP7_75t_R output2378 (.A(net2378),
    .Y(io_outs_down_4[18]));
 BUFx2_ASAP7_75t_R output2379 (.A(net2379),
    .Y(io_outs_down_4[19]));
 BUFx2_ASAP7_75t_R output2380 (.A(net2380),
    .Y(io_outs_down_4[1]));
 BUFx2_ASAP7_75t_R output2381 (.A(net2381),
    .Y(io_outs_down_4[20]));
 BUFx2_ASAP7_75t_R output2382 (.A(net2382),
    .Y(io_outs_down_4[21]));
 BUFx2_ASAP7_75t_R output2383 (.A(net2383),
    .Y(io_outs_down_4[22]));
 BUFx2_ASAP7_75t_R output2384 (.A(net2384),
    .Y(io_outs_down_4[23]));
 BUFx2_ASAP7_75t_R output2385 (.A(net2385),
    .Y(io_outs_down_4[24]));
 BUFx2_ASAP7_75t_R output2386 (.A(net2386),
    .Y(io_outs_down_4[25]));
 BUFx2_ASAP7_75t_R output2387 (.A(net2387),
    .Y(io_outs_down_4[26]));
 BUFx2_ASAP7_75t_R output2388 (.A(net2388),
    .Y(io_outs_down_4[27]));
 BUFx2_ASAP7_75t_R output2389 (.A(net2389),
    .Y(io_outs_down_4[28]));
 BUFx2_ASAP7_75t_R output2390 (.A(net2390),
    .Y(io_outs_down_4[29]));
 BUFx2_ASAP7_75t_R output2391 (.A(net2391),
    .Y(io_outs_down_4[2]));
 BUFx2_ASAP7_75t_R output2392 (.A(net2392),
    .Y(io_outs_down_4[30]));
 BUFx2_ASAP7_75t_R output2393 (.A(net2393),
    .Y(io_outs_down_4[31]));
 BUFx2_ASAP7_75t_R output2394 (.A(net2394),
    .Y(io_outs_down_4[32]));
 BUFx2_ASAP7_75t_R output2395 (.A(net2395),
    .Y(io_outs_down_4[33]));
 BUFx2_ASAP7_75t_R output2396 (.A(net2396),
    .Y(io_outs_down_4[34]));
 BUFx2_ASAP7_75t_R output2397 (.A(net2397),
    .Y(io_outs_down_4[35]));
 BUFx2_ASAP7_75t_R output2398 (.A(net2398),
    .Y(io_outs_down_4[36]));
 BUFx2_ASAP7_75t_R output2399 (.A(net2399),
    .Y(io_outs_down_4[37]));
 BUFx2_ASAP7_75t_R output2400 (.A(net2400),
    .Y(io_outs_down_4[38]));
 BUFx2_ASAP7_75t_R output2401 (.A(net2401),
    .Y(io_outs_down_4[39]));
 BUFx2_ASAP7_75t_R output2402 (.A(net2402),
    .Y(io_outs_down_4[3]));
 BUFx2_ASAP7_75t_R output2403 (.A(net2403),
    .Y(io_outs_down_4[40]));
 BUFx2_ASAP7_75t_R output2404 (.A(net2404),
    .Y(io_outs_down_4[41]));
 BUFx2_ASAP7_75t_R output2405 (.A(net2405),
    .Y(io_outs_down_4[42]));
 BUFx2_ASAP7_75t_R output2406 (.A(net2406),
    .Y(io_outs_down_4[43]));
 BUFx2_ASAP7_75t_R output2407 (.A(net2407),
    .Y(io_outs_down_4[44]));
 BUFx2_ASAP7_75t_R output2408 (.A(net2408),
    .Y(io_outs_down_4[45]));
 BUFx2_ASAP7_75t_R output2409 (.A(net2409),
    .Y(io_outs_down_4[46]));
 BUFx2_ASAP7_75t_R output2410 (.A(net2410),
    .Y(io_outs_down_4[47]));
 BUFx2_ASAP7_75t_R output2411 (.A(net2411),
    .Y(io_outs_down_4[48]));
 BUFx2_ASAP7_75t_R output2412 (.A(net2412),
    .Y(io_outs_down_4[49]));
 BUFx2_ASAP7_75t_R output2413 (.A(net2413),
    .Y(io_outs_down_4[4]));
 BUFx2_ASAP7_75t_R output2414 (.A(net2414),
    .Y(io_outs_down_4[50]));
 BUFx2_ASAP7_75t_R output2415 (.A(net2415),
    .Y(io_outs_down_4[51]));
 BUFx2_ASAP7_75t_R output2416 (.A(net2416),
    .Y(io_outs_down_4[52]));
 BUFx2_ASAP7_75t_R output2417 (.A(net2417),
    .Y(io_outs_down_4[53]));
 BUFx2_ASAP7_75t_R output2418 (.A(net2418),
    .Y(io_outs_down_4[54]));
 BUFx2_ASAP7_75t_R output2419 (.A(net2419),
    .Y(io_outs_down_4[55]));
 BUFx2_ASAP7_75t_R output2420 (.A(net2420),
    .Y(io_outs_down_4[56]));
 BUFx2_ASAP7_75t_R output2421 (.A(net2421),
    .Y(io_outs_down_4[57]));
 BUFx2_ASAP7_75t_R output2422 (.A(net2422),
    .Y(io_outs_down_4[58]));
 BUFx2_ASAP7_75t_R output2423 (.A(net2423),
    .Y(io_outs_down_4[59]));
 BUFx2_ASAP7_75t_R output2424 (.A(net2424),
    .Y(io_outs_down_4[5]));
 BUFx2_ASAP7_75t_R output2425 (.A(net2425),
    .Y(io_outs_down_4[60]));
 BUFx2_ASAP7_75t_R output2426 (.A(net2426),
    .Y(io_outs_down_4[61]));
 BUFx2_ASAP7_75t_R output2427 (.A(net2427),
    .Y(io_outs_down_4[62]));
 BUFx2_ASAP7_75t_R output2428 (.A(net2428),
    .Y(io_outs_down_4[63]));
 BUFx2_ASAP7_75t_R output2429 (.A(net2429),
    .Y(io_outs_down_4[6]));
 BUFx2_ASAP7_75t_R output2430 (.A(net2430),
    .Y(io_outs_down_4[7]));
 BUFx2_ASAP7_75t_R output2431 (.A(net2431),
    .Y(io_outs_down_4[8]));
 BUFx2_ASAP7_75t_R output2432 (.A(net2432),
    .Y(io_outs_down_4[9]));
 BUFx2_ASAP7_75t_R output2433 (.A(net2433),
    .Y(io_outs_down_5[0]));
 BUFx2_ASAP7_75t_R output2434 (.A(net2434),
    .Y(io_outs_down_5[10]));
 BUFx2_ASAP7_75t_R output2435 (.A(net2435),
    .Y(io_outs_down_5[11]));
 BUFx2_ASAP7_75t_R output2436 (.A(net2436),
    .Y(io_outs_down_5[12]));
 BUFx2_ASAP7_75t_R output2437 (.A(net2437),
    .Y(io_outs_down_5[13]));
 BUFx2_ASAP7_75t_R output2438 (.A(net2438),
    .Y(io_outs_down_5[14]));
 BUFx2_ASAP7_75t_R output2439 (.A(net2439),
    .Y(io_outs_down_5[15]));
 BUFx2_ASAP7_75t_R output2440 (.A(net2440),
    .Y(io_outs_down_5[16]));
 BUFx2_ASAP7_75t_R output2441 (.A(net2441),
    .Y(io_outs_down_5[17]));
 BUFx2_ASAP7_75t_R output2442 (.A(net2442),
    .Y(io_outs_down_5[18]));
 BUFx2_ASAP7_75t_R output2443 (.A(net2443),
    .Y(io_outs_down_5[19]));
 BUFx2_ASAP7_75t_R output2444 (.A(net2444),
    .Y(io_outs_down_5[1]));
 BUFx2_ASAP7_75t_R output2445 (.A(net2445),
    .Y(io_outs_down_5[20]));
 BUFx2_ASAP7_75t_R output2446 (.A(net2446),
    .Y(io_outs_down_5[21]));
 BUFx2_ASAP7_75t_R output2447 (.A(net2447),
    .Y(io_outs_down_5[22]));
 BUFx2_ASAP7_75t_R output2448 (.A(net2448),
    .Y(io_outs_down_5[23]));
 BUFx2_ASAP7_75t_R output2449 (.A(net2449),
    .Y(io_outs_down_5[24]));
 BUFx2_ASAP7_75t_R output2450 (.A(net2450),
    .Y(io_outs_down_5[25]));
 BUFx2_ASAP7_75t_R output2451 (.A(net2451),
    .Y(io_outs_down_5[26]));
 BUFx2_ASAP7_75t_R output2452 (.A(net2452),
    .Y(io_outs_down_5[27]));
 BUFx2_ASAP7_75t_R output2453 (.A(net2453),
    .Y(io_outs_down_5[28]));
 BUFx2_ASAP7_75t_R output2454 (.A(net2454),
    .Y(io_outs_down_5[29]));
 BUFx2_ASAP7_75t_R output2455 (.A(net2455),
    .Y(io_outs_down_5[2]));
 BUFx2_ASAP7_75t_R output2456 (.A(net2456),
    .Y(io_outs_down_5[30]));
 BUFx2_ASAP7_75t_R output2457 (.A(net2457),
    .Y(io_outs_down_5[31]));
 BUFx2_ASAP7_75t_R output2458 (.A(net2458),
    .Y(io_outs_down_5[32]));
 BUFx2_ASAP7_75t_R output2459 (.A(net2459),
    .Y(io_outs_down_5[33]));
 BUFx2_ASAP7_75t_R output2460 (.A(net2460),
    .Y(io_outs_down_5[34]));
 BUFx2_ASAP7_75t_R output2461 (.A(net2461),
    .Y(io_outs_down_5[35]));
 BUFx2_ASAP7_75t_R output2462 (.A(net2462),
    .Y(io_outs_down_5[36]));
 BUFx2_ASAP7_75t_R output2463 (.A(net2463),
    .Y(io_outs_down_5[37]));
 BUFx2_ASAP7_75t_R output2464 (.A(net2464),
    .Y(io_outs_down_5[38]));
 BUFx2_ASAP7_75t_R output2465 (.A(net2465),
    .Y(io_outs_down_5[39]));
 BUFx2_ASAP7_75t_R output2466 (.A(net2466),
    .Y(io_outs_down_5[3]));
 BUFx2_ASAP7_75t_R output2467 (.A(net2467),
    .Y(io_outs_down_5[40]));
 BUFx2_ASAP7_75t_R output2468 (.A(net2468),
    .Y(io_outs_down_5[41]));
 BUFx2_ASAP7_75t_R output2469 (.A(net2469),
    .Y(io_outs_down_5[42]));
 BUFx2_ASAP7_75t_R output2470 (.A(net2470),
    .Y(io_outs_down_5[43]));
 BUFx2_ASAP7_75t_R output2471 (.A(net2471),
    .Y(io_outs_down_5[44]));
 BUFx2_ASAP7_75t_R output2472 (.A(net2472),
    .Y(io_outs_down_5[45]));
 BUFx2_ASAP7_75t_R output2473 (.A(net2473),
    .Y(io_outs_down_5[46]));
 BUFx2_ASAP7_75t_R output2474 (.A(net2474),
    .Y(io_outs_down_5[47]));
 BUFx2_ASAP7_75t_R output2475 (.A(net2475),
    .Y(io_outs_down_5[48]));
 BUFx2_ASAP7_75t_R output2476 (.A(net2476),
    .Y(io_outs_down_5[49]));
 BUFx2_ASAP7_75t_R output2477 (.A(net2477),
    .Y(io_outs_down_5[4]));
 BUFx2_ASAP7_75t_R output2478 (.A(net2478),
    .Y(io_outs_down_5[50]));
 BUFx2_ASAP7_75t_R output2479 (.A(net2479),
    .Y(io_outs_down_5[51]));
 BUFx2_ASAP7_75t_R output2480 (.A(net2480),
    .Y(io_outs_down_5[52]));
 BUFx2_ASAP7_75t_R output2481 (.A(net2481),
    .Y(io_outs_down_5[53]));
 BUFx2_ASAP7_75t_R output2482 (.A(net2482),
    .Y(io_outs_down_5[54]));
 BUFx2_ASAP7_75t_R output2483 (.A(net2483),
    .Y(io_outs_down_5[55]));
 BUFx2_ASAP7_75t_R output2484 (.A(net2484),
    .Y(io_outs_down_5[56]));
 BUFx2_ASAP7_75t_R output2485 (.A(net2485),
    .Y(io_outs_down_5[57]));
 BUFx2_ASAP7_75t_R output2486 (.A(net2486),
    .Y(io_outs_down_5[58]));
 BUFx2_ASAP7_75t_R output2487 (.A(net2487),
    .Y(io_outs_down_5[59]));
 BUFx2_ASAP7_75t_R output2488 (.A(net2488),
    .Y(io_outs_down_5[5]));
 BUFx2_ASAP7_75t_R output2489 (.A(net2489),
    .Y(io_outs_down_5[60]));
 BUFx2_ASAP7_75t_R output2490 (.A(net2490),
    .Y(io_outs_down_5[61]));
 BUFx2_ASAP7_75t_R output2491 (.A(net2491),
    .Y(io_outs_down_5[62]));
 BUFx2_ASAP7_75t_R output2492 (.A(net2492),
    .Y(io_outs_down_5[63]));
 BUFx2_ASAP7_75t_R output2493 (.A(net2493),
    .Y(io_outs_down_5[6]));
 BUFx2_ASAP7_75t_R output2494 (.A(net2494),
    .Y(io_outs_down_5[7]));
 BUFx2_ASAP7_75t_R output2495 (.A(net2495),
    .Y(io_outs_down_5[8]));
 BUFx2_ASAP7_75t_R output2496 (.A(net2496),
    .Y(io_outs_down_5[9]));
 BUFx2_ASAP7_75t_R output2497 (.A(net2497),
    .Y(io_outs_down_6[0]));
 BUFx2_ASAP7_75t_R output2498 (.A(net2498),
    .Y(io_outs_down_6[10]));
 BUFx2_ASAP7_75t_R output2499 (.A(net2499),
    .Y(io_outs_down_6[11]));
 BUFx2_ASAP7_75t_R output2500 (.A(net2500),
    .Y(io_outs_down_6[12]));
 BUFx2_ASAP7_75t_R output2501 (.A(net2501),
    .Y(io_outs_down_6[13]));
 BUFx2_ASAP7_75t_R output2502 (.A(net2502),
    .Y(io_outs_down_6[14]));
 BUFx2_ASAP7_75t_R output2503 (.A(net2503),
    .Y(io_outs_down_6[15]));
 BUFx2_ASAP7_75t_R output2504 (.A(net2504),
    .Y(io_outs_down_6[16]));
 BUFx2_ASAP7_75t_R output2505 (.A(net2505),
    .Y(io_outs_down_6[17]));
 BUFx2_ASAP7_75t_R output2506 (.A(net2506),
    .Y(io_outs_down_6[18]));
 BUFx2_ASAP7_75t_R output2507 (.A(net2507),
    .Y(io_outs_down_6[19]));
 BUFx2_ASAP7_75t_R output2508 (.A(net2508),
    .Y(io_outs_down_6[1]));
 BUFx2_ASAP7_75t_R output2509 (.A(net2509),
    .Y(io_outs_down_6[20]));
 BUFx2_ASAP7_75t_R output2510 (.A(net2510),
    .Y(io_outs_down_6[21]));
 BUFx2_ASAP7_75t_R output2511 (.A(net2511),
    .Y(io_outs_down_6[22]));
 BUFx2_ASAP7_75t_R output2512 (.A(net2512),
    .Y(io_outs_down_6[23]));
 BUFx2_ASAP7_75t_R output2513 (.A(net2513),
    .Y(io_outs_down_6[24]));
 BUFx2_ASAP7_75t_R output2514 (.A(net2514),
    .Y(io_outs_down_6[25]));
 BUFx2_ASAP7_75t_R output2515 (.A(net2515),
    .Y(io_outs_down_6[26]));
 BUFx2_ASAP7_75t_R output2516 (.A(net2516),
    .Y(io_outs_down_6[27]));
 BUFx2_ASAP7_75t_R output2517 (.A(net2517),
    .Y(io_outs_down_6[28]));
 BUFx2_ASAP7_75t_R output2518 (.A(net2518),
    .Y(io_outs_down_6[29]));
 BUFx2_ASAP7_75t_R output2519 (.A(net2519),
    .Y(io_outs_down_6[2]));
 BUFx2_ASAP7_75t_R output2520 (.A(net2520),
    .Y(io_outs_down_6[30]));
 BUFx2_ASAP7_75t_R output2521 (.A(net2521),
    .Y(io_outs_down_6[31]));
 BUFx2_ASAP7_75t_R output2522 (.A(net2522),
    .Y(io_outs_down_6[32]));
 BUFx2_ASAP7_75t_R output2523 (.A(net2523),
    .Y(io_outs_down_6[33]));
 BUFx2_ASAP7_75t_R output2524 (.A(net2524),
    .Y(io_outs_down_6[34]));
 BUFx2_ASAP7_75t_R output2525 (.A(net2525),
    .Y(io_outs_down_6[35]));
 BUFx2_ASAP7_75t_R output2526 (.A(net2526),
    .Y(io_outs_down_6[36]));
 BUFx2_ASAP7_75t_R output2527 (.A(net2527),
    .Y(io_outs_down_6[37]));
 BUFx2_ASAP7_75t_R output2528 (.A(net2528),
    .Y(io_outs_down_6[38]));
 BUFx2_ASAP7_75t_R output2529 (.A(net2529),
    .Y(io_outs_down_6[39]));
 BUFx2_ASAP7_75t_R output2530 (.A(net2530),
    .Y(io_outs_down_6[3]));
 BUFx2_ASAP7_75t_R output2531 (.A(net2531),
    .Y(io_outs_down_6[40]));
 BUFx2_ASAP7_75t_R output2532 (.A(net2532),
    .Y(io_outs_down_6[41]));
 BUFx2_ASAP7_75t_R output2533 (.A(net2533),
    .Y(io_outs_down_6[42]));
 BUFx2_ASAP7_75t_R output2534 (.A(net2534),
    .Y(io_outs_down_6[43]));
 BUFx2_ASAP7_75t_R output2535 (.A(net2535),
    .Y(io_outs_down_6[44]));
 BUFx2_ASAP7_75t_R output2536 (.A(net2536),
    .Y(io_outs_down_6[45]));
 BUFx2_ASAP7_75t_R output2537 (.A(net2537),
    .Y(io_outs_down_6[46]));
 BUFx2_ASAP7_75t_R output2538 (.A(net2538),
    .Y(io_outs_down_6[47]));
 BUFx2_ASAP7_75t_R output2539 (.A(net2539),
    .Y(io_outs_down_6[48]));
 BUFx2_ASAP7_75t_R output2540 (.A(net2540),
    .Y(io_outs_down_6[49]));
 BUFx2_ASAP7_75t_R output2541 (.A(net2541),
    .Y(io_outs_down_6[4]));
 BUFx2_ASAP7_75t_R output2542 (.A(net2542),
    .Y(io_outs_down_6[50]));
 BUFx2_ASAP7_75t_R output2543 (.A(net2543),
    .Y(io_outs_down_6[51]));
 BUFx2_ASAP7_75t_R output2544 (.A(net2544),
    .Y(io_outs_down_6[52]));
 BUFx2_ASAP7_75t_R output2545 (.A(net2545),
    .Y(io_outs_down_6[53]));
 BUFx2_ASAP7_75t_R output2546 (.A(net2546),
    .Y(io_outs_down_6[54]));
 BUFx2_ASAP7_75t_R output2547 (.A(net2547),
    .Y(io_outs_down_6[55]));
 BUFx2_ASAP7_75t_R output2548 (.A(net2548),
    .Y(io_outs_down_6[56]));
 BUFx2_ASAP7_75t_R output2549 (.A(net2549),
    .Y(io_outs_down_6[57]));
 BUFx2_ASAP7_75t_R output2550 (.A(net2550),
    .Y(io_outs_down_6[58]));
 BUFx2_ASAP7_75t_R output2551 (.A(net2551),
    .Y(io_outs_down_6[59]));
 BUFx2_ASAP7_75t_R output2552 (.A(net2552),
    .Y(io_outs_down_6[5]));
 BUFx2_ASAP7_75t_R output2553 (.A(net2553),
    .Y(io_outs_down_6[60]));
 BUFx2_ASAP7_75t_R output2554 (.A(net2554),
    .Y(io_outs_down_6[61]));
 BUFx2_ASAP7_75t_R output2555 (.A(net2555),
    .Y(io_outs_down_6[62]));
 BUFx2_ASAP7_75t_R output2556 (.A(net2556),
    .Y(io_outs_down_6[63]));
 BUFx2_ASAP7_75t_R output2557 (.A(net2557),
    .Y(io_outs_down_6[6]));
 BUFx2_ASAP7_75t_R output2558 (.A(net2558),
    .Y(io_outs_down_6[7]));
 BUFx2_ASAP7_75t_R output2559 (.A(net2559),
    .Y(io_outs_down_6[8]));
 BUFx2_ASAP7_75t_R output2560 (.A(net2560),
    .Y(io_outs_down_6[9]));
 BUFx2_ASAP7_75t_R output2561 (.A(net2561),
    .Y(io_outs_down_7[0]));
 BUFx2_ASAP7_75t_R output2562 (.A(net2562),
    .Y(io_outs_down_7[10]));
 BUFx2_ASAP7_75t_R output2563 (.A(net2563),
    .Y(io_outs_down_7[11]));
 BUFx2_ASAP7_75t_R output2564 (.A(net2564),
    .Y(io_outs_down_7[12]));
 BUFx2_ASAP7_75t_R output2565 (.A(net2565),
    .Y(io_outs_down_7[13]));
 BUFx2_ASAP7_75t_R output2566 (.A(net2566),
    .Y(io_outs_down_7[14]));
 BUFx2_ASAP7_75t_R output2567 (.A(net2567),
    .Y(io_outs_down_7[15]));
 BUFx2_ASAP7_75t_R output2568 (.A(net2568),
    .Y(io_outs_down_7[16]));
 BUFx2_ASAP7_75t_R output2569 (.A(net2569),
    .Y(io_outs_down_7[17]));
 BUFx2_ASAP7_75t_R output2570 (.A(net2570),
    .Y(io_outs_down_7[18]));
 BUFx2_ASAP7_75t_R output2571 (.A(net2571),
    .Y(io_outs_down_7[19]));
 BUFx2_ASAP7_75t_R output2572 (.A(net2572),
    .Y(io_outs_down_7[1]));
 BUFx2_ASAP7_75t_R output2573 (.A(net2573),
    .Y(io_outs_down_7[20]));
 BUFx2_ASAP7_75t_R output2574 (.A(net2574),
    .Y(io_outs_down_7[21]));
 BUFx2_ASAP7_75t_R output2575 (.A(net2575),
    .Y(io_outs_down_7[22]));
 BUFx2_ASAP7_75t_R output2576 (.A(net2576),
    .Y(io_outs_down_7[23]));
 BUFx2_ASAP7_75t_R output2577 (.A(net2577),
    .Y(io_outs_down_7[24]));
 BUFx2_ASAP7_75t_R output2578 (.A(net2578),
    .Y(io_outs_down_7[25]));
 BUFx2_ASAP7_75t_R output2579 (.A(net2579),
    .Y(io_outs_down_7[26]));
 BUFx2_ASAP7_75t_R output2580 (.A(net2580),
    .Y(io_outs_down_7[27]));
 BUFx2_ASAP7_75t_R output2581 (.A(net2581),
    .Y(io_outs_down_7[28]));
 BUFx2_ASAP7_75t_R output2582 (.A(net2582),
    .Y(io_outs_down_7[29]));
 BUFx2_ASAP7_75t_R output2583 (.A(net2583),
    .Y(io_outs_down_7[2]));
 BUFx2_ASAP7_75t_R output2584 (.A(net2584),
    .Y(io_outs_down_7[30]));
 BUFx2_ASAP7_75t_R output2585 (.A(net2585),
    .Y(io_outs_down_7[31]));
 BUFx2_ASAP7_75t_R output2586 (.A(net2586),
    .Y(io_outs_down_7[32]));
 BUFx2_ASAP7_75t_R output2587 (.A(net2587),
    .Y(io_outs_down_7[33]));
 BUFx2_ASAP7_75t_R output2588 (.A(net2588),
    .Y(io_outs_down_7[34]));
 BUFx2_ASAP7_75t_R output2589 (.A(net2589),
    .Y(io_outs_down_7[35]));
 BUFx2_ASAP7_75t_R output2590 (.A(net2590),
    .Y(io_outs_down_7[36]));
 BUFx2_ASAP7_75t_R output2591 (.A(net2591),
    .Y(io_outs_down_7[37]));
 BUFx2_ASAP7_75t_R output2592 (.A(net2592),
    .Y(io_outs_down_7[38]));
 BUFx2_ASAP7_75t_R output2593 (.A(net2593),
    .Y(io_outs_down_7[39]));
 BUFx2_ASAP7_75t_R output2594 (.A(net2594),
    .Y(io_outs_down_7[3]));
 BUFx2_ASAP7_75t_R output2595 (.A(net2595),
    .Y(io_outs_down_7[40]));
 BUFx2_ASAP7_75t_R output2596 (.A(net2596),
    .Y(io_outs_down_7[41]));
 BUFx2_ASAP7_75t_R output2597 (.A(net2597),
    .Y(io_outs_down_7[42]));
 BUFx2_ASAP7_75t_R output2598 (.A(net2598),
    .Y(io_outs_down_7[43]));
 BUFx2_ASAP7_75t_R output2599 (.A(net2599),
    .Y(io_outs_down_7[44]));
 BUFx2_ASAP7_75t_R output2600 (.A(net2600),
    .Y(io_outs_down_7[45]));
 BUFx2_ASAP7_75t_R output2601 (.A(net2601),
    .Y(io_outs_down_7[46]));
 BUFx2_ASAP7_75t_R output2602 (.A(net2602),
    .Y(io_outs_down_7[47]));
 BUFx2_ASAP7_75t_R output2603 (.A(net2603),
    .Y(io_outs_down_7[48]));
 BUFx2_ASAP7_75t_R output2604 (.A(net2604),
    .Y(io_outs_down_7[49]));
 BUFx2_ASAP7_75t_R output2605 (.A(net2605),
    .Y(io_outs_down_7[4]));
 BUFx2_ASAP7_75t_R output2606 (.A(net2606),
    .Y(io_outs_down_7[50]));
 BUFx2_ASAP7_75t_R output2607 (.A(net2607),
    .Y(io_outs_down_7[51]));
 BUFx2_ASAP7_75t_R output2608 (.A(net2608),
    .Y(io_outs_down_7[52]));
 BUFx2_ASAP7_75t_R output2609 (.A(net2609),
    .Y(io_outs_down_7[53]));
 BUFx2_ASAP7_75t_R output2610 (.A(net2610),
    .Y(io_outs_down_7[54]));
 BUFx2_ASAP7_75t_R output2611 (.A(net2611),
    .Y(io_outs_down_7[55]));
 BUFx2_ASAP7_75t_R output2612 (.A(net2612),
    .Y(io_outs_down_7[56]));
 BUFx2_ASAP7_75t_R output2613 (.A(net2613),
    .Y(io_outs_down_7[57]));
 BUFx2_ASAP7_75t_R output2614 (.A(net2614),
    .Y(io_outs_down_7[58]));
 BUFx2_ASAP7_75t_R output2615 (.A(net2615),
    .Y(io_outs_down_7[59]));
 BUFx2_ASAP7_75t_R output2616 (.A(net2616),
    .Y(io_outs_down_7[5]));
 BUFx2_ASAP7_75t_R output2617 (.A(net2617),
    .Y(io_outs_down_7[60]));
 BUFx2_ASAP7_75t_R output2618 (.A(net2618),
    .Y(io_outs_down_7[61]));
 BUFx2_ASAP7_75t_R output2619 (.A(net2619),
    .Y(io_outs_down_7[62]));
 BUFx2_ASAP7_75t_R output2620 (.A(net2620),
    .Y(io_outs_down_7[63]));
 BUFx2_ASAP7_75t_R output2621 (.A(net2621),
    .Y(io_outs_down_7[6]));
 BUFx2_ASAP7_75t_R output2622 (.A(net2622),
    .Y(io_outs_down_7[7]));
 BUFx2_ASAP7_75t_R output2623 (.A(net2623),
    .Y(io_outs_down_7[8]));
 BUFx2_ASAP7_75t_R output2624 (.A(net2624),
    .Y(io_outs_down_7[9]));
 BUFx2_ASAP7_75t_R output2625 (.A(net2625),
    .Y(io_outs_left_0[0]));
 BUFx2_ASAP7_75t_R output2626 (.A(net2626),
    .Y(io_outs_left_0[10]));
 BUFx2_ASAP7_75t_R output2627 (.A(net2627),
    .Y(io_outs_left_0[11]));
 BUFx2_ASAP7_75t_R output2628 (.A(net2628),
    .Y(io_outs_left_0[12]));
 BUFx2_ASAP7_75t_R output2629 (.A(net2629),
    .Y(io_outs_left_0[13]));
 BUFx2_ASAP7_75t_R output2630 (.A(net2630),
    .Y(io_outs_left_0[14]));
 BUFx2_ASAP7_75t_R output2631 (.A(net2631),
    .Y(io_outs_left_0[15]));
 BUFx2_ASAP7_75t_R output2632 (.A(net2632),
    .Y(io_outs_left_0[16]));
 BUFx2_ASAP7_75t_R output2633 (.A(net2633),
    .Y(io_outs_left_0[17]));
 BUFx2_ASAP7_75t_R output2634 (.A(net2634),
    .Y(io_outs_left_0[18]));
 BUFx2_ASAP7_75t_R output2635 (.A(net2635),
    .Y(io_outs_left_0[19]));
 BUFx2_ASAP7_75t_R output2636 (.A(net2636),
    .Y(io_outs_left_0[1]));
 BUFx2_ASAP7_75t_R output2637 (.A(net2637),
    .Y(io_outs_left_0[20]));
 BUFx2_ASAP7_75t_R output2638 (.A(net2638),
    .Y(io_outs_left_0[21]));
 BUFx2_ASAP7_75t_R output2639 (.A(net2639),
    .Y(io_outs_left_0[22]));
 BUFx2_ASAP7_75t_R output2640 (.A(net2640),
    .Y(io_outs_left_0[23]));
 BUFx2_ASAP7_75t_R output2641 (.A(net2641),
    .Y(io_outs_left_0[24]));
 BUFx2_ASAP7_75t_R output2642 (.A(net2642),
    .Y(io_outs_left_0[25]));
 BUFx2_ASAP7_75t_R output2643 (.A(net2643),
    .Y(io_outs_left_0[26]));
 BUFx2_ASAP7_75t_R output2644 (.A(net2644),
    .Y(io_outs_left_0[27]));
 BUFx2_ASAP7_75t_R output2645 (.A(net2645),
    .Y(io_outs_left_0[28]));
 BUFx2_ASAP7_75t_R output2646 (.A(net2646),
    .Y(io_outs_left_0[29]));
 BUFx2_ASAP7_75t_R output2647 (.A(net2647),
    .Y(io_outs_left_0[2]));
 BUFx2_ASAP7_75t_R output2648 (.A(net2648),
    .Y(io_outs_left_0[30]));
 BUFx2_ASAP7_75t_R output2649 (.A(net2649),
    .Y(io_outs_left_0[31]));
 BUFx2_ASAP7_75t_R output2650 (.A(net2650),
    .Y(io_outs_left_0[32]));
 BUFx2_ASAP7_75t_R output2651 (.A(net2651),
    .Y(io_outs_left_0[33]));
 BUFx2_ASAP7_75t_R output2652 (.A(net2652),
    .Y(io_outs_left_0[34]));
 BUFx2_ASAP7_75t_R output2653 (.A(net2653),
    .Y(io_outs_left_0[35]));
 BUFx2_ASAP7_75t_R output2654 (.A(net2654),
    .Y(io_outs_left_0[36]));
 BUFx2_ASAP7_75t_R output2655 (.A(net2655),
    .Y(io_outs_left_0[37]));
 BUFx2_ASAP7_75t_R output2656 (.A(net2656),
    .Y(io_outs_left_0[38]));
 BUFx2_ASAP7_75t_R output2657 (.A(net2657),
    .Y(io_outs_left_0[39]));
 BUFx2_ASAP7_75t_R output2658 (.A(net2658),
    .Y(io_outs_left_0[3]));
 BUFx2_ASAP7_75t_R output2659 (.A(net2659),
    .Y(io_outs_left_0[40]));
 BUFx2_ASAP7_75t_R output2660 (.A(net2660),
    .Y(io_outs_left_0[41]));
 BUFx2_ASAP7_75t_R output2661 (.A(net2661),
    .Y(io_outs_left_0[42]));
 BUFx2_ASAP7_75t_R output2662 (.A(net2662),
    .Y(io_outs_left_0[43]));
 BUFx2_ASAP7_75t_R output2663 (.A(net2663),
    .Y(io_outs_left_0[44]));
 BUFx2_ASAP7_75t_R output2664 (.A(net2664),
    .Y(io_outs_left_0[45]));
 BUFx2_ASAP7_75t_R output2665 (.A(net2665),
    .Y(io_outs_left_0[46]));
 BUFx2_ASAP7_75t_R output2666 (.A(net2666),
    .Y(io_outs_left_0[47]));
 BUFx2_ASAP7_75t_R output2667 (.A(net2667),
    .Y(io_outs_left_0[48]));
 BUFx2_ASAP7_75t_R output2668 (.A(net2668),
    .Y(io_outs_left_0[49]));
 BUFx2_ASAP7_75t_R output2669 (.A(net2669),
    .Y(io_outs_left_0[4]));
 BUFx2_ASAP7_75t_R output2670 (.A(net2670),
    .Y(io_outs_left_0[50]));
 BUFx2_ASAP7_75t_R output2671 (.A(net2671),
    .Y(io_outs_left_0[51]));
 BUFx2_ASAP7_75t_R output2672 (.A(net2672),
    .Y(io_outs_left_0[52]));
 BUFx2_ASAP7_75t_R output2673 (.A(net2673),
    .Y(io_outs_left_0[53]));
 BUFx2_ASAP7_75t_R output2674 (.A(net2674),
    .Y(io_outs_left_0[54]));
 BUFx2_ASAP7_75t_R output2675 (.A(net2675),
    .Y(io_outs_left_0[55]));
 BUFx2_ASAP7_75t_R output2676 (.A(net2676),
    .Y(io_outs_left_0[56]));
 BUFx2_ASAP7_75t_R output2677 (.A(net2677),
    .Y(io_outs_left_0[57]));
 BUFx2_ASAP7_75t_R output2678 (.A(net2678),
    .Y(io_outs_left_0[58]));
 BUFx2_ASAP7_75t_R output2679 (.A(net2679),
    .Y(io_outs_left_0[59]));
 BUFx2_ASAP7_75t_R output2680 (.A(net2680),
    .Y(io_outs_left_0[5]));
 BUFx2_ASAP7_75t_R output2681 (.A(net2681),
    .Y(io_outs_left_0[60]));
 BUFx2_ASAP7_75t_R output2682 (.A(net2682),
    .Y(io_outs_left_0[61]));
 BUFx2_ASAP7_75t_R output2683 (.A(net2683),
    .Y(io_outs_left_0[62]));
 BUFx2_ASAP7_75t_R output2684 (.A(net2684),
    .Y(io_outs_left_0[63]));
 BUFx2_ASAP7_75t_R output2685 (.A(net2685),
    .Y(io_outs_left_0[6]));
 BUFx2_ASAP7_75t_R output2686 (.A(net2686),
    .Y(io_outs_left_0[7]));
 BUFx2_ASAP7_75t_R output2687 (.A(net2687),
    .Y(io_outs_left_0[8]));
 BUFx2_ASAP7_75t_R output2688 (.A(net2688),
    .Y(io_outs_left_0[9]));
 BUFx2_ASAP7_75t_R output2689 (.A(net2689),
    .Y(io_outs_left_1[0]));
 BUFx2_ASAP7_75t_R output2690 (.A(net2690),
    .Y(io_outs_left_1[10]));
 BUFx2_ASAP7_75t_R output2691 (.A(net2691),
    .Y(io_outs_left_1[11]));
 BUFx2_ASAP7_75t_R output2692 (.A(net2692),
    .Y(io_outs_left_1[12]));
 BUFx2_ASAP7_75t_R output2693 (.A(net2693),
    .Y(io_outs_left_1[13]));
 BUFx2_ASAP7_75t_R output2694 (.A(net2694),
    .Y(io_outs_left_1[14]));
 BUFx2_ASAP7_75t_R output2695 (.A(net2695),
    .Y(io_outs_left_1[15]));
 BUFx2_ASAP7_75t_R output2696 (.A(net2696),
    .Y(io_outs_left_1[16]));
 BUFx2_ASAP7_75t_R output2697 (.A(net2697),
    .Y(io_outs_left_1[17]));
 BUFx2_ASAP7_75t_R output2698 (.A(net2698),
    .Y(io_outs_left_1[18]));
 BUFx2_ASAP7_75t_R output2699 (.A(net2699),
    .Y(io_outs_left_1[19]));
 BUFx2_ASAP7_75t_R output2700 (.A(net2700),
    .Y(io_outs_left_1[1]));
 BUFx2_ASAP7_75t_R output2701 (.A(net2701),
    .Y(io_outs_left_1[20]));
 BUFx2_ASAP7_75t_R output2702 (.A(net2702),
    .Y(io_outs_left_1[21]));
 BUFx2_ASAP7_75t_R output2703 (.A(net2703),
    .Y(io_outs_left_1[22]));
 BUFx2_ASAP7_75t_R output2704 (.A(net2704),
    .Y(io_outs_left_1[23]));
 BUFx2_ASAP7_75t_R output2705 (.A(net2705),
    .Y(io_outs_left_1[24]));
 BUFx2_ASAP7_75t_R output2706 (.A(net2706),
    .Y(io_outs_left_1[25]));
 BUFx2_ASAP7_75t_R output2707 (.A(net2707),
    .Y(io_outs_left_1[26]));
 BUFx2_ASAP7_75t_R output2708 (.A(net2708),
    .Y(io_outs_left_1[27]));
 BUFx2_ASAP7_75t_R output2709 (.A(net2709),
    .Y(io_outs_left_1[28]));
 BUFx2_ASAP7_75t_R output2710 (.A(net2710),
    .Y(io_outs_left_1[29]));
 BUFx2_ASAP7_75t_R output2711 (.A(net2711),
    .Y(io_outs_left_1[2]));
 BUFx2_ASAP7_75t_R output2712 (.A(net2712),
    .Y(io_outs_left_1[30]));
 BUFx2_ASAP7_75t_R output2713 (.A(net2713),
    .Y(io_outs_left_1[31]));
 BUFx2_ASAP7_75t_R output2714 (.A(net2714),
    .Y(io_outs_left_1[32]));
 BUFx2_ASAP7_75t_R output2715 (.A(net2715),
    .Y(io_outs_left_1[33]));
 BUFx2_ASAP7_75t_R output2716 (.A(net2716),
    .Y(io_outs_left_1[34]));
 BUFx2_ASAP7_75t_R output2717 (.A(net2717),
    .Y(io_outs_left_1[35]));
 BUFx2_ASAP7_75t_R output2718 (.A(net2718),
    .Y(io_outs_left_1[36]));
 BUFx2_ASAP7_75t_R output2719 (.A(net2719),
    .Y(io_outs_left_1[37]));
 BUFx2_ASAP7_75t_R output2720 (.A(net2720),
    .Y(io_outs_left_1[38]));
 BUFx2_ASAP7_75t_R output2721 (.A(net2721),
    .Y(io_outs_left_1[39]));
 BUFx2_ASAP7_75t_R output2722 (.A(net2722),
    .Y(io_outs_left_1[3]));
 BUFx2_ASAP7_75t_R output2723 (.A(net2723),
    .Y(io_outs_left_1[40]));
 BUFx2_ASAP7_75t_R output2724 (.A(net2724),
    .Y(io_outs_left_1[41]));
 BUFx2_ASAP7_75t_R output2725 (.A(net2725),
    .Y(io_outs_left_1[42]));
 BUFx2_ASAP7_75t_R output2726 (.A(net2726),
    .Y(io_outs_left_1[43]));
 BUFx2_ASAP7_75t_R output2727 (.A(net2727),
    .Y(io_outs_left_1[44]));
 BUFx2_ASAP7_75t_R output2728 (.A(net2728),
    .Y(io_outs_left_1[45]));
 BUFx2_ASAP7_75t_R output2729 (.A(net2729),
    .Y(io_outs_left_1[46]));
 BUFx2_ASAP7_75t_R output2730 (.A(net2730),
    .Y(io_outs_left_1[47]));
 BUFx2_ASAP7_75t_R output2731 (.A(net2731),
    .Y(io_outs_left_1[48]));
 BUFx2_ASAP7_75t_R output2732 (.A(net2732),
    .Y(io_outs_left_1[49]));
 BUFx2_ASAP7_75t_R output2733 (.A(net2733),
    .Y(io_outs_left_1[4]));
 BUFx2_ASAP7_75t_R output2734 (.A(net2734),
    .Y(io_outs_left_1[50]));
 BUFx2_ASAP7_75t_R output2735 (.A(net2735),
    .Y(io_outs_left_1[51]));
 BUFx2_ASAP7_75t_R output2736 (.A(net2736),
    .Y(io_outs_left_1[52]));
 BUFx2_ASAP7_75t_R output2737 (.A(net2737),
    .Y(io_outs_left_1[53]));
 BUFx2_ASAP7_75t_R output2738 (.A(net2738),
    .Y(io_outs_left_1[54]));
 BUFx2_ASAP7_75t_R output2739 (.A(net2739),
    .Y(io_outs_left_1[55]));
 BUFx2_ASAP7_75t_R output2740 (.A(net2740),
    .Y(io_outs_left_1[56]));
 BUFx2_ASAP7_75t_R output2741 (.A(net2741),
    .Y(io_outs_left_1[57]));
 BUFx2_ASAP7_75t_R output2742 (.A(net2742),
    .Y(io_outs_left_1[58]));
 BUFx2_ASAP7_75t_R output2743 (.A(net2743),
    .Y(io_outs_left_1[59]));
 BUFx2_ASAP7_75t_R output2744 (.A(net2744),
    .Y(io_outs_left_1[5]));
 BUFx2_ASAP7_75t_R output2745 (.A(net2745),
    .Y(io_outs_left_1[60]));
 BUFx2_ASAP7_75t_R output2746 (.A(net2746),
    .Y(io_outs_left_1[61]));
 BUFx2_ASAP7_75t_R output2747 (.A(net2747),
    .Y(io_outs_left_1[62]));
 BUFx2_ASAP7_75t_R output2748 (.A(net2748),
    .Y(io_outs_left_1[63]));
 BUFx2_ASAP7_75t_R output2749 (.A(net2749),
    .Y(io_outs_left_1[6]));
 BUFx2_ASAP7_75t_R output2750 (.A(net2750),
    .Y(io_outs_left_1[7]));
 BUFx2_ASAP7_75t_R output2751 (.A(net2751),
    .Y(io_outs_left_1[8]));
 BUFx2_ASAP7_75t_R output2752 (.A(net2752),
    .Y(io_outs_left_1[9]));
 BUFx2_ASAP7_75t_R output2753 (.A(net2753),
    .Y(io_outs_left_2[0]));
 BUFx2_ASAP7_75t_R output2754 (.A(net2754),
    .Y(io_outs_left_2[10]));
 BUFx2_ASAP7_75t_R output2755 (.A(net2755),
    .Y(io_outs_left_2[11]));
 BUFx2_ASAP7_75t_R output2756 (.A(net2756),
    .Y(io_outs_left_2[12]));
 BUFx2_ASAP7_75t_R output2757 (.A(net2757),
    .Y(io_outs_left_2[13]));
 BUFx2_ASAP7_75t_R output2758 (.A(net2758),
    .Y(io_outs_left_2[14]));
 BUFx2_ASAP7_75t_R output2759 (.A(net2759),
    .Y(io_outs_left_2[15]));
 BUFx2_ASAP7_75t_R output2760 (.A(net2760),
    .Y(io_outs_left_2[16]));
 BUFx2_ASAP7_75t_R output2761 (.A(net2761),
    .Y(io_outs_left_2[17]));
 BUFx2_ASAP7_75t_R output2762 (.A(net2762),
    .Y(io_outs_left_2[18]));
 BUFx2_ASAP7_75t_R output2763 (.A(net2763),
    .Y(io_outs_left_2[19]));
 BUFx2_ASAP7_75t_R output2764 (.A(net2764),
    .Y(io_outs_left_2[1]));
 BUFx2_ASAP7_75t_R output2765 (.A(net2765),
    .Y(io_outs_left_2[20]));
 BUFx2_ASAP7_75t_R output2766 (.A(net2766),
    .Y(io_outs_left_2[21]));
 BUFx2_ASAP7_75t_R output2767 (.A(net2767),
    .Y(io_outs_left_2[22]));
 BUFx2_ASAP7_75t_R output2768 (.A(net2768),
    .Y(io_outs_left_2[23]));
 BUFx2_ASAP7_75t_R output2769 (.A(net2769),
    .Y(io_outs_left_2[24]));
 BUFx2_ASAP7_75t_R output2770 (.A(net2770),
    .Y(io_outs_left_2[25]));
 BUFx2_ASAP7_75t_R output2771 (.A(net2771),
    .Y(io_outs_left_2[26]));
 BUFx2_ASAP7_75t_R output2772 (.A(net2772),
    .Y(io_outs_left_2[27]));
 BUFx2_ASAP7_75t_R output2773 (.A(net2773),
    .Y(io_outs_left_2[28]));
 BUFx2_ASAP7_75t_R output2774 (.A(net2774),
    .Y(io_outs_left_2[29]));
 BUFx2_ASAP7_75t_R output2775 (.A(net2775),
    .Y(io_outs_left_2[2]));
 BUFx2_ASAP7_75t_R output2776 (.A(net2776),
    .Y(io_outs_left_2[30]));
 BUFx2_ASAP7_75t_R output2777 (.A(net2777),
    .Y(io_outs_left_2[31]));
 BUFx2_ASAP7_75t_R output2778 (.A(net2778),
    .Y(io_outs_left_2[32]));
 BUFx2_ASAP7_75t_R output2779 (.A(net2779),
    .Y(io_outs_left_2[33]));
 BUFx2_ASAP7_75t_R output2780 (.A(net2780),
    .Y(io_outs_left_2[34]));
 BUFx2_ASAP7_75t_R output2781 (.A(net2781),
    .Y(io_outs_left_2[35]));
 BUFx2_ASAP7_75t_R output2782 (.A(net2782),
    .Y(io_outs_left_2[36]));
 BUFx2_ASAP7_75t_R output2783 (.A(net2783),
    .Y(io_outs_left_2[37]));
 BUFx2_ASAP7_75t_R output2784 (.A(net2784),
    .Y(io_outs_left_2[38]));
 BUFx2_ASAP7_75t_R output2785 (.A(net2785),
    .Y(io_outs_left_2[39]));
 BUFx2_ASAP7_75t_R output2786 (.A(net2786),
    .Y(io_outs_left_2[3]));
 BUFx2_ASAP7_75t_R output2787 (.A(net2787),
    .Y(io_outs_left_2[40]));
 BUFx2_ASAP7_75t_R output2788 (.A(net2788),
    .Y(io_outs_left_2[41]));
 BUFx2_ASAP7_75t_R output2789 (.A(net2789),
    .Y(io_outs_left_2[42]));
 BUFx2_ASAP7_75t_R output2790 (.A(net2790),
    .Y(io_outs_left_2[43]));
 BUFx2_ASAP7_75t_R output2791 (.A(net2791),
    .Y(io_outs_left_2[44]));
 BUFx2_ASAP7_75t_R output2792 (.A(net2792),
    .Y(io_outs_left_2[45]));
 BUFx2_ASAP7_75t_R output2793 (.A(net2793),
    .Y(io_outs_left_2[46]));
 BUFx2_ASAP7_75t_R output2794 (.A(net2794),
    .Y(io_outs_left_2[47]));
 BUFx2_ASAP7_75t_R output2795 (.A(net2795),
    .Y(io_outs_left_2[48]));
 BUFx2_ASAP7_75t_R output2796 (.A(net2796),
    .Y(io_outs_left_2[49]));
 BUFx2_ASAP7_75t_R output2797 (.A(net2797),
    .Y(io_outs_left_2[4]));
 BUFx2_ASAP7_75t_R output2798 (.A(net2798),
    .Y(io_outs_left_2[50]));
 BUFx2_ASAP7_75t_R output2799 (.A(net2799),
    .Y(io_outs_left_2[51]));
 BUFx2_ASAP7_75t_R output2800 (.A(net2800),
    .Y(io_outs_left_2[52]));
 BUFx2_ASAP7_75t_R output2801 (.A(net2801),
    .Y(io_outs_left_2[53]));
 BUFx2_ASAP7_75t_R output2802 (.A(net2802),
    .Y(io_outs_left_2[54]));
 BUFx2_ASAP7_75t_R output2803 (.A(net2803),
    .Y(io_outs_left_2[55]));
 BUFx2_ASAP7_75t_R output2804 (.A(net2804),
    .Y(io_outs_left_2[56]));
 BUFx2_ASAP7_75t_R output2805 (.A(net2805),
    .Y(io_outs_left_2[57]));
 BUFx2_ASAP7_75t_R output2806 (.A(net2806),
    .Y(io_outs_left_2[58]));
 BUFx2_ASAP7_75t_R output2807 (.A(net2807),
    .Y(io_outs_left_2[59]));
 BUFx2_ASAP7_75t_R output2808 (.A(net2808),
    .Y(io_outs_left_2[5]));
 BUFx2_ASAP7_75t_R output2809 (.A(net2809),
    .Y(io_outs_left_2[60]));
 BUFx2_ASAP7_75t_R output2810 (.A(net2810),
    .Y(io_outs_left_2[61]));
 BUFx2_ASAP7_75t_R output2811 (.A(net2811),
    .Y(io_outs_left_2[62]));
 BUFx2_ASAP7_75t_R output2812 (.A(net2812),
    .Y(io_outs_left_2[63]));
 BUFx2_ASAP7_75t_R output2813 (.A(net2813),
    .Y(io_outs_left_2[6]));
 BUFx2_ASAP7_75t_R output2814 (.A(net2814),
    .Y(io_outs_left_2[7]));
 BUFx2_ASAP7_75t_R output2815 (.A(net2815),
    .Y(io_outs_left_2[8]));
 BUFx2_ASAP7_75t_R output2816 (.A(net2816),
    .Y(io_outs_left_2[9]));
 BUFx2_ASAP7_75t_R output2817 (.A(net2817),
    .Y(io_outs_left_3[0]));
 BUFx2_ASAP7_75t_R output2818 (.A(net2818),
    .Y(io_outs_left_3[10]));
 BUFx2_ASAP7_75t_R output2819 (.A(net2819),
    .Y(io_outs_left_3[11]));
 BUFx2_ASAP7_75t_R output2820 (.A(net2820),
    .Y(io_outs_left_3[12]));
 BUFx2_ASAP7_75t_R output2821 (.A(net2821),
    .Y(io_outs_left_3[13]));
 BUFx2_ASAP7_75t_R output2822 (.A(net2822),
    .Y(io_outs_left_3[14]));
 BUFx2_ASAP7_75t_R output2823 (.A(net2823),
    .Y(io_outs_left_3[15]));
 BUFx2_ASAP7_75t_R output2824 (.A(net2824),
    .Y(io_outs_left_3[16]));
 BUFx2_ASAP7_75t_R output2825 (.A(net2825),
    .Y(io_outs_left_3[17]));
 BUFx2_ASAP7_75t_R output2826 (.A(net2826),
    .Y(io_outs_left_3[18]));
 BUFx2_ASAP7_75t_R output2827 (.A(net2827),
    .Y(io_outs_left_3[19]));
 BUFx2_ASAP7_75t_R output2828 (.A(net2828),
    .Y(io_outs_left_3[1]));
 BUFx2_ASAP7_75t_R output2829 (.A(net2829),
    .Y(io_outs_left_3[20]));
 BUFx2_ASAP7_75t_R output2830 (.A(net2830),
    .Y(io_outs_left_3[21]));
 BUFx2_ASAP7_75t_R output2831 (.A(net2831),
    .Y(io_outs_left_3[22]));
 BUFx2_ASAP7_75t_R output2832 (.A(net2832),
    .Y(io_outs_left_3[23]));
 BUFx2_ASAP7_75t_R output2833 (.A(net2833),
    .Y(io_outs_left_3[24]));
 BUFx2_ASAP7_75t_R output2834 (.A(net2834),
    .Y(io_outs_left_3[25]));
 BUFx2_ASAP7_75t_R output2835 (.A(net2835),
    .Y(io_outs_left_3[26]));
 BUFx2_ASAP7_75t_R output2836 (.A(net2836),
    .Y(io_outs_left_3[27]));
 BUFx2_ASAP7_75t_R output2837 (.A(net2837),
    .Y(io_outs_left_3[28]));
 BUFx2_ASAP7_75t_R output2838 (.A(net2838),
    .Y(io_outs_left_3[29]));
 BUFx2_ASAP7_75t_R output2839 (.A(net2839),
    .Y(io_outs_left_3[2]));
 BUFx2_ASAP7_75t_R output2840 (.A(net2840),
    .Y(io_outs_left_3[30]));
 BUFx2_ASAP7_75t_R output2841 (.A(net2841),
    .Y(io_outs_left_3[31]));
 BUFx2_ASAP7_75t_R output2842 (.A(net2842),
    .Y(io_outs_left_3[32]));
 BUFx2_ASAP7_75t_R output2843 (.A(net2843),
    .Y(io_outs_left_3[33]));
 BUFx2_ASAP7_75t_R output2844 (.A(net2844),
    .Y(io_outs_left_3[34]));
 BUFx2_ASAP7_75t_R output2845 (.A(net2845),
    .Y(io_outs_left_3[35]));
 BUFx2_ASAP7_75t_R output2846 (.A(net2846),
    .Y(io_outs_left_3[36]));
 BUFx2_ASAP7_75t_R output2847 (.A(net2847),
    .Y(io_outs_left_3[37]));
 BUFx2_ASAP7_75t_R output2848 (.A(net2848),
    .Y(io_outs_left_3[38]));
 BUFx2_ASAP7_75t_R output2849 (.A(net2849),
    .Y(io_outs_left_3[39]));
 BUFx2_ASAP7_75t_R output2850 (.A(net2850),
    .Y(io_outs_left_3[3]));
 BUFx2_ASAP7_75t_R output2851 (.A(net2851),
    .Y(io_outs_left_3[40]));
 BUFx2_ASAP7_75t_R output2852 (.A(net2852),
    .Y(io_outs_left_3[41]));
 BUFx2_ASAP7_75t_R output2853 (.A(net2853),
    .Y(io_outs_left_3[42]));
 BUFx2_ASAP7_75t_R output2854 (.A(net2854),
    .Y(io_outs_left_3[43]));
 BUFx2_ASAP7_75t_R output2855 (.A(net2855),
    .Y(io_outs_left_3[44]));
 BUFx2_ASAP7_75t_R output2856 (.A(net2856),
    .Y(io_outs_left_3[45]));
 BUFx2_ASAP7_75t_R output2857 (.A(net2857),
    .Y(io_outs_left_3[46]));
 BUFx2_ASAP7_75t_R output2858 (.A(net2858),
    .Y(io_outs_left_3[47]));
 BUFx2_ASAP7_75t_R output2859 (.A(net2859),
    .Y(io_outs_left_3[48]));
 BUFx2_ASAP7_75t_R output2860 (.A(net2860),
    .Y(io_outs_left_3[49]));
 BUFx2_ASAP7_75t_R output2861 (.A(net2861),
    .Y(io_outs_left_3[4]));
 BUFx2_ASAP7_75t_R output2862 (.A(net2862),
    .Y(io_outs_left_3[50]));
 BUFx2_ASAP7_75t_R output2863 (.A(net2863),
    .Y(io_outs_left_3[51]));
 BUFx2_ASAP7_75t_R output2864 (.A(net2864),
    .Y(io_outs_left_3[52]));
 BUFx2_ASAP7_75t_R output2865 (.A(net2865),
    .Y(io_outs_left_3[53]));
 BUFx2_ASAP7_75t_R output2866 (.A(net2866),
    .Y(io_outs_left_3[54]));
 BUFx2_ASAP7_75t_R output2867 (.A(net2867),
    .Y(io_outs_left_3[55]));
 BUFx2_ASAP7_75t_R output2868 (.A(net2868),
    .Y(io_outs_left_3[56]));
 BUFx2_ASAP7_75t_R output2869 (.A(net2869),
    .Y(io_outs_left_3[57]));
 BUFx2_ASAP7_75t_R output2870 (.A(net2870),
    .Y(io_outs_left_3[58]));
 BUFx2_ASAP7_75t_R output2871 (.A(net2871),
    .Y(io_outs_left_3[59]));
 BUFx2_ASAP7_75t_R output2872 (.A(net2872),
    .Y(io_outs_left_3[5]));
 BUFx2_ASAP7_75t_R output2873 (.A(net2873),
    .Y(io_outs_left_3[60]));
 BUFx2_ASAP7_75t_R output2874 (.A(net2874),
    .Y(io_outs_left_3[61]));
 BUFx2_ASAP7_75t_R output2875 (.A(net2875),
    .Y(io_outs_left_3[62]));
 BUFx2_ASAP7_75t_R output2876 (.A(net2876),
    .Y(io_outs_left_3[63]));
 BUFx2_ASAP7_75t_R output2877 (.A(net2877),
    .Y(io_outs_left_3[6]));
 BUFx2_ASAP7_75t_R output2878 (.A(net2878),
    .Y(io_outs_left_3[7]));
 BUFx2_ASAP7_75t_R output2879 (.A(net2879),
    .Y(io_outs_left_3[8]));
 BUFx2_ASAP7_75t_R output2880 (.A(net2880),
    .Y(io_outs_left_3[9]));
 BUFx2_ASAP7_75t_R output2881 (.A(net2881),
    .Y(io_outs_left_4[0]));
 BUFx2_ASAP7_75t_R output2882 (.A(net2882),
    .Y(io_outs_left_4[10]));
 BUFx2_ASAP7_75t_R output2883 (.A(net2883),
    .Y(io_outs_left_4[11]));
 BUFx2_ASAP7_75t_R output2884 (.A(net2884),
    .Y(io_outs_left_4[12]));
 BUFx2_ASAP7_75t_R output2885 (.A(net2885),
    .Y(io_outs_left_4[13]));
 BUFx2_ASAP7_75t_R output2886 (.A(net2886),
    .Y(io_outs_left_4[14]));
 BUFx2_ASAP7_75t_R output2887 (.A(net2887),
    .Y(io_outs_left_4[15]));
 BUFx2_ASAP7_75t_R output2888 (.A(net2888),
    .Y(io_outs_left_4[16]));
 BUFx2_ASAP7_75t_R output2889 (.A(net2889),
    .Y(io_outs_left_4[17]));
 BUFx2_ASAP7_75t_R output2890 (.A(net2890),
    .Y(io_outs_left_4[18]));
 BUFx2_ASAP7_75t_R output2891 (.A(net2891),
    .Y(io_outs_left_4[19]));
 BUFx2_ASAP7_75t_R output2892 (.A(net2892),
    .Y(io_outs_left_4[1]));
 BUFx2_ASAP7_75t_R output2893 (.A(net2893),
    .Y(io_outs_left_4[20]));
 BUFx2_ASAP7_75t_R output2894 (.A(net2894),
    .Y(io_outs_left_4[21]));
 BUFx2_ASAP7_75t_R output2895 (.A(net2895),
    .Y(io_outs_left_4[22]));
 BUFx2_ASAP7_75t_R output2896 (.A(net2896),
    .Y(io_outs_left_4[23]));
 BUFx2_ASAP7_75t_R output2897 (.A(net2897),
    .Y(io_outs_left_4[24]));
 BUFx2_ASAP7_75t_R output2898 (.A(net2898),
    .Y(io_outs_left_4[25]));
 BUFx2_ASAP7_75t_R output2899 (.A(net2899),
    .Y(io_outs_left_4[26]));
 BUFx2_ASAP7_75t_R output2900 (.A(net2900),
    .Y(io_outs_left_4[27]));
 BUFx2_ASAP7_75t_R output2901 (.A(net2901),
    .Y(io_outs_left_4[28]));
 BUFx2_ASAP7_75t_R output2902 (.A(net2902),
    .Y(io_outs_left_4[29]));
 BUFx2_ASAP7_75t_R output2903 (.A(net2903),
    .Y(io_outs_left_4[2]));
 BUFx2_ASAP7_75t_R output2904 (.A(net2904),
    .Y(io_outs_left_4[30]));
 BUFx2_ASAP7_75t_R output2905 (.A(net2905),
    .Y(io_outs_left_4[31]));
 BUFx2_ASAP7_75t_R output2906 (.A(net2906),
    .Y(io_outs_left_4[32]));
 BUFx2_ASAP7_75t_R output2907 (.A(net2907),
    .Y(io_outs_left_4[33]));
 BUFx2_ASAP7_75t_R output2908 (.A(net2908),
    .Y(io_outs_left_4[34]));
 BUFx2_ASAP7_75t_R output2909 (.A(net2909),
    .Y(io_outs_left_4[35]));
 BUFx2_ASAP7_75t_R output2910 (.A(net2910),
    .Y(io_outs_left_4[36]));
 BUFx2_ASAP7_75t_R output2911 (.A(net2911),
    .Y(io_outs_left_4[37]));
 BUFx2_ASAP7_75t_R output2912 (.A(net2912),
    .Y(io_outs_left_4[38]));
 BUFx2_ASAP7_75t_R output2913 (.A(net2913),
    .Y(io_outs_left_4[39]));
 BUFx2_ASAP7_75t_R output2914 (.A(net2914),
    .Y(io_outs_left_4[3]));
 BUFx2_ASAP7_75t_R output2915 (.A(net2915),
    .Y(io_outs_left_4[40]));
 BUFx2_ASAP7_75t_R output2916 (.A(net2916),
    .Y(io_outs_left_4[41]));
 BUFx2_ASAP7_75t_R output2917 (.A(net2917),
    .Y(io_outs_left_4[42]));
 BUFx2_ASAP7_75t_R output2918 (.A(net2918),
    .Y(io_outs_left_4[43]));
 BUFx2_ASAP7_75t_R output2919 (.A(net2919),
    .Y(io_outs_left_4[44]));
 BUFx2_ASAP7_75t_R output2920 (.A(net2920),
    .Y(io_outs_left_4[45]));
 BUFx2_ASAP7_75t_R output2921 (.A(net2921),
    .Y(io_outs_left_4[46]));
 BUFx2_ASAP7_75t_R output2922 (.A(net2922),
    .Y(io_outs_left_4[47]));
 BUFx2_ASAP7_75t_R output2923 (.A(net2923),
    .Y(io_outs_left_4[48]));
 BUFx2_ASAP7_75t_R output2924 (.A(net2924),
    .Y(io_outs_left_4[49]));
 BUFx2_ASAP7_75t_R output2925 (.A(net2925),
    .Y(io_outs_left_4[4]));
 BUFx2_ASAP7_75t_R output2926 (.A(net2926),
    .Y(io_outs_left_4[50]));
 BUFx2_ASAP7_75t_R output2927 (.A(net2927),
    .Y(io_outs_left_4[51]));
 BUFx2_ASAP7_75t_R output2928 (.A(net2928),
    .Y(io_outs_left_4[52]));
 BUFx2_ASAP7_75t_R output2929 (.A(net2929),
    .Y(io_outs_left_4[53]));
 BUFx2_ASAP7_75t_R output2930 (.A(net2930),
    .Y(io_outs_left_4[54]));
 BUFx2_ASAP7_75t_R output2931 (.A(net2931),
    .Y(io_outs_left_4[55]));
 BUFx2_ASAP7_75t_R output2932 (.A(net2932),
    .Y(io_outs_left_4[56]));
 BUFx2_ASAP7_75t_R output2933 (.A(net2933),
    .Y(io_outs_left_4[57]));
 BUFx2_ASAP7_75t_R output2934 (.A(net2934),
    .Y(io_outs_left_4[58]));
 BUFx2_ASAP7_75t_R output2935 (.A(net2935),
    .Y(io_outs_left_4[59]));
 BUFx2_ASAP7_75t_R output2936 (.A(net2936),
    .Y(io_outs_left_4[5]));
 BUFx2_ASAP7_75t_R output2937 (.A(net2937),
    .Y(io_outs_left_4[60]));
 BUFx2_ASAP7_75t_R output2938 (.A(net2938),
    .Y(io_outs_left_4[61]));
 BUFx2_ASAP7_75t_R output2939 (.A(net2939),
    .Y(io_outs_left_4[62]));
 BUFx2_ASAP7_75t_R output2940 (.A(net2940),
    .Y(io_outs_left_4[63]));
 BUFx2_ASAP7_75t_R output2941 (.A(net2941),
    .Y(io_outs_left_4[6]));
 BUFx2_ASAP7_75t_R output2942 (.A(net2942),
    .Y(io_outs_left_4[7]));
 BUFx2_ASAP7_75t_R output2943 (.A(net2943),
    .Y(io_outs_left_4[8]));
 BUFx2_ASAP7_75t_R output2944 (.A(net2944),
    .Y(io_outs_left_4[9]));
 BUFx2_ASAP7_75t_R output2945 (.A(net2945),
    .Y(io_outs_left_5[0]));
 BUFx2_ASAP7_75t_R output2946 (.A(net2946),
    .Y(io_outs_left_5[10]));
 BUFx2_ASAP7_75t_R output2947 (.A(net2947),
    .Y(io_outs_left_5[11]));
 BUFx2_ASAP7_75t_R output2948 (.A(net2948),
    .Y(io_outs_left_5[12]));
 BUFx2_ASAP7_75t_R output2949 (.A(net2949),
    .Y(io_outs_left_5[13]));
 BUFx2_ASAP7_75t_R output2950 (.A(net2950),
    .Y(io_outs_left_5[14]));
 BUFx2_ASAP7_75t_R output2951 (.A(net2951),
    .Y(io_outs_left_5[15]));
 BUFx2_ASAP7_75t_R output2952 (.A(net2952),
    .Y(io_outs_left_5[16]));
 BUFx2_ASAP7_75t_R output2953 (.A(net2953),
    .Y(io_outs_left_5[17]));
 BUFx2_ASAP7_75t_R output2954 (.A(net2954),
    .Y(io_outs_left_5[18]));
 BUFx2_ASAP7_75t_R output2955 (.A(net2955),
    .Y(io_outs_left_5[19]));
 BUFx2_ASAP7_75t_R output2956 (.A(net2956),
    .Y(io_outs_left_5[1]));
 BUFx2_ASAP7_75t_R output2957 (.A(net2957),
    .Y(io_outs_left_5[20]));
 BUFx2_ASAP7_75t_R output2958 (.A(net2958),
    .Y(io_outs_left_5[21]));
 BUFx2_ASAP7_75t_R output2959 (.A(net2959),
    .Y(io_outs_left_5[22]));
 BUFx2_ASAP7_75t_R output2960 (.A(net2960),
    .Y(io_outs_left_5[23]));
 BUFx2_ASAP7_75t_R output2961 (.A(net2961),
    .Y(io_outs_left_5[24]));
 BUFx2_ASAP7_75t_R output2962 (.A(net2962),
    .Y(io_outs_left_5[25]));
 BUFx2_ASAP7_75t_R output2963 (.A(net2963),
    .Y(io_outs_left_5[26]));
 BUFx2_ASAP7_75t_R output2964 (.A(net2964),
    .Y(io_outs_left_5[27]));
 BUFx2_ASAP7_75t_R output2965 (.A(net2965),
    .Y(io_outs_left_5[28]));
 BUFx2_ASAP7_75t_R output2966 (.A(net2966),
    .Y(io_outs_left_5[29]));
 BUFx2_ASAP7_75t_R output2967 (.A(net2967),
    .Y(io_outs_left_5[2]));
 BUFx2_ASAP7_75t_R output2968 (.A(net2968),
    .Y(io_outs_left_5[30]));
 BUFx2_ASAP7_75t_R output2969 (.A(net2969),
    .Y(io_outs_left_5[31]));
 BUFx2_ASAP7_75t_R output2970 (.A(net2970),
    .Y(io_outs_left_5[32]));
 BUFx2_ASAP7_75t_R output2971 (.A(net2971),
    .Y(io_outs_left_5[33]));
 BUFx2_ASAP7_75t_R output2972 (.A(net2972),
    .Y(io_outs_left_5[34]));
 BUFx2_ASAP7_75t_R output2973 (.A(net2973),
    .Y(io_outs_left_5[35]));
 BUFx2_ASAP7_75t_R output2974 (.A(net2974),
    .Y(io_outs_left_5[36]));
 BUFx2_ASAP7_75t_R output2975 (.A(net2975),
    .Y(io_outs_left_5[37]));
 BUFx2_ASAP7_75t_R output2976 (.A(net2976),
    .Y(io_outs_left_5[38]));
 BUFx2_ASAP7_75t_R output2977 (.A(net2977),
    .Y(io_outs_left_5[39]));
 BUFx2_ASAP7_75t_R output2978 (.A(net2978),
    .Y(io_outs_left_5[3]));
 BUFx2_ASAP7_75t_R output2979 (.A(net2979),
    .Y(io_outs_left_5[40]));
 BUFx2_ASAP7_75t_R output2980 (.A(net2980),
    .Y(io_outs_left_5[41]));
 BUFx2_ASAP7_75t_R output2981 (.A(net2981),
    .Y(io_outs_left_5[42]));
 BUFx2_ASAP7_75t_R output2982 (.A(net2982),
    .Y(io_outs_left_5[43]));
 BUFx2_ASAP7_75t_R output2983 (.A(net2983),
    .Y(io_outs_left_5[44]));
 BUFx2_ASAP7_75t_R output2984 (.A(net2984),
    .Y(io_outs_left_5[45]));
 BUFx2_ASAP7_75t_R output2985 (.A(net2985),
    .Y(io_outs_left_5[46]));
 BUFx2_ASAP7_75t_R output2986 (.A(net2986),
    .Y(io_outs_left_5[47]));
 BUFx2_ASAP7_75t_R output2987 (.A(net2987),
    .Y(io_outs_left_5[48]));
 BUFx2_ASAP7_75t_R output2988 (.A(net2988),
    .Y(io_outs_left_5[49]));
 BUFx2_ASAP7_75t_R output2989 (.A(net2989),
    .Y(io_outs_left_5[4]));
 BUFx2_ASAP7_75t_R output2990 (.A(net2990),
    .Y(io_outs_left_5[50]));
 BUFx2_ASAP7_75t_R output2991 (.A(net2991),
    .Y(io_outs_left_5[51]));
 BUFx2_ASAP7_75t_R output2992 (.A(net2992),
    .Y(io_outs_left_5[52]));
 BUFx2_ASAP7_75t_R output2993 (.A(net2993),
    .Y(io_outs_left_5[53]));
 BUFx2_ASAP7_75t_R output2994 (.A(net2994),
    .Y(io_outs_left_5[54]));
 BUFx2_ASAP7_75t_R output2995 (.A(net2995),
    .Y(io_outs_left_5[55]));
 BUFx2_ASAP7_75t_R output2996 (.A(net2996),
    .Y(io_outs_left_5[56]));
 BUFx2_ASAP7_75t_R output2997 (.A(net2997),
    .Y(io_outs_left_5[57]));
 BUFx2_ASAP7_75t_R output2998 (.A(net2998),
    .Y(io_outs_left_5[58]));
 BUFx2_ASAP7_75t_R output2999 (.A(net2999),
    .Y(io_outs_left_5[59]));
 BUFx2_ASAP7_75t_R output3000 (.A(net3000),
    .Y(io_outs_left_5[5]));
 BUFx2_ASAP7_75t_R output3001 (.A(net3001),
    .Y(io_outs_left_5[60]));
 BUFx2_ASAP7_75t_R output3002 (.A(net3002),
    .Y(io_outs_left_5[61]));
 BUFx2_ASAP7_75t_R output3003 (.A(net3003),
    .Y(io_outs_left_5[62]));
 BUFx2_ASAP7_75t_R output3004 (.A(net3004),
    .Y(io_outs_left_5[63]));
 BUFx2_ASAP7_75t_R output3005 (.A(net3005),
    .Y(io_outs_left_5[6]));
 BUFx2_ASAP7_75t_R output3006 (.A(net3006),
    .Y(io_outs_left_5[7]));
 BUFx2_ASAP7_75t_R output3007 (.A(net3007),
    .Y(io_outs_left_5[8]));
 BUFx2_ASAP7_75t_R output3008 (.A(net3008),
    .Y(io_outs_left_5[9]));
 BUFx2_ASAP7_75t_R output3009 (.A(net3009),
    .Y(io_outs_left_6[0]));
 BUFx2_ASAP7_75t_R output3010 (.A(net3010),
    .Y(io_outs_left_6[10]));
 BUFx2_ASAP7_75t_R output3011 (.A(net3011),
    .Y(io_outs_left_6[11]));
 BUFx2_ASAP7_75t_R output3012 (.A(net3012),
    .Y(io_outs_left_6[12]));
 BUFx2_ASAP7_75t_R output3013 (.A(net3013),
    .Y(io_outs_left_6[13]));
 BUFx2_ASAP7_75t_R output3014 (.A(net3014),
    .Y(io_outs_left_6[14]));
 BUFx2_ASAP7_75t_R output3015 (.A(net3015),
    .Y(io_outs_left_6[15]));
 BUFx2_ASAP7_75t_R output3016 (.A(net3016),
    .Y(io_outs_left_6[16]));
 BUFx2_ASAP7_75t_R output3017 (.A(net3017),
    .Y(io_outs_left_6[17]));
 BUFx2_ASAP7_75t_R output3018 (.A(net3018),
    .Y(io_outs_left_6[18]));
 BUFx2_ASAP7_75t_R output3019 (.A(net3019),
    .Y(io_outs_left_6[19]));
 BUFx2_ASAP7_75t_R output3020 (.A(net3020),
    .Y(io_outs_left_6[1]));
 BUFx2_ASAP7_75t_R output3021 (.A(net3021),
    .Y(io_outs_left_6[20]));
 BUFx2_ASAP7_75t_R output3022 (.A(net3022),
    .Y(io_outs_left_6[21]));
 BUFx2_ASAP7_75t_R output3023 (.A(net3023),
    .Y(io_outs_left_6[22]));
 BUFx2_ASAP7_75t_R output3024 (.A(net3024),
    .Y(io_outs_left_6[23]));
 BUFx2_ASAP7_75t_R output3025 (.A(net3025),
    .Y(io_outs_left_6[24]));
 BUFx2_ASAP7_75t_R output3026 (.A(net3026),
    .Y(io_outs_left_6[25]));
 BUFx2_ASAP7_75t_R output3027 (.A(net3027),
    .Y(io_outs_left_6[26]));
 BUFx2_ASAP7_75t_R output3028 (.A(net3028),
    .Y(io_outs_left_6[27]));
 BUFx2_ASAP7_75t_R output3029 (.A(net3029),
    .Y(io_outs_left_6[28]));
 BUFx2_ASAP7_75t_R output3030 (.A(net3030),
    .Y(io_outs_left_6[29]));
 BUFx2_ASAP7_75t_R output3031 (.A(net3031),
    .Y(io_outs_left_6[2]));
 BUFx2_ASAP7_75t_R output3032 (.A(net3032),
    .Y(io_outs_left_6[30]));
 BUFx2_ASAP7_75t_R output3033 (.A(net3033),
    .Y(io_outs_left_6[31]));
 BUFx2_ASAP7_75t_R output3034 (.A(net3034),
    .Y(io_outs_left_6[32]));
 BUFx2_ASAP7_75t_R output3035 (.A(net3035),
    .Y(io_outs_left_6[33]));
 BUFx2_ASAP7_75t_R output3036 (.A(net3036),
    .Y(io_outs_left_6[34]));
 BUFx2_ASAP7_75t_R output3037 (.A(net3037),
    .Y(io_outs_left_6[35]));
 BUFx2_ASAP7_75t_R output3038 (.A(net3038),
    .Y(io_outs_left_6[36]));
 BUFx2_ASAP7_75t_R output3039 (.A(net3039),
    .Y(io_outs_left_6[37]));
 BUFx2_ASAP7_75t_R output3040 (.A(net3040),
    .Y(io_outs_left_6[38]));
 BUFx2_ASAP7_75t_R output3041 (.A(net3041),
    .Y(io_outs_left_6[39]));
 BUFx2_ASAP7_75t_R output3042 (.A(net3042),
    .Y(io_outs_left_6[3]));
 BUFx2_ASAP7_75t_R output3043 (.A(net3043),
    .Y(io_outs_left_6[40]));
 BUFx2_ASAP7_75t_R output3044 (.A(net3044),
    .Y(io_outs_left_6[41]));
 BUFx2_ASAP7_75t_R output3045 (.A(net3045),
    .Y(io_outs_left_6[42]));
 BUFx2_ASAP7_75t_R output3046 (.A(net3046),
    .Y(io_outs_left_6[43]));
 BUFx2_ASAP7_75t_R output3047 (.A(net3047),
    .Y(io_outs_left_6[44]));
 BUFx2_ASAP7_75t_R output3048 (.A(net3048),
    .Y(io_outs_left_6[45]));
 BUFx2_ASAP7_75t_R output3049 (.A(net3049),
    .Y(io_outs_left_6[46]));
 BUFx2_ASAP7_75t_R output3050 (.A(net3050),
    .Y(io_outs_left_6[47]));
 BUFx2_ASAP7_75t_R output3051 (.A(net3051),
    .Y(io_outs_left_6[48]));
 BUFx2_ASAP7_75t_R output3052 (.A(net3052),
    .Y(io_outs_left_6[49]));
 BUFx2_ASAP7_75t_R output3053 (.A(net3053),
    .Y(io_outs_left_6[4]));
 BUFx2_ASAP7_75t_R output3054 (.A(net3054),
    .Y(io_outs_left_6[50]));
 BUFx2_ASAP7_75t_R output3055 (.A(net3055),
    .Y(io_outs_left_6[51]));
 BUFx2_ASAP7_75t_R output3056 (.A(net3056),
    .Y(io_outs_left_6[52]));
 BUFx2_ASAP7_75t_R output3057 (.A(net3057),
    .Y(io_outs_left_6[53]));
 BUFx2_ASAP7_75t_R output3058 (.A(net3058),
    .Y(io_outs_left_6[54]));
 BUFx2_ASAP7_75t_R output3059 (.A(net3059),
    .Y(io_outs_left_6[55]));
 BUFx2_ASAP7_75t_R output3060 (.A(net3060),
    .Y(io_outs_left_6[56]));
 BUFx2_ASAP7_75t_R output3061 (.A(net3061),
    .Y(io_outs_left_6[57]));
 BUFx2_ASAP7_75t_R output3062 (.A(net3062),
    .Y(io_outs_left_6[58]));
 BUFx2_ASAP7_75t_R output3063 (.A(net3063),
    .Y(io_outs_left_6[59]));
 BUFx2_ASAP7_75t_R output3064 (.A(net3064),
    .Y(io_outs_left_6[5]));
 BUFx2_ASAP7_75t_R output3065 (.A(net3065),
    .Y(io_outs_left_6[60]));
 BUFx2_ASAP7_75t_R output3066 (.A(net3066),
    .Y(io_outs_left_6[61]));
 BUFx2_ASAP7_75t_R output3067 (.A(net3067),
    .Y(io_outs_left_6[62]));
 BUFx2_ASAP7_75t_R output3068 (.A(net3068),
    .Y(io_outs_left_6[63]));
 BUFx2_ASAP7_75t_R output3069 (.A(net3069),
    .Y(io_outs_left_6[6]));
 BUFx2_ASAP7_75t_R output3070 (.A(net3070),
    .Y(io_outs_left_6[7]));
 BUFx2_ASAP7_75t_R output3071 (.A(net3071),
    .Y(io_outs_left_6[8]));
 BUFx2_ASAP7_75t_R output3072 (.A(net3072),
    .Y(io_outs_left_6[9]));
 BUFx2_ASAP7_75t_R output3073 (.A(net3073),
    .Y(io_outs_left_7[0]));
 BUFx2_ASAP7_75t_R output3074 (.A(net3074),
    .Y(io_outs_left_7[10]));
 BUFx2_ASAP7_75t_R output3075 (.A(net3075),
    .Y(io_outs_left_7[11]));
 BUFx2_ASAP7_75t_R output3076 (.A(net3076),
    .Y(io_outs_left_7[12]));
 BUFx2_ASAP7_75t_R output3077 (.A(net3077),
    .Y(io_outs_left_7[13]));
 BUFx2_ASAP7_75t_R output3078 (.A(net3078),
    .Y(io_outs_left_7[14]));
 BUFx2_ASAP7_75t_R output3079 (.A(net3079),
    .Y(io_outs_left_7[15]));
 BUFx2_ASAP7_75t_R output3080 (.A(net3080),
    .Y(io_outs_left_7[16]));
 BUFx2_ASAP7_75t_R output3081 (.A(net3081),
    .Y(io_outs_left_7[17]));
 BUFx2_ASAP7_75t_R output3082 (.A(net3082),
    .Y(io_outs_left_7[18]));
 BUFx2_ASAP7_75t_R output3083 (.A(net3083),
    .Y(io_outs_left_7[19]));
 BUFx2_ASAP7_75t_R output3084 (.A(net3084),
    .Y(io_outs_left_7[1]));
 BUFx2_ASAP7_75t_R output3085 (.A(net3085),
    .Y(io_outs_left_7[20]));
 BUFx2_ASAP7_75t_R output3086 (.A(net3086),
    .Y(io_outs_left_7[21]));
 BUFx2_ASAP7_75t_R output3087 (.A(net3087),
    .Y(io_outs_left_7[22]));
 BUFx2_ASAP7_75t_R output3088 (.A(net3088),
    .Y(io_outs_left_7[23]));
 BUFx2_ASAP7_75t_R output3089 (.A(net3089),
    .Y(io_outs_left_7[24]));
 BUFx2_ASAP7_75t_R output3090 (.A(net3090),
    .Y(io_outs_left_7[25]));
 BUFx2_ASAP7_75t_R output3091 (.A(net3091),
    .Y(io_outs_left_7[26]));
 BUFx2_ASAP7_75t_R output3092 (.A(net3092),
    .Y(io_outs_left_7[27]));
 BUFx2_ASAP7_75t_R output3093 (.A(net3093),
    .Y(io_outs_left_7[28]));
 BUFx2_ASAP7_75t_R output3094 (.A(net3094),
    .Y(io_outs_left_7[29]));
 BUFx2_ASAP7_75t_R output3095 (.A(net3095),
    .Y(io_outs_left_7[2]));
 BUFx2_ASAP7_75t_R output3096 (.A(net3096),
    .Y(io_outs_left_7[30]));
 BUFx2_ASAP7_75t_R output3097 (.A(net3097),
    .Y(io_outs_left_7[31]));
 BUFx2_ASAP7_75t_R output3098 (.A(net3098),
    .Y(io_outs_left_7[32]));
 BUFx2_ASAP7_75t_R output3099 (.A(net3099),
    .Y(io_outs_left_7[33]));
 BUFx2_ASAP7_75t_R output3100 (.A(net3100),
    .Y(io_outs_left_7[34]));
 BUFx2_ASAP7_75t_R output3101 (.A(net3101),
    .Y(io_outs_left_7[35]));
 BUFx2_ASAP7_75t_R output3102 (.A(net3102),
    .Y(io_outs_left_7[36]));
 BUFx2_ASAP7_75t_R output3103 (.A(net3103),
    .Y(io_outs_left_7[37]));
 BUFx2_ASAP7_75t_R output3104 (.A(net3104),
    .Y(io_outs_left_7[38]));
 BUFx2_ASAP7_75t_R output3105 (.A(net3105),
    .Y(io_outs_left_7[39]));
 BUFx2_ASAP7_75t_R output3106 (.A(net3106),
    .Y(io_outs_left_7[3]));
 BUFx2_ASAP7_75t_R output3107 (.A(net3107),
    .Y(io_outs_left_7[40]));
 BUFx2_ASAP7_75t_R output3108 (.A(net3108),
    .Y(io_outs_left_7[41]));
 BUFx2_ASAP7_75t_R output3109 (.A(net3109),
    .Y(io_outs_left_7[42]));
 BUFx2_ASAP7_75t_R output3110 (.A(net3110),
    .Y(io_outs_left_7[43]));
 BUFx2_ASAP7_75t_R output3111 (.A(net3111),
    .Y(io_outs_left_7[44]));
 BUFx2_ASAP7_75t_R output3112 (.A(net3112),
    .Y(io_outs_left_7[45]));
 BUFx2_ASAP7_75t_R output3113 (.A(net3113),
    .Y(io_outs_left_7[46]));
 BUFx2_ASAP7_75t_R output3114 (.A(net3114),
    .Y(io_outs_left_7[47]));
 BUFx2_ASAP7_75t_R output3115 (.A(net3115),
    .Y(io_outs_left_7[48]));
 BUFx2_ASAP7_75t_R output3116 (.A(net3116),
    .Y(io_outs_left_7[49]));
 BUFx2_ASAP7_75t_R output3117 (.A(net3117),
    .Y(io_outs_left_7[4]));
 BUFx2_ASAP7_75t_R output3118 (.A(net3118),
    .Y(io_outs_left_7[50]));
 BUFx2_ASAP7_75t_R output3119 (.A(net3119),
    .Y(io_outs_left_7[51]));
 BUFx2_ASAP7_75t_R output3120 (.A(net3120),
    .Y(io_outs_left_7[52]));
 BUFx2_ASAP7_75t_R output3121 (.A(net3121),
    .Y(io_outs_left_7[53]));
 BUFx2_ASAP7_75t_R output3122 (.A(net3122),
    .Y(io_outs_left_7[54]));
 BUFx2_ASAP7_75t_R output3123 (.A(net3123),
    .Y(io_outs_left_7[55]));
 BUFx2_ASAP7_75t_R output3124 (.A(net3124),
    .Y(io_outs_left_7[56]));
 BUFx2_ASAP7_75t_R output3125 (.A(net3125),
    .Y(io_outs_left_7[57]));
 BUFx2_ASAP7_75t_R output3126 (.A(net3126),
    .Y(io_outs_left_7[58]));
 BUFx2_ASAP7_75t_R output3127 (.A(net3127),
    .Y(io_outs_left_7[59]));
 BUFx2_ASAP7_75t_R output3128 (.A(net3128),
    .Y(io_outs_left_7[5]));
 BUFx2_ASAP7_75t_R output3129 (.A(net3129),
    .Y(io_outs_left_7[60]));
 BUFx2_ASAP7_75t_R output3130 (.A(net3130),
    .Y(io_outs_left_7[61]));
 BUFx2_ASAP7_75t_R output3131 (.A(net3131),
    .Y(io_outs_left_7[62]));
 BUFx2_ASAP7_75t_R output3132 (.A(net3132),
    .Y(io_outs_left_7[63]));
 BUFx2_ASAP7_75t_R output3133 (.A(net3133),
    .Y(io_outs_left_7[6]));
 BUFx2_ASAP7_75t_R output3134 (.A(net3134),
    .Y(io_outs_left_7[7]));
 BUFx2_ASAP7_75t_R output3135 (.A(net3135),
    .Y(io_outs_left_7[8]));
 BUFx2_ASAP7_75t_R output3136 (.A(net3136),
    .Y(io_outs_left_7[9]));
 BUFx2_ASAP7_75t_R output3137 (.A(net3137),
    .Y(io_outs_right_0[0]));
 BUFx2_ASAP7_75t_R output3138 (.A(net3138),
    .Y(io_outs_right_0[10]));
 BUFx2_ASAP7_75t_R output3139 (.A(net3139),
    .Y(io_outs_right_0[11]));
 BUFx2_ASAP7_75t_R output3140 (.A(net3140),
    .Y(io_outs_right_0[12]));
 BUFx2_ASAP7_75t_R output3141 (.A(net3141),
    .Y(io_outs_right_0[13]));
 BUFx2_ASAP7_75t_R output3142 (.A(net3142),
    .Y(io_outs_right_0[14]));
 BUFx2_ASAP7_75t_R output3143 (.A(net3143),
    .Y(io_outs_right_0[15]));
 BUFx2_ASAP7_75t_R output3144 (.A(net3144),
    .Y(io_outs_right_0[16]));
 BUFx2_ASAP7_75t_R output3145 (.A(net3145),
    .Y(io_outs_right_0[17]));
 BUFx2_ASAP7_75t_R output3146 (.A(net3146),
    .Y(io_outs_right_0[18]));
 BUFx2_ASAP7_75t_R output3147 (.A(net3147),
    .Y(io_outs_right_0[19]));
 BUFx2_ASAP7_75t_R output3148 (.A(net3148),
    .Y(io_outs_right_0[1]));
 BUFx2_ASAP7_75t_R output3149 (.A(net3149),
    .Y(io_outs_right_0[20]));
 BUFx2_ASAP7_75t_R output3150 (.A(net3150),
    .Y(io_outs_right_0[21]));
 BUFx2_ASAP7_75t_R output3151 (.A(net3151),
    .Y(io_outs_right_0[22]));
 BUFx2_ASAP7_75t_R output3152 (.A(net3152),
    .Y(io_outs_right_0[23]));
 BUFx2_ASAP7_75t_R output3153 (.A(net3153),
    .Y(io_outs_right_0[24]));
 BUFx2_ASAP7_75t_R output3154 (.A(net3154),
    .Y(io_outs_right_0[25]));
 BUFx2_ASAP7_75t_R output3155 (.A(net3155),
    .Y(io_outs_right_0[26]));
 BUFx2_ASAP7_75t_R output3156 (.A(net3156),
    .Y(io_outs_right_0[27]));
 BUFx2_ASAP7_75t_R output3157 (.A(net3157),
    .Y(io_outs_right_0[28]));
 BUFx2_ASAP7_75t_R output3158 (.A(net3158),
    .Y(io_outs_right_0[29]));
 BUFx2_ASAP7_75t_R output3159 (.A(net3159),
    .Y(io_outs_right_0[2]));
 BUFx2_ASAP7_75t_R output3160 (.A(net3160),
    .Y(io_outs_right_0[30]));
 BUFx2_ASAP7_75t_R output3161 (.A(net3161),
    .Y(io_outs_right_0[31]));
 BUFx2_ASAP7_75t_R output3162 (.A(net3162),
    .Y(io_outs_right_0[32]));
 BUFx2_ASAP7_75t_R output3163 (.A(net3163),
    .Y(io_outs_right_0[33]));
 BUFx2_ASAP7_75t_R output3164 (.A(net3164),
    .Y(io_outs_right_0[34]));
 BUFx2_ASAP7_75t_R output3165 (.A(net3165),
    .Y(io_outs_right_0[35]));
 BUFx2_ASAP7_75t_R output3166 (.A(net3166),
    .Y(io_outs_right_0[36]));
 BUFx2_ASAP7_75t_R output3167 (.A(net3167),
    .Y(io_outs_right_0[37]));
 BUFx2_ASAP7_75t_R output3168 (.A(net3168),
    .Y(io_outs_right_0[38]));
 BUFx2_ASAP7_75t_R output3169 (.A(net3169),
    .Y(io_outs_right_0[39]));
 BUFx2_ASAP7_75t_R output3170 (.A(net3170),
    .Y(io_outs_right_0[3]));
 BUFx2_ASAP7_75t_R output3171 (.A(net3171),
    .Y(io_outs_right_0[40]));
 BUFx2_ASAP7_75t_R output3172 (.A(net3172),
    .Y(io_outs_right_0[41]));
 BUFx2_ASAP7_75t_R output3173 (.A(net3173),
    .Y(io_outs_right_0[42]));
 BUFx2_ASAP7_75t_R output3174 (.A(net3174),
    .Y(io_outs_right_0[43]));
 BUFx2_ASAP7_75t_R output3175 (.A(net3175),
    .Y(io_outs_right_0[44]));
 BUFx2_ASAP7_75t_R output3176 (.A(net3176),
    .Y(io_outs_right_0[45]));
 BUFx2_ASAP7_75t_R output3177 (.A(net3177),
    .Y(io_outs_right_0[46]));
 BUFx2_ASAP7_75t_R output3178 (.A(net3178),
    .Y(io_outs_right_0[47]));
 BUFx2_ASAP7_75t_R output3179 (.A(net3179),
    .Y(io_outs_right_0[48]));
 BUFx2_ASAP7_75t_R output3180 (.A(net3180),
    .Y(io_outs_right_0[49]));
 BUFx2_ASAP7_75t_R output3181 (.A(net3181),
    .Y(io_outs_right_0[4]));
 BUFx2_ASAP7_75t_R output3182 (.A(net3182),
    .Y(io_outs_right_0[50]));
 BUFx2_ASAP7_75t_R output3183 (.A(net3183),
    .Y(io_outs_right_0[51]));
 BUFx2_ASAP7_75t_R output3184 (.A(net3184),
    .Y(io_outs_right_0[52]));
 BUFx2_ASAP7_75t_R output3185 (.A(net3185),
    .Y(io_outs_right_0[53]));
 BUFx2_ASAP7_75t_R output3186 (.A(net3186),
    .Y(io_outs_right_0[54]));
 BUFx2_ASAP7_75t_R output3187 (.A(net3187),
    .Y(io_outs_right_0[55]));
 BUFx2_ASAP7_75t_R output3188 (.A(net3188),
    .Y(io_outs_right_0[56]));
 BUFx2_ASAP7_75t_R output3189 (.A(net3189),
    .Y(io_outs_right_0[57]));
 BUFx2_ASAP7_75t_R output3190 (.A(net3190),
    .Y(io_outs_right_0[58]));
 BUFx2_ASAP7_75t_R output3191 (.A(net3191),
    .Y(io_outs_right_0[59]));
 BUFx2_ASAP7_75t_R output3192 (.A(net3192),
    .Y(io_outs_right_0[5]));
 BUFx2_ASAP7_75t_R output3193 (.A(net3193),
    .Y(io_outs_right_0[60]));
 BUFx2_ASAP7_75t_R output3194 (.A(net3194),
    .Y(io_outs_right_0[61]));
 BUFx2_ASAP7_75t_R output3195 (.A(net3195),
    .Y(io_outs_right_0[62]));
 BUFx2_ASAP7_75t_R output3196 (.A(net3196),
    .Y(io_outs_right_0[63]));
 BUFx2_ASAP7_75t_R output3197 (.A(net3197),
    .Y(io_outs_right_0[6]));
 BUFx2_ASAP7_75t_R output3198 (.A(net3198),
    .Y(io_outs_right_0[7]));
 BUFx2_ASAP7_75t_R output3199 (.A(net3199),
    .Y(io_outs_right_0[8]));
 BUFx2_ASAP7_75t_R output3200 (.A(net3200),
    .Y(io_outs_right_0[9]));
 BUFx2_ASAP7_75t_R output3201 (.A(net3201),
    .Y(io_outs_right_1[0]));
 BUFx2_ASAP7_75t_R output3202 (.A(net3202),
    .Y(io_outs_right_1[10]));
 BUFx2_ASAP7_75t_R output3203 (.A(net3203),
    .Y(io_outs_right_1[11]));
 BUFx2_ASAP7_75t_R output3204 (.A(net3204),
    .Y(io_outs_right_1[12]));
 BUFx2_ASAP7_75t_R output3205 (.A(net3205),
    .Y(io_outs_right_1[13]));
 BUFx2_ASAP7_75t_R output3206 (.A(net3206),
    .Y(io_outs_right_1[14]));
 BUFx2_ASAP7_75t_R output3207 (.A(net3207),
    .Y(io_outs_right_1[15]));
 BUFx2_ASAP7_75t_R output3208 (.A(net3208),
    .Y(io_outs_right_1[16]));
 BUFx2_ASAP7_75t_R output3209 (.A(net3209),
    .Y(io_outs_right_1[17]));
 BUFx2_ASAP7_75t_R output3210 (.A(net3210),
    .Y(io_outs_right_1[18]));
 BUFx2_ASAP7_75t_R output3211 (.A(net3211),
    .Y(io_outs_right_1[19]));
 BUFx2_ASAP7_75t_R output3212 (.A(net3212),
    .Y(io_outs_right_1[1]));
 BUFx2_ASAP7_75t_R output3213 (.A(net3213),
    .Y(io_outs_right_1[20]));
 BUFx2_ASAP7_75t_R output3214 (.A(net3214),
    .Y(io_outs_right_1[21]));
 BUFx2_ASAP7_75t_R output3215 (.A(net3215),
    .Y(io_outs_right_1[22]));
 BUFx2_ASAP7_75t_R output3216 (.A(net3216),
    .Y(io_outs_right_1[23]));
 BUFx2_ASAP7_75t_R output3217 (.A(net3217),
    .Y(io_outs_right_1[24]));
 BUFx2_ASAP7_75t_R output3218 (.A(net3218),
    .Y(io_outs_right_1[25]));
 BUFx2_ASAP7_75t_R output3219 (.A(net3219),
    .Y(io_outs_right_1[26]));
 BUFx2_ASAP7_75t_R output3220 (.A(net3220),
    .Y(io_outs_right_1[27]));
 BUFx2_ASAP7_75t_R output3221 (.A(net3221),
    .Y(io_outs_right_1[28]));
 BUFx2_ASAP7_75t_R output3222 (.A(net3222),
    .Y(io_outs_right_1[29]));
 BUFx2_ASAP7_75t_R output3223 (.A(net3223),
    .Y(io_outs_right_1[2]));
 BUFx2_ASAP7_75t_R output3224 (.A(net3224),
    .Y(io_outs_right_1[30]));
 BUFx2_ASAP7_75t_R output3225 (.A(net3225),
    .Y(io_outs_right_1[31]));
 BUFx2_ASAP7_75t_R output3226 (.A(net3226),
    .Y(io_outs_right_1[32]));
 BUFx2_ASAP7_75t_R output3227 (.A(net3227),
    .Y(io_outs_right_1[33]));
 BUFx2_ASAP7_75t_R output3228 (.A(net3228),
    .Y(io_outs_right_1[34]));
 BUFx2_ASAP7_75t_R output3229 (.A(net3229),
    .Y(io_outs_right_1[35]));
 BUFx2_ASAP7_75t_R output3230 (.A(net3230),
    .Y(io_outs_right_1[36]));
 BUFx2_ASAP7_75t_R output3231 (.A(net3231),
    .Y(io_outs_right_1[37]));
 BUFx2_ASAP7_75t_R output3232 (.A(net3232),
    .Y(io_outs_right_1[38]));
 BUFx2_ASAP7_75t_R output3233 (.A(net3233),
    .Y(io_outs_right_1[39]));
 BUFx2_ASAP7_75t_R output3234 (.A(net3234),
    .Y(io_outs_right_1[3]));
 BUFx2_ASAP7_75t_R output3235 (.A(net3235),
    .Y(io_outs_right_1[40]));
 BUFx2_ASAP7_75t_R output3236 (.A(net3236),
    .Y(io_outs_right_1[41]));
 BUFx2_ASAP7_75t_R output3237 (.A(net3237),
    .Y(io_outs_right_1[42]));
 BUFx2_ASAP7_75t_R output3238 (.A(net3238),
    .Y(io_outs_right_1[43]));
 BUFx2_ASAP7_75t_R output3239 (.A(net3239),
    .Y(io_outs_right_1[44]));
 BUFx2_ASAP7_75t_R output3240 (.A(net3240),
    .Y(io_outs_right_1[45]));
 BUFx2_ASAP7_75t_R output3241 (.A(net3241),
    .Y(io_outs_right_1[46]));
 BUFx2_ASAP7_75t_R output3242 (.A(net3242),
    .Y(io_outs_right_1[47]));
 BUFx2_ASAP7_75t_R output3243 (.A(net3243),
    .Y(io_outs_right_1[48]));
 BUFx2_ASAP7_75t_R output3244 (.A(net3244),
    .Y(io_outs_right_1[49]));
 BUFx2_ASAP7_75t_R output3245 (.A(net3245),
    .Y(io_outs_right_1[4]));
 BUFx2_ASAP7_75t_R output3246 (.A(net3246),
    .Y(io_outs_right_1[50]));
 BUFx2_ASAP7_75t_R output3247 (.A(net3247),
    .Y(io_outs_right_1[51]));
 BUFx2_ASAP7_75t_R output3248 (.A(net3248),
    .Y(io_outs_right_1[52]));
 BUFx2_ASAP7_75t_R output3249 (.A(net3249),
    .Y(io_outs_right_1[53]));
 BUFx2_ASAP7_75t_R output3250 (.A(net3250),
    .Y(io_outs_right_1[54]));
 BUFx2_ASAP7_75t_R output3251 (.A(net3251),
    .Y(io_outs_right_1[55]));
 BUFx2_ASAP7_75t_R output3252 (.A(net3252),
    .Y(io_outs_right_1[56]));
 BUFx2_ASAP7_75t_R output3253 (.A(net3253),
    .Y(io_outs_right_1[57]));
 BUFx2_ASAP7_75t_R output3254 (.A(net3254),
    .Y(io_outs_right_1[58]));
 BUFx2_ASAP7_75t_R output3255 (.A(net3255),
    .Y(io_outs_right_1[59]));
 BUFx2_ASAP7_75t_R output3256 (.A(net3256),
    .Y(io_outs_right_1[5]));
 BUFx2_ASAP7_75t_R output3257 (.A(net3257),
    .Y(io_outs_right_1[60]));
 BUFx2_ASAP7_75t_R output3258 (.A(net3258),
    .Y(io_outs_right_1[61]));
 BUFx2_ASAP7_75t_R output3259 (.A(net3259),
    .Y(io_outs_right_1[62]));
 BUFx2_ASAP7_75t_R output3260 (.A(net3260),
    .Y(io_outs_right_1[63]));
 BUFx2_ASAP7_75t_R output3261 (.A(net3261),
    .Y(io_outs_right_1[6]));
 BUFx2_ASAP7_75t_R output3262 (.A(net3262),
    .Y(io_outs_right_1[7]));
 BUFx2_ASAP7_75t_R output3263 (.A(net3263),
    .Y(io_outs_right_1[8]));
 BUFx2_ASAP7_75t_R output3264 (.A(net3264),
    .Y(io_outs_right_1[9]));
 BUFx2_ASAP7_75t_R output3265 (.A(net3265),
    .Y(io_outs_right_2[0]));
 BUFx2_ASAP7_75t_R output3266 (.A(net3266),
    .Y(io_outs_right_2[10]));
 BUFx2_ASAP7_75t_R output3267 (.A(net3267),
    .Y(io_outs_right_2[11]));
 BUFx2_ASAP7_75t_R output3268 (.A(net3268),
    .Y(io_outs_right_2[12]));
 BUFx2_ASAP7_75t_R output3269 (.A(net3269),
    .Y(io_outs_right_2[13]));
 BUFx2_ASAP7_75t_R output3270 (.A(net3270),
    .Y(io_outs_right_2[14]));
 BUFx2_ASAP7_75t_R output3271 (.A(net3271),
    .Y(io_outs_right_2[15]));
 BUFx2_ASAP7_75t_R output3272 (.A(net3272),
    .Y(io_outs_right_2[16]));
 BUFx2_ASAP7_75t_R output3273 (.A(net3273),
    .Y(io_outs_right_2[17]));
 BUFx2_ASAP7_75t_R output3274 (.A(net3274),
    .Y(io_outs_right_2[18]));
 BUFx2_ASAP7_75t_R output3275 (.A(net3275),
    .Y(io_outs_right_2[19]));
 BUFx2_ASAP7_75t_R output3276 (.A(net3276),
    .Y(io_outs_right_2[1]));
 BUFx2_ASAP7_75t_R output3277 (.A(net3277),
    .Y(io_outs_right_2[20]));
 BUFx2_ASAP7_75t_R output3278 (.A(net3278),
    .Y(io_outs_right_2[21]));
 BUFx2_ASAP7_75t_R output3279 (.A(net3279),
    .Y(io_outs_right_2[22]));
 BUFx2_ASAP7_75t_R output3280 (.A(net3280),
    .Y(io_outs_right_2[23]));
 BUFx2_ASAP7_75t_R output3281 (.A(net3281),
    .Y(io_outs_right_2[24]));
 BUFx2_ASAP7_75t_R output3282 (.A(net3282),
    .Y(io_outs_right_2[25]));
 BUFx2_ASAP7_75t_R output3283 (.A(net3283),
    .Y(io_outs_right_2[26]));
 BUFx2_ASAP7_75t_R output3284 (.A(net3284),
    .Y(io_outs_right_2[27]));
 BUFx2_ASAP7_75t_R output3285 (.A(net3285),
    .Y(io_outs_right_2[28]));
 BUFx2_ASAP7_75t_R output3286 (.A(net3286),
    .Y(io_outs_right_2[29]));
 BUFx2_ASAP7_75t_R output3287 (.A(net3287),
    .Y(io_outs_right_2[2]));
 BUFx2_ASAP7_75t_R output3288 (.A(net3288),
    .Y(io_outs_right_2[30]));
 BUFx2_ASAP7_75t_R output3289 (.A(net3289),
    .Y(io_outs_right_2[31]));
 BUFx2_ASAP7_75t_R output3290 (.A(net3290),
    .Y(io_outs_right_2[32]));
 BUFx2_ASAP7_75t_R output3291 (.A(net3291),
    .Y(io_outs_right_2[33]));
 BUFx2_ASAP7_75t_R output3292 (.A(net3292),
    .Y(io_outs_right_2[34]));
 BUFx2_ASAP7_75t_R output3293 (.A(net3293),
    .Y(io_outs_right_2[35]));
 BUFx2_ASAP7_75t_R output3294 (.A(net3294),
    .Y(io_outs_right_2[36]));
 BUFx2_ASAP7_75t_R output3295 (.A(net3295),
    .Y(io_outs_right_2[37]));
 BUFx2_ASAP7_75t_R output3296 (.A(net3296),
    .Y(io_outs_right_2[38]));
 BUFx2_ASAP7_75t_R output3297 (.A(net3297),
    .Y(io_outs_right_2[39]));
 BUFx2_ASAP7_75t_R output3298 (.A(net3298),
    .Y(io_outs_right_2[3]));
 BUFx2_ASAP7_75t_R output3299 (.A(net3299),
    .Y(io_outs_right_2[40]));
 BUFx2_ASAP7_75t_R output3300 (.A(net3300),
    .Y(io_outs_right_2[41]));
 BUFx2_ASAP7_75t_R output3301 (.A(net3301),
    .Y(io_outs_right_2[42]));
 BUFx2_ASAP7_75t_R output3302 (.A(net3302),
    .Y(io_outs_right_2[43]));
 BUFx2_ASAP7_75t_R output3303 (.A(net3303),
    .Y(io_outs_right_2[44]));
 BUFx2_ASAP7_75t_R output3304 (.A(net3304),
    .Y(io_outs_right_2[45]));
 BUFx2_ASAP7_75t_R output3305 (.A(net3305),
    .Y(io_outs_right_2[46]));
 BUFx2_ASAP7_75t_R output3306 (.A(net3306),
    .Y(io_outs_right_2[47]));
 BUFx2_ASAP7_75t_R output3307 (.A(net3307),
    .Y(io_outs_right_2[48]));
 BUFx2_ASAP7_75t_R output3308 (.A(net3308),
    .Y(io_outs_right_2[49]));
 BUFx2_ASAP7_75t_R output3309 (.A(net3309),
    .Y(io_outs_right_2[4]));
 BUFx2_ASAP7_75t_R output3310 (.A(net3310),
    .Y(io_outs_right_2[50]));
 BUFx2_ASAP7_75t_R output3311 (.A(net3311),
    .Y(io_outs_right_2[51]));
 BUFx2_ASAP7_75t_R output3312 (.A(net3312),
    .Y(io_outs_right_2[52]));
 BUFx2_ASAP7_75t_R output3313 (.A(net3313),
    .Y(io_outs_right_2[53]));
 BUFx2_ASAP7_75t_R output3314 (.A(net3314),
    .Y(io_outs_right_2[54]));
 BUFx2_ASAP7_75t_R output3315 (.A(net3315),
    .Y(io_outs_right_2[55]));
 BUFx2_ASAP7_75t_R output3316 (.A(net3316),
    .Y(io_outs_right_2[56]));
 BUFx2_ASAP7_75t_R output3317 (.A(net3317),
    .Y(io_outs_right_2[57]));
 BUFx2_ASAP7_75t_R output3318 (.A(net3318),
    .Y(io_outs_right_2[58]));
 BUFx2_ASAP7_75t_R output3319 (.A(net3319),
    .Y(io_outs_right_2[59]));
 BUFx2_ASAP7_75t_R output3320 (.A(net3320),
    .Y(io_outs_right_2[5]));
 BUFx2_ASAP7_75t_R output3321 (.A(net3321),
    .Y(io_outs_right_2[60]));
 BUFx2_ASAP7_75t_R output3322 (.A(net3322),
    .Y(io_outs_right_2[61]));
 BUFx2_ASAP7_75t_R output3323 (.A(net3323),
    .Y(io_outs_right_2[62]));
 BUFx2_ASAP7_75t_R output3324 (.A(net3324),
    .Y(io_outs_right_2[63]));
 BUFx2_ASAP7_75t_R output3325 (.A(net3325),
    .Y(io_outs_right_2[6]));
 BUFx2_ASAP7_75t_R output3326 (.A(net3326),
    .Y(io_outs_right_2[7]));
 BUFx2_ASAP7_75t_R output3327 (.A(net3327),
    .Y(io_outs_right_2[8]));
 BUFx2_ASAP7_75t_R output3328 (.A(net3328),
    .Y(io_outs_right_2[9]));
 BUFx2_ASAP7_75t_R output3329 (.A(net3329),
    .Y(io_outs_right_3[0]));
 BUFx2_ASAP7_75t_R output3330 (.A(net3330),
    .Y(io_outs_right_3[10]));
 BUFx2_ASAP7_75t_R output3331 (.A(net3331),
    .Y(io_outs_right_3[11]));
 BUFx2_ASAP7_75t_R output3332 (.A(net3332),
    .Y(io_outs_right_3[12]));
 BUFx2_ASAP7_75t_R output3333 (.A(net3333),
    .Y(io_outs_right_3[13]));
 BUFx2_ASAP7_75t_R output3334 (.A(net3334),
    .Y(io_outs_right_3[14]));
 BUFx2_ASAP7_75t_R output3335 (.A(net3335),
    .Y(io_outs_right_3[15]));
 BUFx2_ASAP7_75t_R output3336 (.A(net3336),
    .Y(io_outs_right_3[16]));
 BUFx2_ASAP7_75t_R output3337 (.A(net3337),
    .Y(io_outs_right_3[17]));
 BUFx2_ASAP7_75t_R output3338 (.A(net3338),
    .Y(io_outs_right_3[18]));
 BUFx2_ASAP7_75t_R output3339 (.A(net3339),
    .Y(io_outs_right_3[19]));
 BUFx2_ASAP7_75t_R output3340 (.A(net3340),
    .Y(io_outs_right_3[1]));
 BUFx2_ASAP7_75t_R output3341 (.A(net3341),
    .Y(io_outs_right_3[20]));
 BUFx2_ASAP7_75t_R output3342 (.A(net3342),
    .Y(io_outs_right_3[21]));
 BUFx2_ASAP7_75t_R output3343 (.A(net3343),
    .Y(io_outs_right_3[22]));
 BUFx2_ASAP7_75t_R output3344 (.A(net3344),
    .Y(io_outs_right_3[23]));
 BUFx2_ASAP7_75t_R output3345 (.A(net3345),
    .Y(io_outs_right_3[24]));
 BUFx2_ASAP7_75t_R output3346 (.A(net3346),
    .Y(io_outs_right_3[25]));
 BUFx2_ASAP7_75t_R output3347 (.A(net3347),
    .Y(io_outs_right_3[26]));
 BUFx2_ASAP7_75t_R output3348 (.A(net3348),
    .Y(io_outs_right_3[27]));
 BUFx2_ASAP7_75t_R output3349 (.A(net3349),
    .Y(io_outs_right_3[28]));
 BUFx2_ASAP7_75t_R output3350 (.A(net3350),
    .Y(io_outs_right_3[29]));
 BUFx2_ASAP7_75t_R output3351 (.A(net3351),
    .Y(io_outs_right_3[2]));
 BUFx2_ASAP7_75t_R output3352 (.A(net3352),
    .Y(io_outs_right_3[30]));
 BUFx2_ASAP7_75t_R output3353 (.A(net3353),
    .Y(io_outs_right_3[31]));
 BUFx2_ASAP7_75t_R output3354 (.A(net3354),
    .Y(io_outs_right_3[32]));
 BUFx2_ASAP7_75t_R output3355 (.A(net3355),
    .Y(io_outs_right_3[33]));
 BUFx2_ASAP7_75t_R output3356 (.A(net3356),
    .Y(io_outs_right_3[34]));
 BUFx2_ASAP7_75t_R output3357 (.A(net3357),
    .Y(io_outs_right_3[35]));
 BUFx2_ASAP7_75t_R output3358 (.A(net3358),
    .Y(io_outs_right_3[36]));
 BUFx2_ASAP7_75t_R output3359 (.A(net3359),
    .Y(io_outs_right_3[37]));
 BUFx2_ASAP7_75t_R output3360 (.A(net3360),
    .Y(io_outs_right_3[38]));
 BUFx2_ASAP7_75t_R output3361 (.A(net3361),
    .Y(io_outs_right_3[39]));
 BUFx2_ASAP7_75t_R output3362 (.A(net3362),
    .Y(io_outs_right_3[3]));
 BUFx2_ASAP7_75t_R output3363 (.A(net3363),
    .Y(io_outs_right_3[40]));
 BUFx2_ASAP7_75t_R output3364 (.A(net3364),
    .Y(io_outs_right_3[41]));
 BUFx2_ASAP7_75t_R output3365 (.A(net3365),
    .Y(io_outs_right_3[42]));
 BUFx2_ASAP7_75t_R output3366 (.A(net3366),
    .Y(io_outs_right_3[43]));
 BUFx2_ASAP7_75t_R output3367 (.A(net3367),
    .Y(io_outs_right_3[44]));
 BUFx2_ASAP7_75t_R output3368 (.A(net3368),
    .Y(io_outs_right_3[45]));
 BUFx2_ASAP7_75t_R output3369 (.A(net3369),
    .Y(io_outs_right_3[46]));
 BUFx2_ASAP7_75t_R output3370 (.A(net3370),
    .Y(io_outs_right_3[47]));
 BUFx2_ASAP7_75t_R output3371 (.A(net3371),
    .Y(io_outs_right_3[48]));
 BUFx2_ASAP7_75t_R output3372 (.A(net3372),
    .Y(io_outs_right_3[49]));
 BUFx2_ASAP7_75t_R output3373 (.A(net3373),
    .Y(io_outs_right_3[4]));
 BUFx2_ASAP7_75t_R output3374 (.A(net3374),
    .Y(io_outs_right_3[50]));
 BUFx2_ASAP7_75t_R output3375 (.A(net3375),
    .Y(io_outs_right_3[51]));
 BUFx2_ASAP7_75t_R output3376 (.A(net3376),
    .Y(io_outs_right_3[52]));
 BUFx2_ASAP7_75t_R output3377 (.A(net3377),
    .Y(io_outs_right_3[53]));
 BUFx2_ASAP7_75t_R output3378 (.A(net3378),
    .Y(io_outs_right_3[54]));
 BUFx2_ASAP7_75t_R output3379 (.A(net3379),
    .Y(io_outs_right_3[55]));
 BUFx2_ASAP7_75t_R output3380 (.A(net3380),
    .Y(io_outs_right_3[56]));
 BUFx2_ASAP7_75t_R output3381 (.A(net3381),
    .Y(io_outs_right_3[57]));
 BUFx2_ASAP7_75t_R output3382 (.A(net3382),
    .Y(io_outs_right_3[58]));
 BUFx2_ASAP7_75t_R output3383 (.A(net3383),
    .Y(io_outs_right_3[59]));
 BUFx2_ASAP7_75t_R output3384 (.A(net3384),
    .Y(io_outs_right_3[5]));
 BUFx2_ASAP7_75t_R output3385 (.A(net3385),
    .Y(io_outs_right_3[60]));
 BUFx2_ASAP7_75t_R output3386 (.A(net3386),
    .Y(io_outs_right_3[61]));
 BUFx2_ASAP7_75t_R output3387 (.A(net3387),
    .Y(io_outs_right_3[62]));
 BUFx2_ASAP7_75t_R output3388 (.A(net3388),
    .Y(io_outs_right_3[63]));
 BUFx2_ASAP7_75t_R output3389 (.A(net3389),
    .Y(io_outs_right_3[6]));
 BUFx2_ASAP7_75t_R output3390 (.A(net3390),
    .Y(io_outs_right_3[7]));
 BUFx2_ASAP7_75t_R output3391 (.A(net3391),
    .Y(io_outs_right_3[8]));
 BUFx2_ASAP7_75t_R output3392 (.A(net3392),
    .Y(io_outs_right_3[9]));
 BUFx2_ASAP7_75t_R output3393 (.A(net3393),
    .Y(io_outs_right_4[0]));
 BUFx2_ASAP7_75t_R output3394 (.A(net3394),
    .Y(io_outs_right_4[10]));
 BUFx2_ASAP7_75t_R output3395 (.A(net3395),
    .Y(io_outs_right_4[11]));
 BUFx2_ASAP7_75t_R output3396 (.A(net3396),
    .Y(io_outs_right_4[12]));
 BUFx2_ASAP7_75t_R output3397 (.A(net3397),
    .Y(io_outs_right_4[13]));
 BUFx2_ASAP7_75t_R output3398 (.A(net3398),
    .Y(io_outs_right_4[14]));
 BUFx2_ASAP7_75t_R output3399 (.A(net3399),
    .Y(io_outs_right_4[15]));
 BUFx2_ASAP7_75t_R output3400 (.A(net3400),
    .Y(io_outs_right_4[16]));
 BUFx2_ASAP7_75t_R output3401 (.A(net3401),
    .Y(io_outs_right_4[17]));
 BUFx2_ASAP7_75t_R output3402 (.A(net3402),
    .Y(io_outs_right_4[18]));
 BUFx2_ASAP7_75t_R output3403 (.A(net3403),
    .Y(io_outs_right_4[19]));
 BUFx2_ASAP7_75t_R output3404 (.A(net3404),
    .Y(io_outs_right_4[1]));
 BUFx2_ASAP7_75t_R output3405 (.A(net3405),
    .Y(io_outs_right_4[20]));
 BUFx2_ASAP7_75t_R output3406 (.A(net3406),
    .Y(io_outs_right_4[21]));
 BUFx2_ASAP7_75t_R output3407 (.A(net3407),
    .Y(io_outs_right_4[22]));
 BUFx2_ASAP7_75t_R output3408 (.A(net3408),
    .Y(io_outs_right_4[23]));
 BUFx2_ASAP7_75t_R output3409 (.A(net3409),
    .Y(io_outs_right_4[24]));
 BUFx2_ASAP7_75t_R output3410 (.A(net3410),
    .Y(io_outs_right_4[25]));
 BUFx2_ASAP7_75t_R output3411 (.A(net3411),
    .Y(io_outs_right_4[26]));
 BUFx2_ASAP7_75t_R output3412 (.A(net3412),
    .Y(io_outs_right_4[27]));
 BUFx2_ASAP7_75t_R output3413 (.A(net3413),
    .Y(io_outs_right_4[28]));
 BUFx2_ASAP7_75t_R output3414 (.A(net3414),
    .Y(io_outs_right_4[29]));
 BUFx2_ASAP7_75t_R output3415 (.A(net3415),
    .Y(io_outs_right_4[2]));
 BUFx2_ASAP7_75t_R output3416 (.A(net3416),
    .Y(io_outs_right_4[30]));
 BUFx2_ASAP7_75t_R output3417 (.A(net3417),
    .Y(io_outs_right_4[31]));
 BUFx2_ASAP7_75t_R output3418 (.A(net3418),
    .Y(io_outs_right_4[32]));
 BUFx2_ASAP7_75t_R output3419 (.A(net3419),
    .Y(io_outs_right_4[33]));
 BUFx2_ASAP7_75t_R output3420 (.A(net3420),
    .Y(io_outs_right_4[34]));
 BUFx2_ASAP7_75t_R output3421 (.A(net3421),
    .Y(io_outs_right_4[35]));
 BUFx2_ASAP7_75t_R output3422 (.A(net3422),
    .Y(io_outs_right_4[36]));
 BUFx2_ASAP7_75t_R output3423 (.A(net3423),
    .Y(io_outs_right_4[37]));
 BUFx2_ASAP7_75t_R output3424 (.A(net3424),
    .Y(io_outs_right_4[38]));
 BUFx2_ASAP7_75t_R output3425 (.A(net3425),
    .Y(io_outs_right_4[39]));
 BUFx2_ASAP7_75t_R output3426 (.A(net3426),
    .Y(io_outs_right_4[3]));
 BUFx2_ASAP7_75t_R output3427 (.A(net3427),
    .Y(io_outs_right_4[40]));
 BUFx2_ASAP7_75t_R output3428 (.A(net3428),
    .Y(io_outs_right_4[41]));
 BUFx2_ASAP7_75t_R output3429 (.A(net3429),
    .Y(io_outs_right_4[42]));
 BUFx2_ASAP7_75t_R output3430 (.A(net3430),
    .Y(io_outs_right_4[43]));
 BUFx2_ASAP7_75t_R output3431 (.A(net3431),
    .Y(io_outs_right_4[44]));
 BUFx2_ASAP7_75t_R output3432 (.A(net3432),
    .Y(io_outs_right_4[45]));
 BUFx2_ASAP7_75t_R output3433 (.A(net3433),
    .Y(io_outs_right_4[46]));
 BUFx2_ASAP7_75t_R output3434 (.A(net3434),
    .Y(io_outs_right_4[47]));
 BUFx2_ASAP7_75t_R output3435 (.A(net3435),
    .Y(io_outs_right_4[48]));
 BUFx2_ASAP7_75t_R output3436 (.A(net3436),
    .Y(io_outs_right_4[49]));
 BUFx2_ASAP7_75t_R output3437 (.A(net3437),
    .Y(io_outs_right_4[4]));
 BUFx2_ASAP7_75t_R output3438 (.A(net3438),
    .Y(io_outs_right_4[50]));
 BUFx2_ASAP7_75t_R output3439 (.A(net3439),
    .Y(io_outs_right_4[51]));
 BUFx2_ASAP7_75t_R output3440 (.A(net3440),
    .Y(io_outs_right_4[52]));
 BUFx2_ASAP7_75t_R output3441 (.A(net3441),
    .Y(io_outs_right_4[53]));
 BUFx2_ASAP7_75t_R output3442 (.A(net3442),
    .Y(io_outs_right_4[54]));
 BUFx2_ASAP7_75t_R output3443 (.A(net3443),
    .Y(io_outs_right_4[55]));
 BUFx2_ASAP7_75t_R output3444 (.A(net3444),
    .Y(io_outs_right_4[56]));
 BUFx2_ASAP7_75t_R output3445 (.A(net3445),
    .Y(io_outs_right_4[57]));
 BUFx2_ASAP7_75t_R output3446 (.A(net3446),
    .Y(io_outs_right_4[58]));
 BUFx2_ASAP7_75t_R output3447 (.A(net3447),
    .Y(io_outs_right_4[59]));
 BUFx2_ASAP7_75t_R output3448 (.A(net3448),
    .Y(io_outs_right_4[5]));
 BUFx2_ASAP7_75t_R output3449 (.A(net3449),
    .Y(io_outs_right_4[60]));
 BUFx2_ASAP7_75t_R output3450 (.A(net3450),
    .Y(io_outs_right_4[61]));
 BUFx2_ASAP7_75t_R output3451 (.A(net3451),
    .Y(io_outs_right_4[62]));
 BUFx2_ASAP7_75t_R output3452 (.A(net3452),
    .Y(io_outs_right_4[63]));
 BUFx2_ASAP7_75t_R output3453 (.A(net3453),
    .Y(io_outs_right_4[6]));
 BUFx2_ASAP7_75t_R output3454 (.A(net3454),
    .Y(io_outs_right_4[7]));
 BUFx2_ASAP7_75t_R output3455 (.A(net3455),
    .Y(io_outs_right_4[8]));
 BUFx2_ASAP7_75t_R output3456 (.A(net3456),
    .Y(io_outs_right_4[9]));
 BUFx2_ASAP7_75t_R output3457 (.A(net3457),
    .Y(io_outs_right_5[0]));
 BUFx2_ASAP7_75t_R output3458 (.A(net3458),
    .Y(io_outs_right_5[10]));
 BUFx2_ASAP7_75t_R output3459 (.A(net3459),
    .Y(io_outs_right_5[11]));
 BUFx2_ASAP7_75t_R output3460 (.A(net3460),
    .Y(io_outs_right_5[12]));
 BUFx2_ASAP7_75t_R output3461 (.A(net3461),
    .Y(io_outs_right_5[13]));
 BUFx2_ASAP7_75t_R output3462 (.A(net3462),
    .Y(io_outs_right_5[14]));
 BUFx2_ASAP7_75t_R output3463 (.A(net3463),
    .Y(io_outs_right_5[15]));
 BUFx2_ASAP7_75t_R output3464 (.A(net3464),
    .Y(io_outs_right_5[16]));
 BUFx2_ASAP7_75t_R output3465 (.A(net3465),
    .Y(io_outs_right_5[17]));
 BUFx2_ASAP7_75t_R output3466 (.A(net3466),
    .Y(io_outs_right_5[18]));
 BUFx2_ASAP7_75t_R output3467 (.A(net3467),
    .Y(io_outs_right_5[19]));
 BUFx2_ASAP7_75t_R output3468 (.A(net3468),
    .Y(io_outs_right_5[1]));
 BUFx2_ASAP7_75t_R output3469 (.A(net3469),
    .Y(io_outs_right_5[20]));
 BUFx2_ASAP7_75t_R output3470 (.A(net3470),
    .Y(io_outs_right_5[21]));
 BUFx2_ASAP7_75t_R output3471 (.A(net3471),
    .Y(io_outs_right_5[22]));
 BUFx2_ASAP7_75t_R output3472 (.A(net3472),
    .Y(io_outs_right_5[23]));
 BUFx2_ASAP7_75t_R output3473 (.A(net3473),
    .Y(io_outs_right_5[24]));
 BUFx2_ASAP7_75t_R output3474 (.A(net3474),
    .Y(io_outs_right_5[25]));
 BUFx2_ASAP7_75t_R output3475 (.A(net3475),
    .Y(io_outs_right_5[26]));
 BUFx2_ASAP7_75t_R output3476 (.A(net3476),
    .Y(io_outs_right_5[27]));
 BUFx2_ASAP7_75t_R output3477 (.A(net3477),
    .Y(io_outs_right_5[28]));
 BUFx2_ASAP7_75t_R output3478 (.A(net3478),
    .Y(io_outs_right_5[29]));
 BUFx2_ASAP7_75t_R output3479 (.A(net3479),
    .Y(io_outs_right_5[2]));
 BUFx2_ASAP7_75t_R output3480 (.A(net3480),
    .Y(io_outs_right_5[30]));
 BUFx2_ASAP7_75t_R output3481 (.A(net3481),
    .Y(io_outs_right_5[31]));
 BUFx2_ASAP7_75t_R output3482 (.A(net3482),
    .Y(io_outs_right_5[32]));
 BUFx2_ASAP7_75t_R output3483 (.A(net3483),
    .Y(io_outs_right_5[33]));
 BUFx2_ASAP7_75t_R output3484 (.A(net3484),
    .Y(io_outs_right_5[34]));
 BUFx2_ASAP7_75t_R output3485 (.A(net3485),
    .Y(io_outs_right_5[35]));
 BUFx2_ASAP7_75t_R output3486 (.A(net3486),
    .Y(io_outs_right_5[36]));
 BUFx2_ASAP7_75t_R output3487 (.A(net3487),
    .Y(io_outs_right_5[37]));
 BUFx2_ASAP7_75t_R output3488 (.A(net3488),
    .Y(io_outs_right_5[38]));
 BUFx2_ASAP7_75t_R output3489 (.A(net3489),
    .Y(io_outs_right_5[39]));
 BUFx2_ASAP7_75t_R output3490 (.A(net3490),
    .Y(io_outs_right_5[3]));
 BUFx2_ASAP7_75t_R output3491 (.A(net3491),
    .Y(io_outs_right_5[40]));
 BUFx2_ASAP7_75t_R output3492 (.A(net3492),
    .Y(io_outs_right_5[41]));
 BUFx2_ASAP7_75t_R output3493 (.A(net3493),
    .Y(io_outs_right_5[42]));
 BUFx2_ASAP7_75t_R output3494 (.A(net3494),
    .Y(io_outs_right_5[43]));
 BUFx2_ASAP7_75t_R output3495 (.A(net3495),
    .Y(io_outs_right_5[44]));
 BUFx2_ASAP7_75t_R output3496 (.A(net3496),
    .Y(io_outs_right_5[45]));
 BUFx2_ASAP7_75t_R output3497 (.A(net3497),
    .Y(io_outs_right_5[46]));
 BUFx2_ASAP7_75t_R output3498 (.A(net3498),
    .Y(io_outs_right_5[47]));
 BUFx2_ASAP7_75t_R output3499 (.A(net3499),
    .Y(io_outs_right_5[48]));
 BUFx2_ASAP7_75t_R output3500 (.A(net3500),
    .Y(io_outs_right_5[49]));
 BUFx2_ASAP7_75t_R output3501 (.A(net3501),
    .Y(io_outs_right_5[4]));
 BUFx2_ASAP7_75t_R output3502 (.A(net3502),
    .Y(io_outs_right_5[50]));
 BUFx2_ASAP7_75t_R output3503 (.A(net3503),
    .Y(io_outs_right_5[51]));
 BUFx2_ASAP7_75t_R output3504 (.A(net3504),
    .Y(io_outs_right_5[52]));
 BUFx2_ASAP7_75t_R output3505 (.A(net3505),
    .Y(io_outs_right_5[53]));
 BUFx2_ASAP7_75t_R output3506 (.A(net3506),
    .Y(io_outs_right_5[54]));
 BUFx2_ASAP7_75t_R output3507 (.A(net3507),
    .Y(io_outs_right_5[55]));
 BUFx2_ASAP7_75t_R output3508 (.A(net3508),
    .Y(io_outs_right_5[56]));
 BUFx2_ASAP7_75t_R output3509 (.A(net3509),
    .Y(io_outs_right_5[57]));
 BUFx2_ASAP7_75t_R output3510 (.A(net3510),
    .Y(io_outs_right_5[58]));
 BUFx2_ASAP7_75t_R output3511 (.A(net3511),
    .Y(io_outs_right_5[59]));
 BUFx2_ASAP7_75t_R output3512 (.A(net3512),
    .Y(io_outs_right_5[5]));
 BUFx2_ASAP7_75t_R output3513 (.A(net3513),
    .Y(io_outs_right_5[60]));
 BUFx2_ASAP7_75t_R output3514 (.A(net3514),
    .Y(io_outs_right_5[61]));
 BUFx2_ASAP7_75t_R output3515 (.A(net3515),
    .Y(io_outs_right_5[62]));
 BUFx2_ASAP7_75t_R output3516 (.A(net3516),
    .Y(io_outs_right_5[63]));
 BUFx2_ASAP7_75t_R output3517 (.A(net3517),
    .Y(io_outs_right_5[6]));
 BUFx2_ASAP7_75t_R output3518 (.A(net3518),
    .Y(io_outs_right_5[7]));
 BUFx2_ASAP7_75t_R output3519 (.A(net3519),
    .Y(io_outs_right_5[8]));
 BUFx2_ASAP7_75t_R output3520 (.A(net3520),
    .Y(io_outs_right_5[9]));
 BUFx2_ASAP7_75t_R output3521 (.A(net3521),
    .Y(io_outs_right_6[0]));
 BUFx2_ASAP7_75t_R output3522 (.A(net3522),
    .Y(io_outs_right_6[10]));
 BUFx2_ASAP7_75t_R output3523 (.A(net3523),
    .Y(io_outs_right_6[11]));
 BUFx2_ASAP7_75t_R output3524 (.A(net3524),
    .Y(io_outs_right_6[12]));
 BUFx2_ASAP7_75t_R output3525 (.A(net3525),
    .Y(io_outs_right_6[13]));
 BUFx2_ASAP7_75t_R output3526 (.A(net3526),
    .Y(io_outs_right_6[14]));
 BUFx2_ASAP7_75t_R output3527 (.A(net3527),
    .Y(io_outs_right_6[15]));
 BUFx2_ASAP7_75t_R output3528 (.A(net3528),
    .Y(io_outs_right_6[16]));
 BUFx2_ASAP7_75t_R output3529 (.A(net3529),
    .Y(io_outs_right_6[17]));
 BUFx2_ASAP7_75t_R output3530 (.A(net3530),
    .Y(io_outs_right_6[18]));
 BUFx2_ASAP7_75t_R output3531 (.A(net3531),
    .Y(io_outs_right_6[19]));
 BUFx2_ASAP7_75t_R output3532 (.A(net3532),
    .Y(io_outs_right_6[1]));
 BUFx2_ASAP7_75t_R output3533 (.A(net3533),
    .Y(io_outs_right_6[20]));
 BUFx2_ASAP7_75t_R output3534 (.A(net3534),
    .Y(io_outs_right_6[21]));
 BUFx2_ASAP7_75t_R output3535 (.A(net3535),
    .Y(io_outs_right_6[22]));
 BUFx2_ASAP7_75t_R output3536 (.A(net3536),
    .Y(io_outs_right_6[23]));
 BUFx2_ASAP7_75t_R output3537 (.A(net3537),
    .Y(io_outs_right_6[24]));
 BUFx2_ASAP7_75t_R output3538 (.A(net3538),
    .Y(io_outs_right_6[25]));
 BUFx2_ASAP7_75t_R output3539 (.A(net3539),
    .Y(io_outs_right_6[26]));
 BUFx2_ASAP7_75t_R output3540 (.A(net3540),
    .Y(io_outs_right_6[27]));
 BUFx2_ASAP7_75t_R output3541 (.A(net3541),
    .Y(io_outs_right_6[28]));
 BUFx2_ASAP7_75t_R output3542 (.A(net3542),
    .Y(io_outs_right_6[29]));
 BUFx2_ASAP7_75t_R output3543 (.A(net3543),
    .Y(io_outs_right_6[2]));
 BUFx2_ASAP7_75t_R output3544 (.A(net3544),
    .Y(io_outs_right_6[30]));
 BUFx2_ASAP7_75t_R output3545 (.A(net3545),
    .Y(io_outs_right_6[31]));
 BUFx2_ASAP7_75t_R output3546 (.A(net3546),
    .Y(io_outs_right_6[32]));
 BUFx2_ASAP7_75t_R output3547 (.A(net3547),
    .Y(io_outs_right_6[33]));
 BUFx2_ASAP7_75t_R output3548 (.A(net3548),
    .Y(io_outs_right_6[34]));
 BUFx2_ASAP7_75t_R output3549 (.A(net3549),
    .Y(io_outs_right_6[35]));
 BUFx2_ASAP7_75t_R output3550 (.A(net3550),
    .Y(io_outs_right_6[36]));
 BUFx2_ASAP7_75t_R output3551 (.A(net3551),
    .Y(io_outs_right_6[37]));
 BUFx2_ASAP7_75t_R output3552 (.A(net3552),
    .Y(io_outs_right_6[38]));
 BUFx2_ASAP7_75t_R output3553 (.A(net3553),
    .Y(io_outs_right_6[39]));
 BUFx2_ASAP7_75t_R output3554 (.A(net3554),
    .Y(io_outs_right_6[3]));
 BUFx2_ASAP7_75t_R output3555 (.A(net3555),
    .Y(io_outs_right_6[40]));
 BUFx2_ASAP7_75t_R output3556 (.A(net3556),
    .Y(io_outs_right_6[41]));
 BUFx2_ASAP7_75t_R output3557 (.A(net3557),
    .Y(io_outs_right_6[42]));
 BUFx2_ASAP7_75t_R output3558 (.A(net3558),
    .Y(io_outs_right_6[43]));
 BUFx2_ASAP7_75t_R output3559 (.A(net3559),
    .Y(io_outs_right_6[44]));
 BUFx2_ASAP7_75t_R output3560 (.A(net3560),
    .Y(io_outs_right_6[45]));
 BUFx2_ASAP7_75t_R output3561 (.A(net3561),
    .Y(io_outs_right_6[46]));
 BUFx2_ASAP7_75t_R output3562 (.A(net3562),
    .Y(io_outs_right_6[47]));
 BUFx2_ASAP7_75t_R output3563 (.A(net3563),
    .Y(io_outs_right_6[48]));
 BUFx2_ASAP7_75t_R output3564 (.A(net3564),
    .Y(io_outs_right_6[49]));
 BUFx2_ASAP7_75t_R output3565 (.A(net3565),
    .Y(io_outs_right_6[4]));
 BUFx2_ASAP7_75t_R output3566 (.A(net3566),
    .Y(io_outs_right_6[50]));
 BUFx2_ASAP7_75t_R output3567 (.A(net3567),
    .Y(io_outs_right_6[51]));
 BUFx2_ASAP7_75t_R output3568 (.A(net3568),
    .Y(io_outs_right_6[52]));
 BUFx2_ASAP7_75t_R output3569 (.A(net3569),
    .Y(io_outs_right_6[53]));
 BUFx2_ASAP7_75t_R output3570 (.A(net3570),
    .Y(io_outs_right_6[54]));
 BUFx2_ASAP7_75t_R output3571 (.A(net3571),
    .Y(io_outs_right_6[55]));
 BUFx2_ASAP7_75t_R output3572 (.A(net3572),
    .Y(io_outs_right_6[56]));
 BUFx2_ASAP7_75t_R output3573 (.A(net3573),
    .Y(io_outs_right_6[57]));
 BUFx2_ASAP7_75t_R output3574 (.A(net3574),
    .Y(io_outs_right_6[58]));
 BUFx2_ASAP7_75t_R output3575 (.A(net3575),
    .Y(io_outs_right_6[59]));
 BUFx2_ASAP7_75t_R output3576 (.A(net3576),
    .Y(io_outs_right_6[5]));
 BUFx2_ASAP7_75t_R output3577 (.A(net3577),
    .Y(io_outs_right_6[60]));
 BUFx2_ASAP7_75t_R output3578 (.A(net3578),
    .Y(io_outs_right_6[61]));
 BUFx2_ASAP7_75t_R output3579 (.A(net3579),
    .Y(io_outs_right_6[62]));
 BUFx2_ASAP7_75t_R output3580 (.A(net3580),
    .Y(io_outs_right_6[63]));
 BUFx2_ASAP7_75t_R output3581 (.A(net3581),
    .Y(io_outs_right_6[6]));
 BUFx2_ASAP7_75t_R output3582 (.A(net3582),
    .Y(io_outs_right_6[7]));
 BUFx2_ASAP7_75t_R output3583 (.A(net3583),
    .Y(io_outs_right_6[8]));
 BUFx2_ASAP7_75t_R output3584 (.A(net3584),
    .Y(io_outs_right_6[9]));
 BUFx2_ASAP7_75t_R output3585 (.A(net3585),
    .Y(io_outs_right_7[0]));
 BUFx2_ASAP7_75t_R output3586 (.A(net3586),
    .Y(io_outs_right_7[10]));
 BUFx2_ASAP7_75t_R output3587 (.A(net3587),
    .Y(io_outs_right_7[11]));
 BUFx2_ASAP7_75t_R output3588 (.A(net3588),
    .Y(io_outs_right_7[12]));
 BUFx2_ASAP7_75t_R output3589 (.A(net3589),
    .Y(io_outs_right_7[13]));
 BUFx2_ASAP7_75t_R output3590 (.A(net3590),
    .Y(io_outs_right_7[14]));
 BUFx2_ASAP7_75t_R output3591 (.A(net3591),
    .Y(io_outs_right_7[15]));
 BUFx2_ASAP7_75t_R output3592 (.A(net3592),
    .Y(io_outs_right_7[16]));
 BUFx2_ASAP7_75t_R output3593 (.A(net3593),
    .Y(io_outs_right_7[17]));
 BUFx2_ASAP7_75t_R output3594 (.A(net3594),
    .Y(io_outs_right_7[18]));
 BUFx2_ASAP7_75t_R output3595 (.A(net3595),
    .Y(io_outs_right_7[19]));
 BUFx2_ASAP7_75t_R output3596 (.A(net3596),
    .Y(io_outs_right_7[1]));
 BUFx2_ASAP7_75t_R output3597 (.A(net3597),
    .Y(io_outs_right_7[20]));
 BUFx2_ASAP7_75t_R output3598 (.A(net3598),
    .Y(io_outs_right_7[21]));
 BUFx2_ASAP7_75t_R output3599 (.A(net3599),
    .Y(io_outs_right_7[22]));
 BUFx2_ASAP7_75t_R output3600 (.A(net3600),
    .Y(io_outs_right_7[23]));
 BUFx2_ASAP7_75t_R output3601 (.A(net3601),
    .Y(io_outs_right_7[24]));
 BUFx2_ASAP7_75t_R output3602 (.A(net3602),
    .Y(io_outs_right_7[25]));
 BUFx2_ASAP7_75t_R output3603 (.A(net3603),
    .Y(io_outs_right_7[26]));
 BUFx2_ASAP7_75t_R output3604 (.A(net3604),
    .Y(io_outs_right_7[27]));
 BUFx2_ASAP7_75t_R output3605 (.A(net3605),
    .Y(io_outs_right_7[28]));
 BUFx2_ASAP7_75t_R output3606 (.A(net3606),
    .Y(io_outs_right_7[29]));
 BUFx2_ASAP7_75t_R output3607 (.A(net3607),
    .Y(io_outs_right_7[2]));
 BUFx2_ASAP7_75t_R output3608 (.A(net3608),
    .Y(io_outs_right_7[30]));
 BUFx2_ASAP7_75t_R output3609 (.A(net3609),
    .Y(io_outs_right_7[31]));
 BUFx2_ASAP7_75t_R output3610 (.A(net3610),
    .Y(io_outs_right_7[32]));
 BUFx2_ASAP7_75t_R output3611 (.A(net3611),
    .Y(io_outs_right_7[33]));
 BUFx2_ASAP7_75t_R output3612 (.A(net3612),
    .Y(io_outs_right_7[34]));
 BUFx2_ASAP7_75t_R output3613 (.A(net3613),
    .Y(io_outs_right_7[35]));
 BUFx2_ASAP7_75t_R output3614 (.A(net3614),
    .Y(io_outs_right_7[36]));
 BUFx2_ASAP7_75t_R output3615 (.A(net3615),
    .Y(io_outs_right_7[37]));
 BUFx2_ASAP7_75t_R output3616 (.A(net3616),
    .Y(io_outs_right_7[38]));
 BUFx2_ASAP7_75t_R output3617 (.A(net3617),
    .Y(io_outs_right_7[39]));
 BUFx2_ASAP7_75t_R output3618 (.A(net3618),
    .Y(io_outs_right_7[3]));
 BUFx2_ASAP7_75t_R output3619 (.A(net3619),
    .Y(io_outs_right_7[40]));
 BUFx2_ASAP7_75t_R output3620 (.A(net3620),
    .Y(io_outs_right_7[41]));
 BUFx2_ASAP7_75t_R output3621 (.A(net3621),
    .Y(io_outs_right_7[42]));
 BUFx2_ASAP7_75t_R output3622 (.A(net3622),
    .Y(io_outs_right_7[43]));
 BUFx2_ASAP7_75t_R output3623 (.A(net3623),
    .Y(io_outs_right_7[44]));
 BUFx2_ASAP7_75t_R output3624 (.A(net3624),
    .Y(io_outs_right_7[45]));
 BUFx2_ASAP7_75t_R output3625 (.A(net3625),
    .Y(io_outs_right_7[46]));
 BUFx2_ASAP7_75t_R output3626 (.A(net3626),
    .Y(io_outs_right_7[47]));
 BUFx2_ASAP7_75t_R output3627 (.A(net3627),
    .Y(io_outs_right_7[48]));
 BUFx2_ASAP7_75t_R output3628 (.A(net3628),
    .Y(io_outs_right_7[49]));
 BUFx2_ASAP7_75t_R output3629 (.A(net3629),
    .Y(io_outs_right_7[4]));
 BUFx2_ASAP7_75t_R output3630 (.A(net3630),
    .Y(io_outs_right_7[50]));
 BUFx2_ASAP7_75t_R output3631 (.A(net3631),
    .Y(io_outs_right_7[51]));
 BUFx2_ASAP7_75t_R output3632 (.A(net3632),
    .Y(io_outs_right_7[52]));
 BUFx2_ASAP7_75t_R output3633 (.A(net3633),
    .Y(io_outs_right_7[53]));
 BUFx2_ASAP7_75t_R output3634 (.A(net3634),
    .Y(io_outs_right_7[54]));
 BUFx2_ASAP7_75t_R output3635 (.A(net3635),
    .Y(io_outs_right_7[55]));
 BUFx2_ASAP7_75t_R output3636 (.A(net3636),
    .Y(io_outs_right_7[56]));
 BUFx2_ASAP7_75t_R output3637 (.A(net3637),
    .Y(io_outs_right_7[57]));
 BUFx2_ASAP7_75t_R output3638 (.A(net3638),
    .Y(io_outs_right_7[58]));
 BUFx2_ASAP7_75t_R output3639 (.A(net3639),
    .Y(io_outs_right_7[59]));
 BUFx2_ASAP7_75t_R output3640 (.A(net3640),
    .Y(io_outs_right_7[5]));
 BUFx2_ASAP7_75t_R output3641 (.A(net3641),
    .Y(io_outs_right_7[60]));
 BUFx2_ASAP7_75t_R output3642 (.A(net3642),
    .Y(io_outs_right_7[61]));
 BUFx2_ASAP7_75t_R output3643 (.A(net3643),
    .Y(io_outs_right_7[62]));
 BUFx2_ASAP7_75t_R output3644 (.A(net3644),
    .Y(io_outs_right_7[63]));
 BUFx2_ASAP7_75t_R output3645 (.A(net3645),
    .Y(io_outs_right_7[6]));
 BUFx2_ASAP7_75t_R output3646 (.A(net3646),
    .Y(io_outs_right_7[7]));
 BUFx2_ASAP7_75t_R output3647 (.A(net3647),
    .Y(io_outs_right_7[8]));
 BUFx2_ASAP7_75t_R output3648 (.A(net3648),
    .Y(io_outs_right_7[9]));
 BUFx2_ASAP7_75t_R output3649 (.A(net3649),
    .Y(io_outs_up_0[0]));
 BUFx2_ASAP7_75t_R output3650 (.A(net3650),
    .Y(io_outs_up_0[10]));
 BUFx2_ASAP7_75t_R output3651 (.A(net3651),
    .Y(io_outs_up_0[11]));
 BUFx2_ASAP7_75t_R output3652 (.A(net3652),
    .Y(io_outs_up_0[12]));
 BUFx2_ASAP7_75t_R output3653 (.A(net3653),
    .Y(io_outs_up_0[13]));
 BUFx2_ASAP7_75t_R output3654 (.A(net3654),
    .Y(io_outs_up_0[14]));
 BUFx2_ASAP7_75t_R output3655 (.A(net3655),
    .Y(io_outs_up_0[15]));
 BUFx2_ASAP7_75t_R output3656 (.A(net3656),
    .Y(io_outs_up_0[16]));
 BUFx2_ASAP7_75t_R output3657 (.A(net3657),
    .Y(io_outs_up_0[17]));
 BUFx2_ASAP7_75t_R output3658 (.A(net3658),
    .Y(io_outs_up_0[18]));
 BUFx2_ASAP7_75t_R output3659 (.A(net3659),
    .Y(io_outs_up_0[19]));
 BUFx2_ASAP7_75t_R output3660 (.A(net3660),
    .Y(io_outs_up_0[1]));
 BUFx2_ASAP7_75t_R output3661 (.A(net3661),
    .Y(io_outs_up_0[20]));
 BUFx2_ASAP7_75t_R output3662 (.A(net3662),
    .Y(io_outs_up_0[21]));
 BUFx2_ASAP7_75t_R output3663 (.A(net3663),
    .Y(io_outs_up_0[22]));
 BUFx2_ASAP7_75t_R output3664 (.A(net3664),
    .Y(io_outs_up_0[23]));
 BUFx2_ASAP7_75t_R output3665 (.A(net3665),
    .Y(io_outs_up_0[24]));
 BUFx2_ASAP7_75t_R output3666 (.A(net3666),
    .Y(io_outs_up_0[25]));
 BUFx2_ASAP7_75t_R output3667 (.A(net3667),
    .Y(io_outs_up_0[26]));
 BUFx2_ASAP7_75t_R output3668 (.A(net3668),
    .Y(io_outs_up_0[27]));
 BUFx2_ASAP7_75t_R output3669 (.A(net3669),
    .Y(io_outs_up_0[28]));
 BUFx2_ASAP7_75t_R output3670 (.A(net3670),
    .Y(io_outs_up_0[29]));
 BUFx2_ASAP7_75t_R output3671 (.A(net3671),
    .Y(io_outs_up_0[2]));
 BUFx2_ASAP7_75t_R output3672 (.A(net3672),
    .Y(io_outs_up_0[30]));
 BUFx2_ASAP7_75t_R output3673 (.A(net3673),
    .Y(io_outs_up_0[31]));
 BUFx2_ASAP7_75t_R output3674 (.A(net3674),
    .Y(io_outs_up_0[32]));
 BUFx2_ASAP7_75t_R output3675 (.A(net3675),
    .Y(io_outs_up_0[33]));
 BUFx2_ASAP7_75t_R output3676 (.A(net3676),
    .Y(io_outs_up_0[34]));
 BUFx2_ASAP7_75t_R output3677 (.A(net3677),
    .Y(io_outs_up_0[35]));
 BUFx2_ASAP7_75t_R output3678 (.A(net3678),
    .Y(io_outs_up_0[36]));
 BUFx2_ASAP7_75t_R output3679 (.A(net3679),
    .Y(io_outs_up_0[37]));
 BUFx2_ASAP7_75t_R output3680 (.A(net3680),
    .Y(io_outs_up_0[38]));
 BUFx2_ASAP7_75t_R output3681 (.A(net3681),
    .Y(io_outs_up_0[39]));
 BUFx2_ASAP7_75t_R output3682 (.A(net3682),
    .Y(io_outs_up_0[3]));
 BUFx2_ASAP7_75t_R output3683 (.A(net3683),
    .Y(io_outs_up_0[40]));
 BUFx2_ASAP7_75t_R output3684 (.A(net3684),
    .Y(io_outs_up_0[41]));
 BUFx2_ASAP7_75t_R output3685 (.A(net3685),
    .Y(io_outs_up_0[42]));
 BUFx2_ASAP7_75t_R output3686 (.A(net3686),
    .Y(io_outs_up_0[43]));
 BUFx2_ASAP7_75t_R output3687 (.A(net3687),
    .Y(io_outs_up_0[44]));
 BUFx2_ASAP7_75t_R output3688 (.A(net3688),
    .Y(io_outs_up_0[45]));
 BUFx2_ASAP7_75t_R output3689 (.A(net3689),
    .Y(io_outs_up_0[46]));
 BUFx2_ASAP7_75t_R output3690 (.A(net3690),
    .Y(io_outs_up_0[47]));
 BUFx2_ASAP7_75t_R output3691 (.A(net3691),
    .Y(io_outs_up_0[48]));
 BUFx2_ASAP7_75t_R output3692 (.A(net3692),
    .Y(io_outs_up_0[49]));
 BUFx2_ASAP7_75t_R output3693 (.A(net3693),
    .Y(io_outs_up_0[4]));
 BUFx2_ASAP7_75t_R output3694 (.A(net3694),
    .Y(io_outs_up_0[50]));
 BUFx2_ASAP7_75t_R output3695 (.A(net3695),
    .Y(io_outs_up_0[51]));
 BUFx2_ASAP7_75t_R output3696 (.A(net3696),
    .Y(io_outs_up_0[52]));
 BUFx2_ASAP7_75t_R output3697 (.A(net3697),
    .Y(io_outs_up_0[53]));
 BUFx2_ASAP7_75t_R output3698 (.A(net3698),
    .Y(io_outs_up_0[54]));
 BUFx2_ASAP7_75t_R output3699 (.A(net3699),
    .Y(io_outs_up_0[55]));
 BUFx2_ASAP7_75t_R output3700 (.A(net3700),
    .Y(io_outs_up_0[56]));
 BUFx2_ASAP7_75t_R output3701 (.A(net3701),
    .Y(io_outs_up_0[57]));
 BUFx2_ASAP7_75t_R output3702 (.A(net3702),
    .Y(io_outs_up_0[58]));
 BUFx2_ASAP7_75t_R output3703 (.A(net3703),
    .Y(io_outs_up_0[59]));
 BUFx2_ASAP7_75t_R output3704 (.A(net3704),
    .Y(io_outs_up_0[5]));
 BUFx2_ASAP7_75t_R output3705 (.A(net3705),
    .Y(io_outs_up_0[60]));
 BUFx2_ASAP7_75t_R output3706 (.A(net3706),
    .Y(io_outs_up_0[61]));
 BUFx2_ASAP7_75t_R output3707 (.A(net3707),
    .Y(io_outs_up_0[62]));
 BUFx2_ASAP7_75t_R output3708 (.A(net3708),
    .Y(io_outs_up_0[63]));
 BUFx2_ASAP7_75t_R output3709 (.A(net3709),
    .Y(io_outs_up_0[6]));
 BUFx2_ASAP7_75t_R output3710 (.A(net3710),
    .Y(io_outs_up_0[7]));
 BUFx2_ASAP7_75t_R output3711 (.A(net3711),
    .Y(io_outs_up_0[8]));
 BUFx2_ASAP7_75t_R output3712 (.A(net3712),
    .Y(io_outs_up_0[9]));
 BUFx2_ASAP7_75t_R output3713 (.A(net3713),
    .Y(io_outs_up_1[0]));
 BUFx2_ASAP7_75t_R output3714 (.A(net3714),
    .Y(io_outs_up_1[10]));
 BUFx2_ASAP7_75t_R output3715 (.A(net3715),
    .Y(io_outs_up_1[11]));
 BUFx2_ASAP7_75t_R output3716 (.A(net3716),
    .Y(io_outs_up_1[12]));
 BUFx2_ASAP7_75t_R output3717 (.A(net3717),
    .Y(io_outs_up_1[13]));
 BUFx2_ASAP7_75t_R output3718 (.A(net3718),
    .Y(io_outs_up_1[14]));
 BUFx2_ASAP7_75t_R output3719 (.A(net3719),
    .Y(io_outs_up_1[15]));
 BUFx2_ASAP7_75t_R output3720 (.A(net3720),
    .Y(io_outs_up_1[16]));
 BUFx2_ASAP7_75t_R output3721 (.A(net3721),
    .Y(io_outs_up_1[17]));
 BUFx2_ASAP7_75t_R output3722 (.A(net3722),
    .Y(io_outs_up_1[18]));
 BUFx2_ASAP7_75t_R output3723 (.A(net3723),
    .Y(io_outs_up_1[19]));
 BUFx2_ASAP7_75t_R output3724 (.A(net3724),
    .Y(io_outs_up_1[1]));
 BUFx2_ASAP7_75t_R output3725 (.A(net3725),
    .Y(io_outs_up_1[20]));
 BUFx2_ASAP7_75t_R output3726 (.A(net3726),
    .Y(io_outs_up_1[21]));
 BUFx2_ASAP7_75t_R output3727 (.A(net3727),
    .Y(io_outs_up_1[22]));
 BUFx2_ASAP7_75t_R output3728 (.A(net3728),
    .Y(io_outs_up_1[23]));
 BUFx2_ASAP7_75t_R output3729 (.A(net3729),
    .Y(io_outs_up_1[24]));
 BUFx2_ASAP7_75t_R output3730 (.A(net3730),
    .Y(io_outs_up_1[25]));
 BUFx2_ASAP7_75t_R output3731 (.A(net3731),
    .Y(io_outs_up_1[26]));
 BUFx2_ASAP7_75t_R output3732 (.A(net3732),
    .Y(io_outs_up_1[27]));
 BUFx2_ASAP7_75t_R output3733 (.A(net3733),
    .Y(io_outs_up_1[28]));
 BUFx2_ASAP7_75t_R output3734 (.A(net3734),
    .Y(io_outs_up_1[29]));
 BUFx2_ASAP7_75t_R output3735 (.A(net3735),
    .Y(io_outs_up_1[2]));
 BUFx2_ASAP7_75t_R output3736 (.A(net3736),
    .Y(io_outs_up_1[30]));
 BUFx2_ASAP7_75t_R output3737 (.A(net3737),
    .Y(io_outs_up_1[31]));
 BUFx2_ASAP7_75t_R output3738 (.A(net3738),
    .Y(io_outs_up_1[32]));
 BUFx2_ASAP7_75t_R output3739 (.A(net3739),
    .Y(io_outs_up_1[33]));
 BUFx2_ASAP7_75t_R output3740 (.A(net3740),
    .Y(io_outs_up_1[34]));
 BUFx2_ASAP7_75t_R output3741 (.A(net3741),
    .Y(io_outs_up_1[35]));
 BUFx2_ASAP7_75t_R output3742 (.A(net3742),
    .Y(io_outs_up_1[36]));
 BUFx2_ASAP7_75t_R output3743 (.A(net3743),
    .Y(io_outs_up_1[37]));
 BUFx2_ASAP7_75t_R output3744 (.A(net3744),
    .Y(io_outs_up_1[38]));
 BUFx2_ASAP7_75t_R output3745 (.A(net3745),
    .Y(io_outs_up_1[39]));
 BUFx2_ASAP7_75t_R output3746 (.A(net3746),
    .Y(io_outs_up_1[3]));
 BUFx2_ASAP7_75t_R output3747 (.A(net3747),
    .Y(io_outs_up_1[40]));
 BUFx2_ASAP7_75t_R output3748 (.A(net3748),
    .Y(io_outs_up_1[41]));
 BUFx2_ASAP7_75t_R output3749 (.A(net3749),
    .Y(io_outs_up_1[42]));
 BUFx2_ASAP7_75t_R output3750 (.A(net3750),
    .Y(io_outs_up_1[43]));
 BUFx2_ASAP7_75t_R output3751 (.A(net3751),
    .Y(io_outs_up_1[44]));
 BUFx2_ASAP7_75t_R output3752 (.A(net3752),
    .Y(io_outs_up_1[45]));
 BUFx2_ASAP7_75t_R output3753 (.A(net3753),
    .Y(io_outs_up_1[46]));
 BUFx2_ASAP7_75t_R output3754 (.A(net3754),
    .Y(io_outs_up_1[47]));
 BUFx2_ASAP7_75t_R output3755 (.A(net3755),
    .Y(io_outs_up_1[48]));
 BUFx2_ASAP7_75t_R output3756 (.A(net3756),
    .Y(io_outs_up_1[49]));
 BUFx2_ASAP7_75t_R output3757 (.A(net3757),
    .Y(io_outs_up_1[4]));
 BUFx2_ASAP7_75t_R output3758 (.A(net3758),
    .Y(io_outs_up_1[50]));
 BUFx2_ASAP7_75t_R output3759 (.A(net3759),
    .Y(io_outs_up_1[51]));
 BUFx2_ASAP7_75t_R output3760 (.A(net3760),
    .Y(io_outs_up_1[52]));
 BUFx2_ASAP7_75t_R output3761 (.A(net3761),
    .Y(io_outs_up_1[53]));
 BUFx2_ASAP7_75t_R output3762 (.A(net3762),
    .Y(io_outs_up_1[54]));
 BUFx2_ASAP7_75t_R output3763 (.A(net3763),
    .Y(io_outs_up_1[55]));
 BUFx2_ASAP7_75t_R output3764 (.A(net3764),
    .Y(io_outs_up_1[56]));
 BUFx2_ASAP7_75t_R output3765 (.A(net3765),
    .Y(io_outs_up_1[57]));
 BUFx2_ASAP7_75t_R output3766 (.A(net3766),
    .Y(io_outs_up_1[58]));
 BUFx2_ASAP7_75t_R output3767 (.A(net3767),
    .Y(io_outs_up_1[59]));
 BUFx2_ASAP7_75t_R output3768 (.A(net3768),
    .Y(io_outs_up_1[5]));
 BUFx2_ASAP7_75t_R output3769 (.A(net3769),
    .Y(io_outs_up_1[60]));
 BUFx2_ASAP7_75t_R output3770 (.A(net3770),
    .Y(io_outs_up_1[61]));
 BUFx2_ASAP7_75t_R output3771 (.A(net3771),
    .Y(io_outs_up_1[62]));
 BUFx2_ASAP7_75t_R output3772 (.A(net3772),
    .Y(io_outs_up_1[63]));
 BUFx2_ASAP7_75t_R output3773 (.A(net3773),
    .Y(io_outs_up_1[6]));
 BUFx2_ASAP7_75t_R output3774 (.A(net3774),
    .Y(io_outs_up_1[7]));
 BUFx2_ASAP7_75t_R output3775 (.A(net3775),
    .Y(io_outs_up_1[8]));
 BUFx2_ASAP7_75t_R output3776 (.A(net3776),
    .Y(io_outs_up_1[9]));
 BUFx2_ASAP7_75t_R output3777 (.A(net3777),
    .Y(io_outs_up_2[0]));
 BUFx2_ASAP7_75t_R output3778 (.A(net3778),
    .Y(io_outs_up_2[10]));
 BUFx2_ASAP7_75t_R output3779 (.A(net3779),
    .Y(io_outs_up_2[11]));
 BUFx2_ASAP7_75t_R output3780 (.A(net3780),
    .Y(io_outs_up_2[12]));
 BUFx2_ASAP7_75t_R output3781 (.A(net3781),
    .Y(io_outs_up_2[13]));
 BUFx2_ASAP7_75t_R output3782 (.A(net3782),
    .Y(io_outs_up_2[14]));
 BUFx2_ASAP7_75t_R output3783 (.A(net3783),
    .Y(io_outs_up_2[15]));
 BUFx2_ASAP7_75t_R output3784 (.A(net3784),
    .Y(io_outs_up_2[16]));
 BUFx2_ASAP7_75t_R output3785 (.A(net3785),
    .Y(io_outs_up_2[17]));
 BUFx2_ASAP7_75t_R output3786 (.A(net3786),
    .Y(io_outs_up_2[18]));
 BUFx2_ASAP7_75t_R output3787 (.A(net3787),
    .Y(io_outs_up_2[19]));
 BUFx2_ASAP7_75t_R output3788 (.A(net3788),
    .Y(io_outs_up_2[1]));
 BUFx2_ASAP7_75t_R output3789 (.A(net3789),
    .Y(io_outs_up_2[20]));
 BUFx2_ASAP7_75t_R output3790 (.A(net3790),
    .Y(io_outs_up_2[21]));
 BUFx2_ASAP7_75t_R output3791 (.A(net3791),
    .Y(io_outs_up_2[22]));
 BUFx2_ASAP7_75t_R output3792 (.A(net3792),
    .Y(io_outs_up_2[23]));
 BUFx2_ASAP7_75t_R output3793 (.A(net3793),
    .Y(io_outs_up_2[24]));
 BUFx2_ASAP7_75t_R output3794 (.A(net3794),
    .Y(io_outs_up_2[25]));
 BUFx2_ASAP7_75t_R output3795 (.A(net3795),
    .Y(io_outs_up_2[26]));
 BUFx2_ASAP7_75t_R output3796 (.A(net3796),
    .Y(io_outs_up_2[27]));
 BUFx2_ASAP7_75t_R output3797 (.A(net3797),
    .Y(io_outs_up_2[28]));
 BUFx2_ASAP7_75t_R output3798 (.A(net3798),
    .Y(io_outs_up_2[29]));
 BUFx2_ASAP7_75t_R output3799 (.A(net3799),
    .Y(io_outs_up_2[2]));
 BUFx2_ASAP7_75t_R output3800 (.A(net3800),
    .Y(io_outs_up_2[30]));
 BUFx2_ASAP7_75t_R output3801 (.A(net3801),
    .Y(io_outs_up_2[31]));
 BUFx2_ASAP7_75t_R output3802 (.A(net3802),
    .Y(io_outs_up_2[32]));
 BUFx2_ASAP7_75t_R output3803 (.A(net3803),
    .Y(io_outs_up_2[33]));
 BUFx2_ASAP7_75t_R output3804 (.A(net3804),
    .Y(io_outs_up_2[34]));
 BUFx2_ASAP7_75t_R output3805 (.A(net3805),
    .Y(io_outs_up_2[35]));
 BUFx2_ASAP7_75t_R output3806 (.A(net3806),
    .Y(io_outs_up_2[36]));
 BUFx2_ASAP7_75t_R output3807 (.A(net3807),
    .Y(io_outs_up_2[37]));
 BUFx2_ASAP7_75t_R output3808 (.A(net3808),
    .Y(io_outs_up_2[38]));
 BUFx2_ASAP7_75t_R output3809 (.A(net3809),
    .Y(io_outs_up_2[39]));
 BUFx2_ASAP7_75t_R output3810 (.A(net3810),
    .Y(io_outs_up_2[3]));
 BUFx2_ASAP7_75t_R output3811 (.A(net3811),
    .Y(io_outs_up_2[40]));
 BUFx2_ASAP7_75t_R output3812 (.A(net3812),
    .Y(io_outs_up_2[41]));
 BUFx2_ASAP7_75t_R output3813 (.A(net3813),
    .Y(io_outs_up_2[42]));
 BUFx2_ASAP7_75t_R output3814 (.A(net3814),
    .Y(io_outs_up_2[43]));
 BUFx2_ASAP7_75t_R output3815 (.A(net3815),
    .Y(io_outs_up_2[44]));
 BUFx2_ASAP7_75t_R output3816 (.A(net3816),
    .Y(io_outs_up_2[45]));
 BUFx2_ASAP7_75t_R output3817 (.A(net3817),
    .Y(io_outs_up_2[46]));
 BUFx2_ASAP7_75t_R output3818 (.A(net3818),
    .Y(io_outs_up_2[47]));
 BUFx2_ASAP7_75t_R output3819 (.A(net3819),
    .Y(io_outs_up_2[48]));
 BUFx2_ASAP7_75t_R output3820 (.A(net3820),
    .Y(io_outs_up_2[49]));
 BUFx2_ASAP7_75t_R output3821 (.A(net3821),
    .Y(io_outs_up_2[4]));
 BUFx2_ASAP7_75t_R output3822 (.A(net3822),
    .Y(io_outs_up_2[50]));
 BUFx2_ASAP7_75t_R output3823 (.A(net3823),
    .Y(io_outs_up_2[51]));
 BUFx2_ASAP7_75t_R output3824 (.A(net3824),
    .Y(io_outs_up_2[52]));
 BUFx2_ASAP7_75t_R output3825 (.A(net3825),
    .Y(io_outs_up_2[53]));
 BUFx2_ASAP7_75t_R output3826 (.A(net3826),
    .Y(io_outs_up_2[54]));
 BUFx2_ASAP7_75t_R output3827 (.A(net3827),
    .Y(io_outs_up_2[55]));
 BUFx2_ASAP7_75t_R output3828 (.A(net3828),
    .Y(io_outs_up_2[56]));
 BUFx2_ASAP7_75t_R output3829 (.A(net3829),
    .Y(io_outs_up_2[57]));
 BUFx2_ASAP7_75t_R output3830 (.A(net3830),
    .Y(io_outs_up_2[58]));
 BUFx2_ASAP7_75t_R output3831 (.A(net3831),
    .Y(io_outs_up_2[59]));
 BUFx2_ASAP7_75t_R output3832 (.A(net3832),
    .Y(io_outs_up_2[5]));
 BUFx2_ASAP7_75t_R output3833 (.A(net3833),
    .Y(io_outs_up_2[60]));
 BUFx2_ASAP7_75t_R output3834 (.A(net3834),
    .Y(io_outs_up_2[61]));
 BUFx2_ASAP7_75t_R output3835 (.A(net3835),
    .Y(io_outs_up_2[62]));
 BUFx2_ASAP7_75t_R output3836 (.A(net3836),
    .Y(io_outs_up_2[63]));
 BUFx2_ASAP7_75t_R output3837 (.A(net3837),
    .Y(io_outs_up_2[6]));
 BUFx2_ASAP7_75t_R output3838 (.A(net3838),
    .Y(io_outs_up_2[7]));
 BUFx2_ASAP7_75t_R output3839 (.A(net3839),
    .Y(io_outs_up_2[8]));
 BUFx2_ASAP7_75t_R output3840 (.A(net3840),
    .Y(io_outs_up_2[9]));
 BUFx2_ASAP7_75t_R output3841 (.A(net3841),
    .Y(io_outs_up_3[0]));
 BUFx2_ASAP7_75t_R output3842 (.A(net3842),
    .Y(io_outs_up_3[10]));
 BUFx2_ASAP7_75t_R output3843 (.A(net3843),
    .Y(io_outs_up_3[11]));
 BUFx2_ASAP7_75t_R output3844 (.A(net3844),
    .Y(io_outs_up_3[12]));
 BUFx2_ASAP7_75t_R output3845 (.A(net3845),
    .Y(io_outs_up_3[13]));
 BUFx2_ASAP7_75t_R output3846 (.A(net3846),
    .Y(io_outs_up_3[14]));
 BUFx2_ASAP7_75t_R output3847 (.A(net3847),
    .Y(io_outs_up_3[15]));
 BUFx2_ASAP7_75t_R output3848 (.A(net3848),
    .Y(io_outs_up_3[16]));
 BUFx2_ASAP7_75t_R output3849 (.A(net3849),
    .Y(io_outs_up_3[17]));
 BUFx2_ASAP7_75t_R output3850 (.A(net3850),
    .Y(io_outs_up_3[18]));
 BUFx2_ASAP7_75t_R output3851 (.A(net3851),
    .Y(io_outs_up_3[19]));
 BUFx2_ASAP7_75t_R output3852 (.A(net3852),
    .Y(io_outs_up_3[1]));
 BUFx2_ASAP7_75t_R output3853 (.A(net3853),
    .Y(io_outs_up_3[20]));
 BUFx2_ASAP7_75t_R output3854 (.A(net3854),
    .Y(io_outs_up_3[21]));
 BUFx2_ASAP7_75t_R output3855 (.A(net3855),
    .Y(io_outs_up_3[22]));
 BUFx2_ASAP7_75t_R output3856 (.A(net3856),
    .Y(io_outs_up_3[23]));
 BUFx2_ASAP7_75t_R output3857 (.A(net3857),
    .Y(io_outs_up_3[24]));
 BUFx2_ASAP7_75t_R output3858 (.A(net3858),
    .Y(io_outs_up_3[25]));
 BUFx2_ASAP7_75t_R output3859 (.A(net3859),
    .Y(io_outs_up_3[26]));
 BUFx2_ASAP7_75t_R output3860 (.A(net3860),
    .Y(io_outs_up_3[27]));
 BUFx2_ASAP7_75t_R output3861 (.A(net3861),
    .Y(io_outs_up_3[28]));
 BUFx2_ASAP7_75t_R output3862 (.A(net3862),
    .Y(io_outs_up_3[29]));
 BUFx2_ASAP7_75t_R output3863 (.A(net3863),
    .Y(io_outs_up_3[2]));
 BUFx2_ASAP7_75t_R output3864 (.A(net3864),
    .Y(io_outs_up_3[30]));
 BUFx2_ASAP7_75t_R output3865 (.A(net3865),
    .Y(io_outs_up_3[31]));
 BUFx2_ASAP7_75t_R output3866 (.A(net3866),
    .Y(io_outs_up_3[32]));
 BUFx2_ASAP7_75t_R output3867 (.A(net3867),
    .Y(io_outs_up_3[33]));
 BUFx2_ASAP7_75t_R output3868 (.A(net3868),
    .Y(io_outs_up_3[34]));
 BUFx2_ASAP7_75t_R output3869 (.A(net3869),
    .Y(io_outs_up_3[35]));
 BUFx2_ASAP7_75t_R output3870 (.A(net3870),
    .Y(io_outs_up_3[36]));
 BUFx2_ASAP7_75t_R output3871 (.A(net3871),
    .Y(io_outs_up_3[37]));
 BUFx2_ASAP7_75t_R output3872 (.A(net3872),
    .Y(io_outs_up_3[38]));
 BUFx2_ASAP7_75t_R output3873 (.A(net3873),
    .Y(io_outs_up_3[39]));
 BUFx2_ASAP7_75t_R output3874 (.A(net3874),
    .Y(io_outs_up_3[3]));
 BUFx2_ASAP7_75t_R output3875 (.A(net3875),
    .Y(io_outs_up_3[40]));
 BUFx2_ASAP7_75t_R output3876 (.A(net3876),
    .Y(io_outs_up_3[41]));
 BUFx2_ASAP7_75t_R output3877 (.A(net3877),
    .Y(io_outs_up_3[42]));
 BUFx2_ASAP7_75t_R output3878 (.A(net3878),
    .Y(io_outs_up_3[43]));
 BUFx2_ASAP7_75t_R output3879 (.A(net3879),
    .Y(io_outs_up_3[44]));
 BUFx2_ASAP7_75t_R output3880 (.A(net3880),
    .Y(io_outs_up_3[45]));
 BUFx2_ASAP7_75t_R output3881 (.A(net3881),
    .Y(io_outs_up_3[46]));
 BUFx2_ASAP7_75t_R output3882 (.A(net3882),
    .Y(io_outs_up_3[47]));
 BUFx2_ASAP7_75t_R output3883 (.A(net3883),
    .Y(io_outs_up_3[48]));
 BUFx2_ASAP7_75t_R output3884 (.A(net3884),
    .Y(io_outs_up_3[49]));
 BUFx2_ASAP7_75t_R output3885 (.A(net3885),
    .Y(io_outs_up_3[4]));
 BUFx2_ASAP7_75t_R output3886 (.A(net3886),
    .Y(io_outs_up_3[50]));
 BUFx2_ASAP7_75t_R output3887 (.A(net3887),
    .Y(io_outs_up_3[51]));
 BUFx2_ASAP7_75t_R output3888 (.A(net3888),
    .Y(io_outs_up_3[52]));
 BUFx2_ASAP7_75t_R output3889 (.A(net3889),
    .Y(io_outs_up_3[53]));
 BUFx2_ASAP7_75t_R output3890 (.A(net3890),
    .Y(io_outs_up_3[54]));
 BUFx2_ASAP7_75t_R output3891 (.A(net3891),
    .Y(io_outs_up_3[55]));
 BUFx2_ASAP7_75t_R output3892 (.A(net3892),
    .Y(io_outs_up_3[56]));
 BUFx2_ASAP7_75t_R output3893 (.A(net3893),
    .Y(io_outs_up_3[57]));
 BUFx2_ASAP7_75t_R output3894 (.A(net3894),
    .Y(io_outs_up_3[58]));
 BUFx2_ASAP7_75t_R output3895 (.A(net3895),
    .Y(io_outs_up_3[59]));
 BUFx2_ASAP7_75t_R output3896 (.A(net3896),
    .Y(io_outs_up_3[5]));
 BUFx2_ASAP7_75t_R output3897 (.A(net3897),
    .Y(io_outs_up_3[60]));
 BUFx2_ASAP7_75t_R output3898 (.A(net3898),
    .Y(io_outs_up_3[61]));
 BUFx2_ASAP7_75t_R output3899 (.A(net3899),
    .Y(io_outs_up_3[62]));
 BUFx2_ASAP7_75t_R output3900 (.A(net3900),
    .Y(io_outs_up_3[63]));
 BUFx2_ASAP7_75t_R output3901 (.A(net3901),
    .Y(io_outs_up_3[6]));
 BUFx2_ASAP7_75t_R output3902 (.A(net3902),
    .Y(io_outs_up_3[7]));
 BUFx2_ASAP7_75t_R output3903 (.A(net3903),
    .Y(io_outs_up_3[8]));
 BUFx2_ASAP7_75t_R output3904 (.A(net3904),
    .Y(io_outs_up_3[9]));
 BUFx2_ASAP7_75t_R output3905 (.A(net3905),
    .Y(io_outs_up_4[0]));
 BUFx2_ASAP7_75t_R output3906 (.A(net3906),
    .Y(io_outs_up_4[10]));
 BUFx2_ASAP7_75t_R output3907 (.A(net3907),
    .Y(io_outs_up_4[11]));
 BUFx2_ASAP7_75t_R output3908 (.A(net3908),
    .Y(io_outs_up_4[12]));
 BUFx2_ASAP7_75t_R output3909 (.A(net3909),
    .Y(io_outs_up_4[13]));
 BUFx2_ASAP7_75t_R output3910 (.A(net3910),
    .Y(io_outs_up_4[14]));
 BUFx2_ASAP7_75t_R output3911 (.A(net3911),
    .Y(io_outs_up_4[15]));
 BUFx2_ASAP7_75t_R output3912 (.A(net3912),
    .Y(io_outs_up_4[16]));
 BUFx2_ASAP7_75t_R output3913 (.A(net3913),
    .Y(io_outs_up_4[17]));
 BUFx2_ASAP7_75t_R output3914 (.A(net3914),
    .Y(io_outs_up_4[18]));
 BUFx2_ASAP7_75t_R output3915 (.A(net3915),
    .Y(io_outs_up_4[19]));
 BUFx2_ASAP7_75t_R output3916 (.A(net3916),
    .Y(io_outs_up_4[1]));
 BUFx2_ASAP7_75t_R output3917 (.A(net3917),
    .Y(io_outs_up_4[20]));
 BUFx2_ASAP7_75t_R output3918 (.A(net3918),
    .Y(io_outs_up_4[21]));
 BUFx2_ASAP7_75t_R output3919 (.A(net3919),
    .Y(io_outs_up_4[22]));
 BUFx2_ASAP7_75t_R output3920 (.A(net3920),
    .Y(io_outs_up_4[23]));
 BUFx2_ASAP7_75t_R output3921 (.A(net3921),
    .Y(io_outs_up_4[24]));
 BUFx2_ASAP7_75t_R output3922 (.A(net3922),
    .Y(io_outs_up_4[25]));
 BUFx2_ASAP7_75t_R output3923 (.A(net3923),
    .Y(io_outs_up_4[26]));
 BUFx2_ASAP7_75t_R output3924 (.A(net3924),
    .Y(io_outs_up_4[27]));
 BUFx2_ASAP7_75t_R output3925 (.A(net3925),
    .Y(io_outs_up_4[28]));
 BUFx2_ASAP7_75t_R output3926 (.A(net3926),
    .Y(io_outs_up_4[29]));
 BUFx2_ASAP7_75t_R output3927 (.A(net3927),
    .Y(io_outs_up_4[2]));
 BUFx2_ASAP7_75t_R output3928 (.A(net3928),
    .Y(io_outs_up_4[30]));
 BUFx2_ASAP7_75t_R output3929 (.A(net3929),
    .Y(io_outs_up_4[31]));
 BUFx2_ASAP7_75t_R output3930 (.A(net3930),
    .Y(io_outs_up_4[32]));
 BUFx2_ASAP7_75t_R output3931 (.A(net3931),
    .Y(io_outs_up_4[33]));
 BUFx2_ASAP7_75t_R output3932 (.A(net3932),
    .Y(io_outs_up_4[34]));
 BUFx2_ASAP7_75t_R output3933 (.A(net3933),
    .Y(io_outs_up_4[35]));
 BUFx2_ASAP7_75t_R output3934 (.A(net3934),
    .Y(io_outs_up_4[36]));
 BUFx2_ASAP7_75t_R output3935 (.A(net3935),
    .Y(io_outs_up_4[37]));
 BUFx2_ASAP7_75t_R output3936 (.A(net3936),
    .Y(io_outs_up_4[38]));
 BUFx2_ASAP7_75t_R output3937 (.A(net3937),
    .Y(io_outs_up_4[39]));
 BUFx2_ASAP7_75t_R output3938 (.A(net3938),
    .Y(io_outs_up_4[3]));
 BUFx2_ASAP7_75t_R output3939 (.A(net3939),
    .Y(io_outs_up_4[40]));
 BUFx2_ASAP7_75t_R output3940 (.A(net3940),
    .Y(io_outs_up_4[41]));
 BUFx2_ASAP7_75t_R output3941 (.A(net3941),
    .Y(io_outs_up_4[42]));
 BUFx2_ASAP7_75t_R output3942 (.A(net3942),
    .Y(io_outs_up_4[43]));
 BUFx2_ASAP7_75t_R output3943 (.A(net3943),
    .Y(io_outs_up_4[44]));
 BUFx2_ASAP7_75t_R output3944 (.A(net3944),
    .Y(io_outs_up_4[45]));
 BUFx2_ASAP7_75t_R output3945 (.A(net3945),
    .Y(io_outs_up_4[46]));
 BUFx2_ASAP7_75t_R output3946 (.A(net3946),
    .Y(io_outs_up_4[47]));
 BUFx2_ASAP7_75t_R output3947 (.A(net3947),
    .Y(io_outs_up_4[48]));
 BUFx2_ASAP7_75t_R output3948 (.A(net3948),
    .Y(io_outs_up_4[49]));
 BUFx2_ASAP7_75t_R output3949 (.A(net3949),
    .Y(io_outs_up_4[4]));
 BUFx2_ASAP7_75t_R output3950 (.A(net3950),
    .Y(io_outs_up_4[50]));
 BUFx2_ASAP7_75t_R output3951 (.A(net3951),
    .Y(io_outs_up_4[51]));
 BUFx2_ASAP7_75t_R output3952 (.A(net3952),
    .Y(io_outs_up_4[52]));
 BUFx2_ASAP7_75t_R output3953 (.A(net3953),
    .Y(io_outs_up_4[53]));
 BUFx2_ASAP7_75t_R output3954 (.A(net3954),
    .Y(io_outs_up_4[54]));
 BUFx2_ASAP7_75t_R output3955 (.A(net3955),
    .Y(io_outs_up_4[55]));
 BUFx2_ASAP7_75t_R output3956 (.A(net3956),
    .Y(io_outs_up_4[56]));
 BUFx2_ASAP7_75t_R output3957 (.A(net3957),
    .Y(io_outs_up_4[57]));
 BUFx2_ASAP7_75t_R output3958 (.A(net3958),
    .Y(io_outs_up_4[58]));
 BUFx2_ASAP7_75t_R output3959 (.A(net3959),
    .Y(io_outs_up_4[59]));
 BUFx2_ASAP7_75t_R output3960 (.A(net3960),
    .Y(io_outs_up_4[5]));
 BUFx2_ASAP7_75t_R output3961 (.A(net3961),
    .Y(io_outs_up_4[60]));
 BUFx2_ASAP7_75t_R output3962 (.A(net3962),
    .Y(io_outs_up_4[61]));
 BUFx2_ASAP7_75t_R output3963 (.A(net3963),
    .Y(io_outs_up_4[62]));
 BUFx2_ASAP7_75t_R output3964 (.A(net3964),
    .Y(io_outs_up_4[63]));
 BUFx2_ASAP7_75t_R output3965 (.A(net3965),
    .Y(io_outs_up_4[6]));
 BUFx2_ASAP7_75t_R output3966 (.A(net3966),
    .Y(io_outs_up_4[7]));
 BUFx2_ASAP7_75t_R output3967 (.A(net3967),
    .Y(io_outs_up_4[8]));
 BUFx2_ASAP7_75t_R output3968 (.A(net3968),
    .Y(io_outs_up_4[9]));
 BUFx2_ASAP7_75t_R output3969 (.A(net3969),
    .Y(io_outs_up_5[0]));
 BUFx2_ASAP7_75t_R output3970 (.A(net3970),
    .Y(io_outs_up_5[10]));
 BUFx2_ASAP7_75t_R output3971 (.A(net3971),
    .Y(io_outs_up_5[11]));
 BUFx2_ASAP7_75t_R output3972 (.A(net3972),
    .Y(io_outs_up_5[12]));
 BUFx2_ASAP7_75t_R output3973 (.A(net3973),
    .Y(io_outs_up_5[13]));
 BUFx2_ASAP7_75t_R output3974 (.A(net3974),
    .Y(io_outs_up_5[14]));
 BUFx2_ASAP7_75t_R output3975 (.A(net3975),
    .Y(io_outs_up_5[15]));
 BUFx2_ASAP7_75t_R output3976 (.A(net3976),
    .Y(io_outs_up_5[16]));
 BUFx2_ASAP7_75t_R output3977 (.A(net3977),
    .Y(io_outs_up_5[17]));
 BUFx2_ASAP7_75t_R output3978 (.A(net3978),
    .Y(io_outs_up_5[18]));
 BUFx2_ASAP7_75t_R output3979 (.A(net3979),
    .Y(io_outs_up_5[19]));
 BUFx2_ASAP7_75t_R output3980 (.A(net3980),
    .Y(io_outs_up_5[1]));
 BUFx2_ASAP7_75t_R output3981 (.A(net3981),
    .Y(io_outs_up_5[20]));
 BUFx2_ASAP7_75t_R output3982 (.A(net3982),
    .Y(io_outs_up_5[21]));
 BUFx2_ASAP7_75t_R output3983 (.A(net3983),
    .Y(io_outs_up_5[22]));
 BUFx2_ASAP7_75t_R output3984 (.A(net3984),
    .Y(io_outs_up_5[23]));
 BUFx2_ASAP7_75t_R output3985 (.A(net3985),
    .Y(io_outs_up_5[24]));
 BUFx2_ASAP7_75t_R output3986 (.A(net3986),
    .Y(io_outs_up_5[25]));
 BUFx2_ASAP7_75t_R output3987 (.A(net3987),
    .Y(io_outs_up_5[26]));
 BUFx2_ASAP7_75t_R output3988 (.A(net3988),
    .Y(io_outs_up_5[27]));
 BUFx2_ASAP7_75t_R output3989 (.A(net3989),
    .Y(io_outs_up_5[28]));
 BUFx2_ASAP7_75t_R output3990 (.A(net3990),
    .Y(io_outs_up_5[29]));
 BUFx2_ASAP7_75t_R output3991 (.A(net3991),
    .Y(io_outs_up_5[2]));
 BUFx2_ASAP7_75t_R output3992 (.A(net3992),
    .Y(io_outs_up_5[30]));
 BUFx2_ASAP7_75t_R output3993 (.A(net3993),
    .Y(io_outs_up_5[31]));
 BUFx2_ASAP7_75t_R output3994 (.A(net3994),
    .Y(io_outs_up_5[32]));
 BUFx2_ASAP7_75t_R output3995 (.A(net3995),
    .Y(io_outs_up_5[33]));
 BUFx2_ASAP7_75t_R output3996 (.A(net3996),
    .Y(io_outs_up_5[34]));
 BUFx2_ASAP7_75t_R output3997 (.A(net3997),
    .Y(io_outs_up_5[35]));
 BUFx2_ASAP7_75t_R output3998 (.A(net3998),
    .Y(io_outs_up_5[36]));
 BUFx2_ASAP7_75t_R output3999 (.A(net3999),
    .Y(io_outs_up_5[37]));
 BUFx2_ASAP7_75t_R output4000 (.A(net4000),
    .Y(io_outs_up_5[38]));
 BUFx2_ASAP7_75t_R output4001 (.A(net4001),
    .Y(io_outs_up_5[39]));
 BUFx2_ASAP7_75t_R output4002 (.A(net4002),
    .Y(io_outs_up_5[3]));
 BUFx2_ASAP7_75t_R output4003 (.A(net4003),
    .Y(io_outs_up_5[40]));
 BUFx2_ASAP7_75t_R output4004 (.A(net4004),
    .Y(io_outs_up_5[41]));
 BUFx2_ASAP7_75t_R output4005 (.A(net4005),
    .Y(io_outs_up_5[42]));
 BUFx2_ASAP7_75t_R output4006 (.A(net4006),
    .Y(io_outs_up_5[43]));
 BUFx2_ASAP7_75t_R output4007 (.A(net4007),
    .Y(io_outs_up_5[44]));
 BUFx2_ASAP7_75t_R output4008 (.A(net4008),
    .Y(io_outs_up_5[45]));
 BUFx2_ASAP7_75t_R output4009 (.A(net4009),
    .Y(io_outs_up_5[46]));
 BUFx2_ASAP7_75t_R output4010 (.A(net4010),
    .Y(io_outs_up_5[47]));
 BUFx2_ASAP7_75t_R output4011 (.A(net4011),
    .Y(io_outs_up_5[48]));
 BUFx2_ASAP7_75t_R output4012 (.A(net4012),
    .Y(io_outs_up_5[49]));
 BUFx2_ASAP7_75t_R output4013 (.A(net4013),
    .Y(io_outs_up_5[4]));
 BUFx2_ASAP7_75t_R output4014 (.A(net4014),
    .Y(io_outs_up_5[50]));
 BUFx2_ASAP7_75t_R output4015 (.A(net4015),
    .Y(io_outs_up_5[51]));
 BUFx2_ASAP7_75t_R output4016 (.A(net4016),
    .Y(io_outs_up_5[52]));
 BUFx2_ASAP7_75t_R output4017 (.A(net4017),
    .Y(io_outs_up_5[53]));
 BUFx2_ASAP7_75t_R output4018 (.A(net4018),
    .Y(io_outs_up_5[54]));
 BUFx2_ASAP7_75t_R output4019 (.A(net4019),
    .Y(io_outs_up_5[55]));
 BUFx2_ASAP7_75t_R output4020 (.A(net4020),
    .Y(io_outs_up_5[56]));
 BUFx2_ASAP7_75t_R output4021 (.A(net4021),
    .Y(io_outs_up_5[57]));
 BUFx2_ASAP7_75t_R output4022 (.A(net4022),
    .Y(io_outs_up_5[58]));
 BUFx2_ASAP7_75t_R output4023 (.A(net4023),
    .Y(io_outs_up_5[59]));
 BUFx2_ASAP7_75t_R output4024 (.A(net4024),
    .Y(io_outs_up_5[5]));
 BUFx2_ASAP7_75t_R output4025 (.A(net4025),
    .Y(io_outs_up_5[60]));
 BUFx2_ASAP7_75t_R output4026 (.A(net4026),
    .Y(io_outs_up_5[61]));
 BUFx2_ASAP7_75t_R output4027 (.A(net4027),
    .Y(io_outs_up_5[62]));
 BUFx2_ASAP7_75t_R output4028 (.A(net4028),
    .Y(io_outs_up_5[63]));
 BUFx2_ASAP7_75t_R output4029 (.A(net4029),
    .Y(io_outs_up_5[6]));
 BUFx2_ASAP7_75t_R output4030 (.A(net4030),
    .Y(io_outs_up_5[7]));
 BUFx2_ASAP7_75t_R output4031 (.A(net4031),
    .Y(io_outs_up_5[8]));
 BUFx2_ASAP7_75t_R output4032 (.A(net4032),
    .Y(io_outs_up_5[9]));
 BUFx2_ASAP7_75t_R output4033 (.A(net4033),
    .Y(io_outs_up_6[0]));
 BUFx2_ASAP7_75t_R output4034 (.A(net4034),
    .Y(io_outs_up_6[10]));
 BUFx2_ASAP7_75t_R output4035 (.A(net4035),
    .Y(io_outs_up_6[11]));
 BUFx2_ASAP7_75t_R output4036 (.A(net4036),
    .Y(io_outs_up_6[12]));
 BUFx2_ASAP7_75t_R output4037 (.A(net4037),
    .Y(io_outs_up_6[13]));
 BUFx2_ASAP7_75t_R output4038 (.A(net4038),
    .Y(io_outs_up_6[14]));
 BUFx2_ASAP7_75t_R output4039 (.A(net4039),
    .Y(io_outs_up_6[15]));
 BUFx2_ASAP7_75t_R output4040 (.A(net4040),
    .Y(io_outs_up_6[16]));
 BUFx2_ASAP7_75t_R output4041 (.A(net4041),
    .Y(io_outs_up_6[17]));
 BUFx2_ASAP7_75t_R output4042 (.A(net4042),
    .Y(io_outs_up_6[18]));
 BUFx2_ASAP7_75t_R output4043 (.A(net4043),
    .Y(io_outs_up_6[19]));
 BUFx2_ASAP7_75t_R output4044 (.A(net4044),
    .Y(io_outs_up_6[1]));
 BUFx2_ASAP7_75t_R output4045 (.A(net4045),
    .Y(io_outs_up_6[20]));
 BUFx2_ASAP7_75t_R output4046 (.A(net4046),
    .Y(io_outs_up_6[21]));
 BUFx2_ASAP7_75t_R output4047 (.A(net4047),
    .Y(io_outs_up_6[22]));
 BUFx2_ASAP7_75t_R output4048 (.A(net4048),
    .Y(io_outs_up_6[23]));
 BUFx2_ASAP7_75t_R output4049 (.A(net4049),
    .Y(io_outs_up_6[24]));
 BUFx2_ASAP7_75t_R output4050 (.A(net4050),
    .Y(io_outs_up_6[25]));
 BUFx2_ASAP7_75t_R output4051 (.A(net4051),
    .Y(io_outs_up_6[26]));
 BUFx2_ASAP7_75t_R output4052 (.A(net4052),
    .Y(io_outs_up_6[27]));
 BUFx2_ASAP7_75t_R output4053 (.A(net4053),
    .Y(io_outs_up_6[28]));
 BUFx2_ASAP7_75t_R output4054 (.A(net4054),
    .Y(io_outs_up_6[29]));
 BUFx2_ASAP7_75t_R output4055 (.A(net4055),
    .Y(io_outs_up_6[2]));
 BUFx2_ASAP7_75t_R output4056 (.A(net4056),
    .Y(io_outs_up_6[30]));
 BUFx2_ASAP7_75t_R output4057 (.A(net4057),
    .Y(io_outs_up_6[31]));
 BUFx2_ASAP7_75t_R output4058 (.A(net4058),
    .Y(io_outs_up_6[32]));
 BUFx2_ASAP7_75t_R output4059 (.A(net4059),
    .Y(io_outs_up_6[33]));
 BUFx2_ASAP7_75t_R output4060 (.A(net4060),
    .Y(io_outs_up_6[34]));
 BUFx2_ASAP7_75t_R output4061 (.A(net4061),
    .Y(io_outs_up_6[35]));
 BUFx2_ASAP7_75t_R output4062 (.A(net4062),
    .Y(io_outs_up_6[36]));
 BUFx2_ASAP7_75t_R output4063 (.A(net4063),
    .Y(io_outs_up_6[37]));
 BUFx2_ASAP7_75t_R output4064 (.A(net4064),
    .Y(io_outs_up_6[38]));
 BUFx2_ASAP7_75t_R output4065 (.A(net4065),
    .Y(io_outs_up_6[39]));
 BUFx2_ASAP7_75t_R output4066 (.A(net4066),
    .Y(io_outs_up_6[3]));
 BUFx2_ASAP7_75t_R output4067 (.A(net4067),
    .Y(io_outs_up_6[40]));
 BUFx2_ASAP7_75t_R output4068 (.A(net4068),
    .Y(io_outs_up_6[41]));
 BUFx2_ASAP7_75t_R output4069 (.A(net4069),
    .Y(io_outs_up_6[42]));
 BUFx2_ASAP7_75t_R output4070 (.A(net4070),
    .Y(io_outs_up_6[43]));
 BUFx2_ASAP7_75t_R output4071 (.A(net4071),
    .Y(io_outs_up_6[44]));
 BUFx2_ASAP7_75t_R output4072 (.A(net4072),
    .Y(io_outs_up_6[45]));
 BUFx2_ASAP7_75t_R output4073 (.A(net4073),
    .Y(io_outs_up_6[46]));
 BUFx2_ASAP7_75t_R output4074 (.A(net4074),
    .Y(io_outs_up_6[47]));
 BUFx2_ASAP7_75t_R output4075 (.A(net4075),
    .Y(io_outs_up_6[48]));
 BUFx2_ASAP7_75t_R output4076 (.A(net4076),
    .Y(io_outs_up_6[49]));
 BUFx2_ASAP7_75t_R output4077 (.A(net4077),
    .Y(io_outs_up_6[4]));
 BUFx2_ASAP7_75t_R output4078 (.A(net4078),
    .Y(io_outs_up_6[50]));
 BUFx2_ASAP7_75t_R output4079 (.A(net4079),
    .Y(io_outs_up_6[51]));
 BUFx2_ASAP7_75t_R output4080 (.A(net4080),
    .Y(io_outs_up_6[52]));
 BUFx2_ASAP7_75t_R output4081 (.A(net4081),
    .Y(io_outs_up_6[53]));
 BUFx2_ASAP7_75t_R output4082 (.A(net4082),
    .Y(io_outs_up_6[54]));
 BUFx2_ASAP7_75t_R output4083 (.A(net4083),
    .Y(io_outs_up_6[55]));
 BUFx2_ASAP7_75t_R output4084 (.A(net4084),
    .Y(io_outs_up_6[56]));
 BUFx2_ASAP7_75t_R output4085 (.A(net4085),
    .Y(io_outs_up_6[57]));
 BUFx2_ASAP7_75t_R output4086 (.A(net4086),
    .Y(io_outs_up_6[58]));
 BUFx2_ASAP7_75t_R output4087 (.A(net4087),
    .Y(io_outs_up_6[59]));
 BUFx2_ASAP7_75t_R output4088 (.A(net4088),
    .Y(io_outs_up_6[5]));
 BUFx2_ASAP7_75t_R output4089 (.A(net4089),
    .Y(io_outs_up_6[60]));
 BUFx2_ASAP7_75t_R output4090 (.A(net4090),
    .Y(io_outs_up_6[61]));
 BUFx2_ASAP7_75t_R output4091 (.A(net4091),
    .Y(io_outs_up_6[62]));
 BUFx2_ASAP7_75t_R output4092 (.A(net4092),
    .Y(io_outs_up_6[63]));
 BUFx2_ASAP7_75t_R output4093 (.A(net4093),
    .Y(io_outs_up_6[6]));
 BUFx2_ASAP7_75t_R output4094 (.A(net4094),
    .Y(io_outs_up_6[7]));
 BUFx2_ASAP7_75t_R output4095 (.A(net4095),
    .Y(io_outs_up_6[8]));
 BUFx2_ASAP7_75t_R output4096 (.A(net4096),
    .Y(io_outs_up_6[9]));
 BUFx2_ASAP7_75t_R output4097 (.A(net4097),
    .Y(io_outs_up_7[0]));
 BUFx2_ASAP7_75t_R output4098 (.A(net4098),
    .Y(io_outs_up_7[10]));
 BUFx2_ASAP7_75t_R output4099 (.A(net4099),
    .Y(io_outs_up_7[11]));
 BUFx2_ASAP7_75t_R output4100 (.A(net4100),
    .Y(io_outs_up_7[12]));
 BUFx2_ASAP7_75t_R output4101 (.A(net4101),
    .Y(io_outs_up_7[13]));
 BUFx2_ASAP7_75t_R output4102 (.A(net4102),
    .Y(io_outs_up_7[14]));
 BUFx2_ASAP7_75t_R output4103 (.A(net4103),
    .Y(io_outs_up_7[15]));
 BUFx2_ASAP7_75t_R output4104 (.A(net4104),
    .Y(io_outs_up_7[16]));
 BUFx2_ASAP7_75t_R output4105 (.A(net4105),
    .Y(io_outs_up_7[17]));
 BUFx2_ASAP7_75t_R output4106 (.A(net4106),
    .Y(io_outs_up_7[18]));
 BUFx2_ASAP7_75t_R output4107 (.A(net4107),
    .Y(io_outs_up_7[19]));
 BUFx2_ASAP7_75t_R output4108 (.A(net4108),
    .Y(io_outs_up_7[1]));
 BUFx2_ASAP7_75t_R output4109 (.A(net4109),
    .Y(io_outs_up_7[20]));
 BUFx2_ASAP7_75t_R output4110 (.A(net4110),
    .Y(io_outs_up_7[21]));
 BUFx2_ASAP7_75t_R output4111 (.A(net4111),
    .Y(io_outs_up_7[22]));
 BUFx2_ASAP7_75t_R output4112 (.A(net4112),
    .Y(io_outs_up_7[23]));
 BUFx2_ASAP7_75t_R output4113 (.A(net4113),
    .Y(io_outs_up_7[24]));
 BUFx2_ASAP7_75t_R output4114 (.A(net4114),
    .Y(io_outs_up_7[25]));
 BUFx2_ASAP7_75t_R output4115 (.A(net4115),
    .Y(io_outs_up_7[26]));
 BUFx2_ASAP7_75t_R output4116 (.A(net4116),
    .Y(io_outs_up_7[27]));
 BUFx2_ASAP7_75t_R output4117 (.A(net4117),
    .Y(io_outs_up_7[28]));
 BUFx2_ASAP7_75t_R output4118 (.A(net4118),
    .Y(io_outs_up_7[29]));
 BUFx2_ASAP7_75t_R output4119 (.A(net4119),
    .Y(io_outs_up_7[2]));
 BUFx2_ASAP7_75t_R output4120 (.A(net4120),
    .Y(io_outs_up_7[30]));
 BUFx2_ASAP7_75t_R output4121 (.A(net4121),
    .Y(io_outs_up_7[31]));
 BUFx2_ASAP7_75t_R output4122 (.A(net4122),
    .Y(io_outs_up_7[32]));
 BUFx2_ASAP7_75t_R output4123 (.A(net4123),
    .Y(io_outs_up_7[33]));
 BUFx2_ASAP7_75t_R output4124 (.A(net4124),
    .Y(io_outs_up_7[34]));
 BUFx2_ASAP7_75t_R output4125 (.A(net4125),
    .Y(io_outs_up_7[35]));
 BUFx2_ASAP7_75t_R output4126 (.A(net4126),
    .Y(io_outs_up_7[36]));
 BUFx2_ASAP7_75t_R output4127 (.A(net4127),
    .Y(io_outs_up_7[37]));
 BUFx2_ASAP7_75t_R output4128 (.A(net4128),
    .Y(io_outs_up_7[38]));
 BUFx2_ASAP7_75t_R output4129 (.A(net4129),
    .Y(io_outs_up_7[39]));
 BUFx2_ASAP7_75t_R output4130 (.A(net4130),
    .Y(io_outs_up_7[3]));
 BUFx2_ASAP7_75t_R output4131 (.A(net4131),
    .Y(io_outs_up_7[40]));
 BUFx2_ASAP7_75t_R output4132 (.A(net4132),
    .Y(io_outs_up_7[41]));
 BUFx2_ASAP7_75t_R output4133 (.A(net4133),
    .Y(io_outs_up_7[42]));
 BUFx2_ASAP7_75t_R output4134 (.A(net4134),
    .Y(io_outs_up_7[43]));
 BUFx2_ASAP7_75t_R output4135 (.A(net4135),
    .Y(io_outs_up_7[44]));
 BUFx2_ASAP7_75t_R output4136 (.A(net4136),
    .Y(io_outs_up_7[45]));
 BUFx2_ASAP7_75t_R output4137 (.A(net4137),
    .Y(io_outs_up_7[46]));
 BUFx2_ASAP7_75t_R output4138 (.A(net4138),
    .Y(io_outs_up_7[47]));
 BUFx2_ASAP7_75t_R output4139 (.A(net4139),
    .Y(io_outs_up_7[48]));
 BUFx2_ASAP7_75t_R output4140 (.A(net4140),
    .Y(io_outs_up_7[49]));
 BUFx2_ASAP7_75t_R output4141 (.A(net4141),
    .Y(io_outs_up_7[4]));
 BUFx2_ASAP7_75t_R output4142 (.A(net4142),
    .Y(io_outs_up_7[50]));
 BUFx2_ASAP7_75t_R output4143 (.A(net4143),
    .Y(io_outs_up_7[51]));
 BUFx2_ASAP7_75t_R output4144 (.A(net4144),
    .Y(io_outs_up_7[52]));
 BUFx2_ASAP7_75t_R output4145 (.A(net4145),
    .Y(io_outs_up_7[53]));
 BUFx2_ASAP7_75t_R output4146 (.A(net4146),
    .Y(io_outs_up_7[54]));
 BUFx2_ASAP7_75t_R output4147 (.A(net4147),
    .Y(io_outs_up_7[55]));
 BUFx2_ASAP7_75t_R output4148 (.A(net4148),
    .Y(io_outs_up_7[56]));
 BUFx2_ASAP7_75t_R output4149 (.A(net4149),
    .Y(io_outs_up_7[57]));
 BUFx2_ASAP7_75t_R output4150 (.A(net4150),
    .Y(io_outs_up_7[58]));
 BUFx2_ASAP7_75t_R output4151 (.A(net4151),
    .Y(io_outs_up_7[59]));
 BUFx2_ASAP7_75t_R output4152 (.A(net4152),
    .Y(io_outs_up_7[5]));
 BUFx2_ASAP7_75t_R output4153 (.A(net4153),
    .Y(io_outs_up_7[60]));
 BUFx2_ASAP7_75t_R output4154 (.A(net4154),
    .Y(io_outs_up_7[61]));
 BUFx2_ASAP7_75t_R output4155 (.A(net4155),
    .Y(io_outs_up_7[62]));
 BUFx2_ASAP7_75t_R output4156 (.A(net4156),
    .Y(io_outs_up_7[63]));
 BUFx2_ASAP7_75t_R output4157 (.A(net4157),
    .Y(io_outs_up_7[6]));
 BUFx2_ASAP7_75t_R output4158 (.A(net4158),
    .Y(io_outs_up_7[7]));
 BUFx2_ASAP7_75t_R output4159 (.A(net4159),
    .Y(io_outs_up_7[8]));
 BUFx2_ASAP7_75t_R output4160 (.A(net4160),
    .Y(io_outs_up_7[9]));
 TIELOx1_ASAP7_75t_R ces_0_0_4161 (.L(net4161));
 TIELOx1_ASAP7_75t_R ces_0_0_4162 (.L(net4162));
 TIELOx1_ASAP7_75t_R ces_0_0_4163 (.L(net4163));
 TIELOx1_ASAP7_75t_R ces_0_0_4164 (.L(net4164));
 TIELOx1_ASAP7_75t_R ces_0_0_4165 (.L(net4165));
 TIELOx1_ASAP7_75t_R ces_0_0_4166 (.L(net4166));
 TIELOx1_ASAP7_75t_R ces_0_0_4167 (.L(net4167));
 TIELOx1_ASAP7_75t_R ces_1_0_4168 (.L(net4168));
 TIELOx1_ASAP7_75t_R ces_1_0_4169 (.L(net4169));
 TIELOx1_ASAP7_75t_R ces_1_0_4170 (.L(net4170));
 TIELOx1_ASAP7_75t_R ces_1_0_4171 (.L(net4171));
 TIELOx1_ASAP7_75t_R ces_1_0_4172 (.L(net4172));
 TIELOx1_ASAP7_75t_R ces_1_0_4173 (.L(net4173));
 TIELOx1_ASAP7_75t_R ces_1_0_4174 (.L(net4174));
 TIELOx1_ASAP7_75t_R ces_2_0_4175 (.L(net4175));
 TIELOx1_ASAP7_75t_R ces_2_0_4176 (.L(net4176));
 TIELOx1_ASAP7_75t_R ces_2_0_4177 (.L(net4177));
 TIELOx1_ASAP7_75t_R ces_2_0_4178 (.L(net4178));
 TIELOx1_ASAP7_75t_R ces_2_0_4179 (.L(net4179));
 TIELOx1_ASAP7_75t_R ces_2_0_4180 (.L(net4180));
 TIELOx1_ASAP7_75t_R ces_2_0_4181 (.L(net4181));
 TIELOx1_ASAP7_75t_R ces_3_0_4182 (.L(net4182));
 TIELOx1_ASAP7_75t_R ces_3_0_4183 (.L(net4183));
 TIELOx1_ASAP7_75t_R ces_3_0_4184 (.L(net4184));
 TIELOx1_ASAP7_75t_R ces_3_0_4185 (.L(net4185));
 TIELOx1_ASAP7_75t_R ces_3_0_4186 (.L(net4186));
 TIELOx1_ASAP7_75t_R ces_3_0_4187 (.L(net4187));
 TIELOx1_ASAP7_75t_R ces_3_0_4188 (.L(net4188));
 TIELOx1_ASAP7_75t_R ces_4_0_4189 (.L(net4189));
 TIELOx1_ASAP7_75t_R ces_4_0_4190 (.L(net4190));
 TIELOx1_ASAP7_75t_R ces_4_0_4191 (.L(net4191));
 TIELOx1_ASAP7_75t_R ces_4_0_4192 (.L(net4192));
 TIELOx1_ASAP7_75t_R ces_4_0_4193 (.L(net4193));
 TIELOx1_ASAP7_75t_R ces_4_0_4194 (.L(net4194));
 TIELOx1_ASAP7_75t_R ces_4_0_4195 (.L(net4195));
 TIELOx1_ASAP7_75t_R ces_5_0_4196 (.L(net4196));
 TIELOx1_ASAP7_75t_R ces_5_0_4197 (.L(net4197));
 TIELOx1_ASAP7_75t_R ces_5_0_4198 (.L(net4198));
 TIELOx1_ASAP7_75t_R ces_5_0_4199 (.L(net4199));
 TIELOx1_ASAP7_75t_R ces_5_0_4200 (.L(net4200));
 TIELOx1_ASAP7_75t_R ces_5_0_4201 (.L(net4201));
 TIELOx1_ASAP7_75t_R ces_5_0_4202 (.L(net4202));
 TIELOx1_ASAP7_75t_R ces_6_0_4203 (.L(net4203));
 TIELOx1_ASAP7_75t_R ces_6_0_4204 (.L(net4204));
 TIELOx1_ASAP7_75t_R ces_6_0_4205 (.L(net4205));
 TIELOx1_ASAP7_75t_R ces_6_0_4206 (.L(net4206));
 TIELOx1_ASAP7_75t_R ces_6_0_4207 (.L(net4207));
 TIELOx1_ASAP7_75t_R ces_6_0_4208 (.L(net4208));
 TIELOx1_ASAP7_75t_R ces_6_0_4209 (.L(net4209));
 TIELOx1_ASAP7_75t_R ces_7_0_4210 (.L(net4210));
 TIELOx1_ASAP7_75t_R ces_7_0_4211 (.L(net4211));
 TIELOx1_ASAP7_75t_R ces_7_0_4212 (.L(net4212));
 TIELOx1_ASAP7_75t_R ces_7_0_4213 (.L(net4213));
 TIELOx1_ASAP7_75t_R ces_7_0_4214 (.L(net4214));
 TIELOx1_ASAP7_75t_R ces_7_0_4215 (.L(net4215));
 TIELOx1_ASAP7_75t_R ces_7_0_4216 (.L(net4216));
 BUFx24_ASAP7_75t_R clkbuf_0_clock (.A(net4217),
    .Y(clknet_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_1_0_0_clock (.A(clknet_0_clock),
    .Y(clknet_1_0_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_1_1_0_clock (.A(clknet_0_clock),
    .Y(clknet_1_1_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_2_0_0_clock (.A(clknet_1_0_0_clock),
    .Y(clknet_2_0_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_2_1_0_clock (.A(clknet_1_0_0_clock),
    .Y(clknet_2_1_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_2_2_0_clock (.A(clknet_1_1_0_clock),
    .Y(clknet_2_2_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_2_3_0_clock (.A(clknet_1_1_0_clock),
    .Y(clknet_2_3_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_3_0_0_clock (.A(clknet_2_0_0_clock),
    .Y(clknet_3_0_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_3_1_0_clock (.A(clknet_2_0_0_clock),
    .Y(clknet_3_1_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_3_2_0_clock (.A(clknet_2_1_0_clock),
    .Y(clknet_3_2_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_3_3_0_clock (.A(clknet_2_1_0_clock),
    .Y(clknet_3_3_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_3_4_0_clock (.A(clknet_2_2_0_clock),
    .Y(clknet_3_4_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_3_5_0_clock (.A(clknet_2_2_0_clock),
    .Y(clknet_3_5_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_3_6_0_clock (.A(clknet_2_3_0_clock),
    .Y(clknet_3_6_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_3_7_0_clock (.A(clknet_2_3_0_clock),
    .Y(clknet_3_7_0_clock));
 BUFx24_ASAP7_75t_R clkbuf_0_clock_regs (.A(clock_regs),
    .Y(clknet_0_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_3_0_0_clock_regs (.A(clknet_0_clock_regs),
    .Y(clknet_3_0_0_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_3_1_0_clock_regs (.A(clknet_0_clock_regs),
    .Y(clknet_3_1_0_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_3_2_0_clock_regs (.A(clknet_0_clock_regs),
    .Y(clknet_3_2_0_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_3_3_0_clock_regs (.A(clknet_0_clock_regs),
    .Y(clknet_3_3_0_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_3_4_0_clock_regs (.A(clknet_0_clock_regs),
    .Y(clknet_3_4_0_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_3_5_0_clock_regs (.A(clknet_0_clock_regs),
    .Y(clknet_3_5_0_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_3_6_0_clock_regs (.A(clknet_0_clock_regs),
    .Y(clknet_3_6_0_clock_regs));
 BUFx24_ASAP7_75t_R clkbuf_3_7_0_clock_regs (.A(clknet_0_clock_regs),
    .Y(clknet_3_7_0_clock_regs));
 INVxp67_ASAP7_75t_R clkload0 (.A(clknet_3_1_0_clock_regs));
 BUFx4f_ASAP7_75t_R clkload1 (.A(clknet_3_2_0_clock_regs));
 INVxp67_ASAP7_75t_R clkload2 (.A(clknet_3_3_0_clock_regs));
 BUFx4f_ASAP7_75t_R clkload3 (.A(clknet_3_4_0_clock_regs));
 BUFx4f_ASAP7_75t_R clkload4 (.A(clknet_3_7_0_clock_regs));
 BUFx24_ASAP7_75t_R delaybuf_0_clock (.A(delaynet_0_clock),
    .Y(delaynet_1_clock));
 BUFx24_ASAP7_75t_R delaybuf_1_clock (.A(delaynet_1_clock),
    .Y(delaynet_2_clock));
 BUFx24_ASAP7_75t_R delaybuf_2_clock (.A(delaynet_2_clock),
    .Y(delaynet_3_clock));
 BUFx24_ASAP7_75t_R delaybuf_3_clock (.A(delaynet_3_clock),
    .Y(delaynet_4_clock));
 BUFx24_ASAP7_75t_R delaybuf_4_clock (.A(delaynet_4_clock),
    .Y(delaynet_5_clock));
 BUFx24_ASAP7_75t_R delaybuf_5_clock (.A(delaynet_5_clock),
    .Y(clock_regs));
 BUFx16f_ASAP7_75t_R wire1 (.A(net4218),
    .Y(net4217));
 BUFx6f_ASAP7_75t_R wire2 (.A(clock),
    .Y(net4218));
 DECAPx10_ASAP7_75t_R FILLER_0_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_332 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_354 ();
 FILLER_ASAP7_75t_R FILLER_0_0_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_382 ();
 FILLER_ASAP7_75t_R FILLER_0_0_393 ();
 FILLER_ASAP7_75t_R FILLER_0_0_405 ();
 FILLER_ASAP7_75t_R FILLER_0_0_412 ();
 FILLER_ASAP7_75t_R FILLER_0_0_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_421 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_461 ();
 FILLER_ASAP7_75t_R FILLER_0_0_464 ();
 FILLER_ASAP7_75t_R FILLER_0_0_476 ();
 FILLER_ASAP7_75t_R FILLER_0_0_488 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_495 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_566 ();
 FILLER_ASAP7_75t_R FILLER_0_0_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_580 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1124 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1201 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1212 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1224 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_1236 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1240 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_1246 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1250 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1271 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_1282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1288 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1294 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_1306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1367 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1380 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1393 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1818 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_1840 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1846 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_1938 ();
 FILLER_ASAP7_75t_R FILLER_0_0_1960 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_1962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2198 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2220 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2242 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2264 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2286 ();
 FILLER_ASAP7_75t_R FILLER_0_0_2308 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2730 ();
 DECAPx4_ASAP7_75t_R FILLER_0_0_2752 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_2767 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_2771 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_2774 ();
 FILLER_ASAP7_75t_R FILLER_0_0_2893 ();
 FILLER_ASAP7_75t_R FILLER_0_0_2910 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_2912 ();
 FILLER_ASAP7_75t_R FILLER_0_0_2978 ();
 FILLER_ASAP7_75t_R FILLER_0_0_2985 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_2987 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_2998 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3020 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3042 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3064 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3086 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3108 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3130 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3174 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3196 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_3218 ();
 FILLER_ASAP7_75t_R FILLER_0_0_3232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3522 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_3544 ();
 FILLER_ASAP7_75t_R FILLER_0_0_3558 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_3560 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_3571 ();
 FILLER_ASAP7_75t_R FILLER_0_0_3577 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_3589 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_3605 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_3624 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_3663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_3679 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_3695 ();
 FILLER_ASAP7_75t_R FILLER_0_0_3763 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3800 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3822 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3844 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3866 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3888 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3910 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3932 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3954 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3976 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_3998 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4020 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4042 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4064 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4086 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4108 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4130 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4336 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_4358 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_4397 ();
 FILLER_ASAP7_75t_R FILLER_0_0_4428 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_4495 ();
 FILLER_ASAP7_75t_R FILLER_0_0_4544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_4546 ();
 FILLER_ASAP7_75t_R FILLER_0_0_4567 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_4569 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_4580 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_4601 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_4615 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_4619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5128 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_5150 ();
 FILLER_ASAP7_75t_R FILLER_0_0_5164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_5196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_5207 ();
 FILLER_ASAP7_75t_R FILLER_0_0_5218 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_5250 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_5254 ();
 FILLER_ASAP7_75t_R FILLER_0_0_5280 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_5287 ();
 DECAPx2_ASAP7_75t_R FILLER_0_0_5308 ();
 DECAPx4_ASAP7_75t_R FILLER_0_0_5324 ();
 FILLER_ASAP7_75t_R FILLER_0_0_5384 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_5386 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5397 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5419 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5441 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5463 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5485 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5507 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_5529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_5543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_5942 ();
 FILLER_ASAP7_75t_R FILLER_0_0_5964 ();
 FILLER_ASAP7_75t_R FILLER_0_0_6193 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6442 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_6464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_332 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_368 ();
 FILLER_ASAP7_75t_R FILLER_0_1_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_411 ();
 FILLER_ASAP7_75t_R FILLER_0_1_417 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_458 ();
 FILLER_ASAP7_75t_R FILLER_0_1_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_476 ();
 FILLER_ASAP7_75t_R FILLER_0_1_487 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_541 ();
 FILLER_ASAP7_75t_R FILLER_0_1_547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_558 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_594 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_638 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_704 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_726 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_748 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_770 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_792 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_814 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_836 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_858 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_880 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_902 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1124 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_1146 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1176 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_1183 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1189 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1191 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_1207 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1216 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1222 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1237 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1243 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1245 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1251 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1258 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_1264 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1309 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1315 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1327 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1333 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_1348 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1352 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1363 ();
 FILLER_ASAP7_75t_R FILLER_0_1_1369 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1387 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1393 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1415 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1437 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1459 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1481 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1503 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1525 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1569 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1591 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1613 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1635 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1657 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1679 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1701 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1723 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1745 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1767 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1789 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1811 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_1833 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1847 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_1938 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1_1960 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1970 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_1981 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_1985 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_2001 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2005 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2016 ();
 FILLER_ASAP7_75t_R FILLER_0_1_2022 ();
 FILLER_ASAP7_75t_R FILLER_0_1_2034 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_2056 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2060 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2066 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2072 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2078 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_2084 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_2093 ();
 FILLER_ASAP7_75t_R FILLER_0_1_2099 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_2116 ();
 FILLER_ASAP7_75t_R FILLER_0_1_2125 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2127 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2133 ();
 FILLER_ASAP7_75t_R FILLER_0_1_2139 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_2156 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2191 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2197 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2219 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2241 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2263 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2285 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2307 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2329 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2351 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2373 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2395 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2417 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2439 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2483 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2505 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2527 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2549 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2571 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2593 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2615 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2637 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2659 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2681 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2703 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2725 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1_2747 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_2762 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2766 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2794 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2800 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_2841 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2845 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1_2896 ();
 FILLER_ASAP7_75t_R FILLER_0_1_2926 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_2933 ();
 FILLER_ASAP7_75t_R FILLER_0_1_2939 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_2946 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2957 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_2963 ();
 FILLER_ASAP7_75t_R FILLER_0_1_2969 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3524 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_3546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_3560 ();
 FILLER_ASAP7_75t_R FILLER_0_1_3626 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_3653 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_3664 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_3680 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_3686 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_3692 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_3713 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_3719 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_3725 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_3729 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_3740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_3744 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_3750 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_3769 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_3775 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_3781 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_3785 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_3994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4324 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_4346 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_4360 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_4371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4375 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_4406 ();
 FILLER_ASAP7_75t_R FILLER_0_1_4412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4414 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_4425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4431 ();
 FILLER_ASAP7_75t_R FILLER_0_1_4437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4439 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4445 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_4451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4455 ();
 FILLER_ASAP7_75t_R FILLER_0_1_4466 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_4478 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_4492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4502 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_4518 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_4549 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_4558 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4564 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_4570 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4576 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_4582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4591 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_4613 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_4619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5128 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_5150 ();
 FILLER_ASAP7_75t_R FILLER_0_1_5164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5191 ();
 FILLER_ASAP7_75t_R FILLER_0_1_5202 ();
 FILLER_ASAP7_75t_R FILLER_0_1_5214 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_5221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5246 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_5252 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5258 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5269 ();
 FILLER_ASAP7_75t_R FILLER_0_1_5290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5303 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_5379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5383 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5389 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5411 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5433 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5455 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5477 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5499 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5521 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_5920 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_5942 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_5956 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5962 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_5968 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1_5999 ();
 FILLER_ASAP7_75t_R FILLER_0_1_6009 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_6011 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_6022 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_6026 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1_6037 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_6047 ();
 FILLER_ASAP7_75t_R FILLER_0_1_6058 ();
 FILLER_ASAP7_75t_R FILLER_0_1_6065 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_6077 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_6081 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_6092 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_6096 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_6107 ();
 FILLER_ASAP7_75t_R FILLER_0_1_6116 ();
 FILLER_ASAP7_75t_R FILLER_0_1_6128 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_6135 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_6151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_6157 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_6163 ();
 FILLER_ASAP7_75t_R FILLER_0_1_6182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6436 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1_6458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_332 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_354 ();
 FILLER_ASAP7_75t_R FILLER_0_2_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_373 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_379 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_393 ();
 FILLER_ASAP7_75t_R FILLER_0_2_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_411 ();
 FILLER_ASAP7_75t_R FILLER_0_2_417 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_429 ();
 FILLER_ASAP7_75t_R FILLER_0_2_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_445 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_451 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_479 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_490 ();
 FILLER_ASAP7_75t_R FILLER_0_2_496 ();
 FILLER_ASAP7_75t_R FILLER_0_2_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_510 ();
 FILLER_ASAP7_75t_R FILLER_0_2_516 ();
 FILLER_ASAP7_75t_R FILLER_0_2_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_525 ();
 FILLER_ASAP7_75t_R FILLER_0_2_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_533 ();
 FILLER_ASAP7_75t_R FILLER_0_2_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_541 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_551 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_562 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_604 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_626 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_648 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_670 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_692 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_714 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_736 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_758 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_780 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_802 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_824 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_846 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_868 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_890 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_912 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_934 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_956 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_978 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1022 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1044 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1066 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1088 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1132 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_1154 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1164 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_1170 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1178 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_1199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1219 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_1226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1232 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_1258 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_1269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1273 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1287 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1293 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_1304 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_1313 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1323 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1325 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1336 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1344 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1350 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_1356 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1385 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_1938 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1960 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1962 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_1968 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1974 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_1993 ();
 FILLER_ASAP7_75t_R FILLER_0_2_1999 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2001 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2007 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_2014 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2018 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2029 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_2035 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2041 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_2062 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2072 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2084 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2108 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2114 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_2126 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2132 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2139 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2145 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_2152 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_2163 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2173 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2179 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2201 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2245 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2267 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_2289 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_2303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2309 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2730 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_2752 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2779 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2801 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2803 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_2809 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2823 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2825 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2831 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2833 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_2839 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2853 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2855 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_2861 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2871 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2873 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2884 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_2890 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2909 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2916 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2918 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2924 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2931 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_2942 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_2951 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2957 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2964 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_2970 ();
 FILLER_ASAP7_75t_R FILLER_0_2_2976 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2978 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_2984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2990 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3012 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3034 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3056 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3078 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3122 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3144 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3166 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3188 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3210 ();
 FILLER_ASAP7_75t_R FILLER_0_2_3232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3544 ();
 FILLER_ASAP7_75t_R FILLER_0_2_3566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_3568 ();
 FILLER_ASAP7_75t_R FILLER_0_2_3574 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_3586 ();
 FILLER_ASAP7_75t_R FILLER_0_2_3592 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_3599 ();
 FILLER_ASAP7_75t_R FILLER_0_2_3620 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_3622 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_3638 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_3657 ();
 FILLER_ASAP7_75t_R FILLER_0_2_3663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_3665 ();
 FILLER_ASAP7_75t_R FILLER_0_2_3681 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_3693 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_3722 ();
 FILLER_ASAP7_75t_R FILLER_0_2_3728 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_3730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_3736 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_3752 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_3768 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3792 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3814 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3836 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3858 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3880 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3902 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3924 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3946 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3968 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_3990 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4012 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4034 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4056 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4078 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4122 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_4144 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4336 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_4358 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4368 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_4374 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_4388 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4398 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_4404 ();
 FILLER_ASAP7_75t_R FILLER_0_2_4418 ();
 FILLER_ASAP7_75t_R FILLER_0_2_4425 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_4437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4441 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4452 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_4458 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4464 ();
 FILLER_ASAP7_75t_R FILLER_0_2_4470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4472 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_4478 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_4489 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4493 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_4504 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4515 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_4526 ();
 FILLER_ASAP7_75t_R FILLER_0_2_4532 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4539 ();
 FILLER_ASAP7_75t_R FILLER_0_2_4545 ();
 FILLER_ASAP7_75t_R FILLER_0_2_4552 ();
 FILLER_ASAP7_75t_R FILLER_0_2_4559 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4561 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_4572 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_4576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4604 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4626 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4648 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4670 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4692 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4714 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4736 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4758 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4780 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4802 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4824 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4846 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4868 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4890 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4912 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4934 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4956 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_4978 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5022 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5044 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_5066 ();
 FILLER_ASAP7_75t_R FILLER_0_2_5080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5150 ();
 FILLER_ASAP7_75t_R FILLER_0_2_5182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_5189 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_5195 ();
 FILLER_ASAP7_75t_R FILLER_0_2_5210 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_5222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_5241 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_5252 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_5263 ();
 FILLER_ASAP7_75t_R FILLER_0_2_5269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_5271 ();
 FILLER_ASAP7_75t_R FILLER_0_2_5277 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_5284 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_5293 ();
 FILLER_ASAP7_75t_R FILLER_0_2_5303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_5305 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_5311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_5315 ();
 FILLER_ASAP7_75t_R FILLER_0_2_5326 ();
 FILLER_ASAP7_75t_R FILLER_0_2_5333 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_5335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_5351 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_5357 ();
 FILLER_ASAP7_75t_R FILLER_0_2_5367 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_5379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_5393 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5399 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5421 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5443 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5465 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5487 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5509 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5531 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5553 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5575 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5597 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5641 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5663 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5685 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5707 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5729 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5751 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5773 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5795 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5817 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5839 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5861 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5883 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5905 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_5927 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_5949 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_5963 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_5974 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_5980 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_5986 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_5990 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_6013 ();
 DECAPx6_ASAP7_75t_R FILLER_0_2_6034 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_6048 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_6054 ();
 FILLER_ASAP7_75t_R FILLER_0_2_6065 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_6067 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_6078 ();
 FILLER_ASAP7_75t_R FILLER_0_2_6084 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_6086 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_6097 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_6103 ();
 FILLER_ASAP7_75t_R FILLER_0_2_6113 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_6115 ();
 FILLER_ASAP7_75t_R FILLER_0_2_6121 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_6128 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_6134 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_6150 ();
 FILLER_ASAP7_75t_R FILLER_0_2_6156 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_6168 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_6183 ();
 FILLER_ASAP7_75t_R FILLER_0_2_6189 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6201 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6245 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6267 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6289 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6311 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6333 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6355 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6377 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6399 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6421 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6443 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6465 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6487 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6509 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_6531 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_332 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_354 ();
 FILLER_ASAP7_75t_R FILLER_0_3_368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_375 ();
 FILLER_ASAP7_75t_R FILLER_0_3_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_389 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_411 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_454 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_460 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_475 ();
 FILLER_ASAP7_75t_R FILLER_0_3_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_494 ();
 FILLER_ASAP7_75t_R FILLER_0_3_505 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_516 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_522 ();
 FILLER_ASAP7_75t_R FILLER_0_3_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_544 ();
 FILLER_ASAP7_75t_R FILLER_0_3_555 ();
 FILLER_ASAP7_75t_R FILLER_0_3_567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1175 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_1191 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1216 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1235 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_1241 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1249 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1260 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1275 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_1296 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1310 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1323 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_1329 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1335 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_1342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_1351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_1360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1816 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_1838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_1938 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_1960 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_1984 ();
 FILLER_ASAP7_75t_R FILLER_0_3_1994 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2001 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_2007 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_2016 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2020 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_2026 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2032 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_2039 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_2053 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2059 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2065 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_2071 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_2090 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2096 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_2102 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2112 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2114 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_2120 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_2136 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2150 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2174 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2218 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2240 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2284 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2350 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2372 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2394 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2416 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2438 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2482 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2504 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2526 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2548 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2570 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2592 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2636 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2658 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2680 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2702 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2724 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2746 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_2768 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2774 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2781 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_2807 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2813 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2815 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_2826 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2840 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2856 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2863 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2870 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_2892 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2906 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_2918 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2928 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2930 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2936 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2943 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2945 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_2961 ();
 FILLER_ASAP7_75t_R FILLER_0_3_2967 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_2969 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2975 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2997 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3019 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3041 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3063 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3085 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3107 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3129 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3151 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3173 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3283 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3327 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3349 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3371 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3393 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3415 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3437 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3459 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3481 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3503 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3525 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3569 ();
 FILLER_ASAP7_75t_R FILLER_0_3_3591 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_3598 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_3604 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_3618 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_3624 ();
 FILLER_ASAP7_75t_R FILLER_0_3_3634 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_3641 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_3647 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_3653 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_3659 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_3673 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_3679 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_3690 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_3698 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_3704 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_3710 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_3721 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_3730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_3741 ();
 FILLER_ASAP7_75t_R FILLER_0_3_3747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_3749 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_3755 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_3769 ();
 FILLER_ASAP7_75t_R FILLER_0_3_3785 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3792 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3814 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3836 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3858 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3880 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3902 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3924 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3946 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3968 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_3990 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4012 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4034 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4056 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4078 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4122 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4144 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4166 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4188 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4210 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4298 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4342 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4364 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_4386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_4392 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_4408 ();
 FILLER_ASAP7_75t_R FILLER_0_3_4418 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_4430 ();
 FILLER_ASAP7_75t_R FILLER_0_3_4436 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_4443 ();
 FILLER_ASAP7_75t_R FILLER_0_3_4449 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_4451 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_4457 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_4468 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_4474 ();
 FILLER_ASAP7_75t_R FILLER_0_3_4485 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_4487 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_4503 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_4512 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_4523 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_4537 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_4558 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_4569 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_4583 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4594 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_4616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5150 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_5172 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_5186 ();
 FILLER_ASAP7_75t_R FILLER_0_3_5197 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_5209 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_5223 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_5229 ();
 FILLER_ASAP7_75t_R FILLER_0_3_5235 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_5237 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_5248 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_5257 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_5268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_5272 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_5278 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_5284 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_5290 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_5304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_5308 ();
 FILLER_ASAP7_75t_R FILLER_0_3_5314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_5316 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_5327 ();
 FILLER_ASAP7_75t_R FILLER_0_3_5333 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_5335 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_5341 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_5355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_5364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_5370 ();
 FILLER_ASAP7_75t_R FILLER_0_3_5376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5520 ();
 FILLER_ASAP7_75t_R FILLER_0_3_5542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_5964 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_5986 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_5992 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_5998 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6009 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_6031 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_6037 ();
 FILLER_ASAP7_75t_R FILLER_0_3_6053 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_6060 ();
 FILLER_ASAP7_75t_R FILLER_0_3_6066 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_6078 ();
 FILLER_ASAP7_75t_R FILLER_0_3_6084 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_6086 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_6092 ();
 FILLER_ASAP7_75t_R FILLER_0_3_6108 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_6115 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_6126 ();
 FILLER_ASAP7_75t_R FILLER_0_3_6136 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_6143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_6152 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_6156 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_6167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_6171 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_6177 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6188 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6210 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6298 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6342 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6364 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6386 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6430 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_6452 ();
 FILLER_ASAP7_75t_R FILLER_0_3_6466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_9_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_13_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_51 ();
 FILLER_ASAP7_75t_R FILLER_0_72_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_72_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_6529 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_73_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_73_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_6552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_2 ();
 FILLER_ASAP7_75t_R FILLER_0_74_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_6523 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_6537 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_75_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_6532 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_6543 ();
 FILLER_ASAP7_75t_R FILLER_0_75_6549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_2 ();
 FILLER_ASAP7_75t_R FILLER_0_76_8 ();
 FILLER_ASAP7_75t_R FILLER_0_76_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_76_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_77_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_77_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_6542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_2 ();
 FILLER_ASAP7_75t_R FILLER_0_78_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_51 ();
 FILLER_ASAP7_75t_R FILLER_0_78_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_78_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_6522 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_6533 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_6557 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_79_13 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_59 ();
 FILLER_ASAP7_75t_R FILLER_0_79_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_79_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_81_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_81_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_81_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_6537 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_83_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_6547 ();
 FILLER_ASAP7_75t_R FILLER_0_84_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_4 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_14 ();
 FILLER_ASAP7_75t_R FILLER_0_84_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_84_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_84_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_85_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_32 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_60 ();
 FILLER_ASAP7_75t_R FILLER_0_86_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_86_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_6528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_6537 ();
 DECAPx1_ASAP7_75t_R FILLER_0_86_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_86_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_44 ();
 FILLER_ASAP7_75t_R FILLER_0_87_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_87_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_87_6524 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_6540 ();
 DECAPx4_ASAP7_75t_R FILLER_0_87_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_87_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_44 ();
 FILLER_ASAP7_75t_R FILLER_0_88_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_88_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_6547 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_56 ();
 FILLER_ASAP7_75t_R FILLER_0_90_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_90_6551 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_12 ();
 FILLER_ASAP7_75t_R FILLER_0_91_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_91_52 ();
 FILLER_ASAP7_75t_R FILLER_0_91_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_6548 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_6547 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_2 ();
 FILLER_ASAP7_75t_R FILLER_0_93_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_93_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_18 ();
 FILLER_ASAP7_75t_R FILLER_0_94_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_8 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_95_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_6522 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_6539 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_17 ();
 FILLER_ASAP7_75t_R FILLER_0_96_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_96_6523 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_6525 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_6531 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_51 ();
 FILLER_ASAP7_75t_R FILLER_0_97_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_6537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_97_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_6 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_98_6546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_13 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_99_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_99_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_6547 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_12 ();
 FILLER_ASAP7_75t_R FILLER_0_100_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_51 ();
 FILLER_ASAP7_75t_R FILLER_0_100_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_43 ();
 FILLER_ASAP7_75t_R FILLER_0_101_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_101_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_101_6542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_6544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_101_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_11 ();
 FILLER_ASAP7_75t_R FILLER_0_102_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_102_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_6529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_6535 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_103_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_14 ();
 FILLER_ASAP7_75t_R FILLER_0_103_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_103_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_103_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_103_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_6530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_103_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_103_6551 ();
 DECAPx4_ASAP7_75t_R FILLER_0_104_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_44 ();
 FILLER_ASAP7_75t_R FILLER_0_104_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_104_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_6 ();
 DECAPx6_ASAP7_75t_R FILLER_0_105_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_105_59 ();
 FILLER_ASAP7_75t_R FILLER_0_105_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_105_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_6537 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_13 ();
 FILLER_ASAP7_75t_R FILLER_0_106_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_106_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_106_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_106_6538 ();
 DECAPx4_ASAP7_75t_R FILLER_0_107_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_107_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_107_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_107_6528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_6535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_6539 ();
 DECAPx4_ASAP7_75t_R FILLER_0_107_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_107_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_108_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_108_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_108_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_6535 ();
 FILLER_ASAP7_75t_R FILLER_0_108_6545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_6547 ();
 FILLER_ASAP7_75t_R FILLER_0_109_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_4 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_109_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_6529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_6533 ();
 DECAPx6_ASAP7_75t_R FILLER_0_109_6539 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_110_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_110_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_111_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_111_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_111_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_112_2 ();
 FILLER_ASAP7_75t_R FILLER_0_112_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_112_51 ();
 FILLER_ASAP7_75t_R FILLER_0_112_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_112_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_112_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_6530 ();
 FILLER_ASAP7_75t_R FILLER_0_112_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_6538 ();
 DECAPx6_ASAP7_75t_R FILLER_0_112_6544 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_44 ();
 FILLER_ASAP7_75t_R FILLER_0_113_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_113_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_2 ();
 FILLER_ASAP7_75t_R FILLER_0_114_8 ();
 FILLER_ASAP7_75t_R FILLER_0_114_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_114_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_114_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_114_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_6530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_114_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_114_6551 ();
 DECAPx6_ASAP7_75t_R FILLER_0_115_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_115_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_115_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_115_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_6546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_116_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_116_6556 ();
 DECAPx6_ASAP7_75t_R FILLER_0_117_7 ();
 FILLER_ASAP7_75t_R FILLER_0_117_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_33 ();
 DECAPx4_ASAP7_75t_R FILLER_0_117_55 ();
 FILLER_ASAP7_75t_R FILLER_0_117_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_117_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_117_6540 ();
 DECAPx4_ASAP7_75t_R FILLER_0_117_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_118_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_34 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_56 ();
 FILLER_ASAP7_75t_R FILLER_0_118_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_118_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_6530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_119_46 ();
 FILLER_ASAP7_75t_R FILLER_0_119_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_24 ();
 DECAPx4_ASAP7_75t_R FILLER_0_120_46 ();
 FILLER_ASAP7_75t_R FILLER_0_120_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_58 ();
 FILLER_ASAP7_75t_R FILLER_0_120_62 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_121_46 ();
 FILLER_ASAP7_75t_R FILLER_0_121_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_152_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_152_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_152_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_152_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_152_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_152_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_153_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_154_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_155_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_157_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_158_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_158_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_158_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_158_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_158_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_158_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_159_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_159_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_159_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_159_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_159_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_159_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_160_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_160_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_160_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_160_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_160_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_160_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_161_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_162_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_163_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_164_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_165_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_166_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_167_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_168_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_169_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_170_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_171_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_172_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_173_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_174_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_175_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_176_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_177_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_178_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_178_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_179_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_179_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_179_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_180_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_180_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_180_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_181_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_181_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_181_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_182_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_182_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_182_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_183_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_183_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_183_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_184_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_184_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_184_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_185_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_185_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_185_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_186_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_186_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_186_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_187_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_187_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_187_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_188_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_188_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_188_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_189_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_189_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_189_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_190_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_191_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_192_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_193_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_194_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_195_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_196_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_197_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_198_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_199_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_201_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_202_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_203_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_204_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_205_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_206_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_207_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_208_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_209_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_210_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_211_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_212_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_213_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_214_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_215_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_216_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_217_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_218_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_219_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_220_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_221_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_223_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_224_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_225_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_225_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_225_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_225_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_225_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_225_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_226_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_227_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_228_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_229_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_230_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_231_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_231_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_231_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_231_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_231_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_231_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_232_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_232_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_232_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_232_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_232_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_232_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_233_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_234_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_235_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_235_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_235_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_235_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_235_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_235_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_236_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_236_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_236_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_236_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_236_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_236_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_237_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_238_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_239_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_240_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_240_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_240_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_240_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_240_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_240_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_241_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_242_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_243_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_244_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_245_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_246_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_247_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_247_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_247_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_247_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_247_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_247_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_248_2 ();
 FILLER_ASAP7_75t_R FILLER_0_248_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_248_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_248_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_248_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_248_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_248_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_248_6522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_248_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_248_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_248_6556 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_2 ();
 FILLER_ASAP7_75t_R FILLER_0_249_8 ();
 DECAPx2_ASAP7_75t_R FILLER_0_249_15 ();
 FILLER_ASAP7_75t_R FILLER_0_249_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_249_56 ();
 FILLER_ASAP7_75t_R FILLER_0_249_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_249_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_249_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_6538 ();
 FILLER_ASAP7_75t_R FILLER_0_249_6549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_249_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_2 ();
 FILLER_ASAP7_75t_R FILLER_0_250_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_250_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_250_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_250_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_250_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_250_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_251_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_251_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_251_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_251_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_251_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_252_12 ();
 FILLER_ASAP7_75t_R FILLER_0_252_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_252_56 ();
 FILLER_ASAP7_75t_R FILLER_0_252_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_252_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_252_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_6537 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_252_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_252_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_253_7 ();
 FILLER_ASAP7_75t_R FILLER_0_253_17 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_253_56 ();
 FILLER_ASAP7_75t_R FILLER_0_253_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_253_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_253_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_253_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_253_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_12 ();
 FILLER_ASAP7_75t_R FILLER_0_254_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_254_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_254_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_254_6536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_254_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_255_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_255_12 ();
 FILLER_ASAP7_75t_R FILLER_0_255_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_24 ();
 DECAPx1_ASAP7_75t_R FILLER_0_255_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_34 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_255_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_255_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_255_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_255_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_255_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_255_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_256_2 ();
 FILLER_ASAP7_75t_R FILLER_0_256_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_256_51 ();
 FILLER_ASAP7_75t_R FILLER_0_256_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_256_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_256_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_256_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_6532 ();
 DECAPx6_ASAP7_75t_R FILLER_0_256_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_256_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_257_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_257_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_257_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_257_6522 ();
 DECAPx4_ASAP7_75t_R FILLER_0_257_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_257_6543 ();
 DECAPx1_ASAP7_75t_R FILLER_0_257_6554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_258_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_43 ();
 FILLER_ASAP7_75t_R FILLER_0_258_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_258_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_258_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_258_6522 ();
 DECAPx6_ASAP7_75t_R FILLER_0_258_6533 ();
 DECAPx2_ASAP7_75t_R FILLER_0_258_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_259_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_259_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_259_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_259_6551 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_260_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_260_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_260_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_260_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_260_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_6540 ();
 DECAPx2_ASAP7_75t_R FILLER_0_260_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_260_6552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_261_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_261_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_261_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_261_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_261_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_261_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_261_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_262_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_262_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_262_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_262_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_262_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_262_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_262_6531 ();
 FILLER_ASAP7_75t_R FILLER_0_262_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_262_6548 ();
 FILLER_ASAP7_75t_R FILLER_0_262_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_262_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_59 ();
 FILLER_ASAP7_75t_R FILLER_0_263_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_263_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_263_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_263_6522 ();
 DECAPx6_ASAP7_75t_R FILLER_0_263_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_263_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_44 ();
 FILLER_ASAP7_75t_R FILLER_0_264_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_264_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_264_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_264_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_264_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_265_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_265_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_265_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_6539 ();
 FILLER_ASAP7_75t_R FILLER_0_265_6545 ();
 DECAPx2_ASAP7_75t_R FILLER_0_265_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_266_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_44 ();
 FILLER_ASAP7_75t_R FILLER_0_266_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_266_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_266_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_266_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_266_6535 ();
 DECAPx1_ASAP7_75t_R FILLER_0_266_6549 ();
 DECAPx1_ASAP7_75t_R FILLER_0_267_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_12 ();
 FILLER_ASAP7_75t_R FILLER_0_267_18 ();
 FILLER_ASAP7_75t_R FILLER_0_267_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_267_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_267_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_267_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_267_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_267_6544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_267_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_267_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_268_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_44 ();
 FILLER_ASAP7_75t_R FILLER_0_268_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_268_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_268_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_268_6524 ();
 DECAPx6_ASAP7_75t_R FILLER_0_268_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_268_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_268_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_44 ();
 FILLER_ASAP7_75t_R FILLER_0_269_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_269_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_269_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_269_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_6522 ();
 DECAPx6_ASAP7_75t_R FILLER_0_269_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_269_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_269_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_270_2 ();
 FILLER_ASAP7_75t_R FILLER_0_270_9 ();
 DECAPx4_ASAP7_75t_R FILLER_0_270_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_270_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_270_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_270_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_270_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_270_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_2 ();
 FILLER_ASAP7_75t_R FILLER_0_271_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_10 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_271_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_271_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_271_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_271_6544 ();
 FILLER_ASAP7_75t_R FILLER_0_271_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_271_6552 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_8 ();
 FILLER_ASAP7_75t_R FILLER_0_272_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_44 ();
 FILLER_ASAP7_75t_R FILLER_0_272_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_272_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_272_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_272_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_272_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_273_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_9 ();
 DECAPx6_ASAP7_75t_R FILLER_0_273_15 ();
 FILLER_ASAP7_75t_R FILLER_0_273_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_273_59 ();
 FILLER_ASAP7_75t_R FILLER_0_273_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_273_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_273_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_273_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_273_6534 ();
 DECAPx2_ASAP7_75t_R FILLER_0_273_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_273_6556 ();
 FILLER_ASAP7_75t_R FILLER_0_274_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_14 ();
 FILLER_ASAP7_75t_R FILLER_0_274_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_274_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_274_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_274_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_274_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_274_6522 ();
 DECAPx6_ASAP7_75t_R FILLER_0_274_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_274_6542 ();
 DECAPx6_ASAP7_75t_R FILLER_0_275_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_16 ();
 FILLER_ASAP7_75t_R FILLER_0_275_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_275_56 ();
 FILLER_ASAP7_75t_R FILLER_0_275_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_275_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_275_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_275_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_275_6534 ();
 DECAPx1_ASAP7_75t_R FILLER_0_276_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_276_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_276_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_276_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_276_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_276_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_276_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_276_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_276_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_276_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_276_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_276_6530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_276_6541 ();
 DECAPx4_ASAP7_75t_R FILLER_0_276_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_276_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_277_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_277_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_277_44 ();
 FILLER_ASAP7_75t_R FILLER_0_277_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_277_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_277_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_277_6529 ();
 FILLER_ASAP7_75t_R FILLER_0_277_6535 ();
 DECAPx6_ASAP7_75t_R FILLER_0_277_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_277_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_278_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_278_6 ();
 FILLER_ASAP7_75t_R FILLER_0_278_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_278_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_278_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_278_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_278_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_278_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_278_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_278_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_278_6538 ();
 DECAPx1_ASAP7_75t_R FILLER_0_278_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_278_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_279_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_279_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_279_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_279_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_279_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_279_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_279_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_279_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_279_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_279_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_279_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_279_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_279_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_280_7 ();
 FILLER_ASAP7_75t_R FILLER_0_280_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_280_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_280_51 ();
 FILLER_ASAP7_75t_R FILLER_0_280_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_280_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_280_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_280_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_280_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_280_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_280_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_280_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_280_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_281_2 ();
 FILLER_ASAP7_75t_R FILLER_0_281_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_281_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_281_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_281_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_281_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_281_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_281_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_281_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_281_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_281_6541 ();
 DECAPx1_ASAP7_75t_R FILLER_0_281_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_281_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_282_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_282_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_282_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_282_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_282_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_282_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_282_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_282_6530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_282_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_282_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_283_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_283_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_283_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_283_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_283_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_283_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_283_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_283_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_283_6522 ();
 DECAPx4_ASAP7_75t_R FILLER_0_283_6528 ();
 FILLER_ASAP7_75t_R FILLER_0_283_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_283_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_283_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_283_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_283_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_284_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_284_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_284_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_284_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_284_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_284_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_284_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_284_6534 ();
 DECAPx1_ASAP7_75t_R FILLER_0_284_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_284_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_285_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_285_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_285_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_285_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_285_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_285_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_285_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_285_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_285_6522 ();
 DECAPx4_ASAP7_75t_R FILLER_0_285_6528 ();
 FILLER_ASAP7_75t_R FILLER_0_285_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_285_6540 ();
 DECAPx4_ASAP7_75t_R FILLER_0_285_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_285_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_286_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_286_11 ();
 DECAPx1_ASAP7_75t_R FILLER_0_286_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_286_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_286_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_286_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_286_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_286_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_286_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_286_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_286_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_286_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_286_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_287_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_287_9 ();
 DECAPx2_ASAP7_75t_R FILLER_0_287_15 ();
 FILLER_ASAP7_75t_R FILLER_0_287_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_287_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_287_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_287_51 ();
 FILLER_ASAP7_75t_R FILLER_0_287_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_287_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_287_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_287_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_287_6518 ();
 DECAPx6_ASAP7_75t_R FILLER_0_287_6524 ();
 DECAPx1_ASAP7_75t_R FILLER_0_287_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_287_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_287_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_287_6552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_288_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_288_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_288_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_288_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_288_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_288_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_288_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_288_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_288_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_288_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_288_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_289_2 ();
 FILLER_ASAP7_75t_R FILLER_0_289_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_289_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_289_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_289_52 ();
 FILLER_ASAP7_75t_R FILLER_0_289_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_289_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_289_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_289_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_289_6532 ();
 DECAPx2_ASAP7_75t_R FILLER_0_289_6538 ();
 FILLER_ASAP7_75t_R FILLER_0_289_6544 ();
 FILLER_ASAP7_75t_R FILLER_0_289_6551 ();
 DECAPx4_ASAP7_75t_R FILLER_0_290_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_290_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_290_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_290_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_290_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_290_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_290_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_290_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_290_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_290_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_290_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_290_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_290_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_291_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_291_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_291_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_291_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_291_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_291_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_291_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_291_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_291_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_291_6532 ();
 DECAPx6_ASAP7_75t_R FILLER_0_291_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_291_6557 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_292_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_292_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_292_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_292_41 ();
 DECAPx1_ASAP7_75t_R FILLER_0_292_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_292_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_292_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_292_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_292_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_292_6530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_292_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_292_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_292_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_293_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_293_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_293_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_293_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_293_51 ();
 FILLER_ASAP7_75t_R FILLER_0_293_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_293_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_293_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_293_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_293_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_293_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_294_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_294_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_294_39 ();
 DECAPx1_ASAP7_75t_R FILLER_0_294_61 ();
 DECAPx10_ASAP7_75t_R FILLER_0_294_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_294_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_294_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_294_6530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_294_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_295_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_295_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_295_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_295_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_295_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_295_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_295_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_295_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_296_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_296_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_296_46 ();
 FILLER_ASAP7_75t_R FILLER_0_296_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_296_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_296_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_296_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_297_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_297_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_297_46 ();
 FILLER_ASAP7_75t_R FILLER_0_297_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_297_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_297_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_297_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_298_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_298_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_298_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_298_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_298_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_298_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_299_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_299_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_299_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_299_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_299_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_299_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_300_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_300_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_300_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_300_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_300_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_300_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_301_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_301_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_301_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_301_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_301_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_301_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_302_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_302_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_302_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_302_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_302_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_302_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_303_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_303_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_303_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_303_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_303_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_303_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_304_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_304_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_304_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_304_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_304_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_304_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_305_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_305_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_305_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_305_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_305_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_305_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_306_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_306_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_306_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_306_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_306_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_306_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_307_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_307_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_307_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_307_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_307_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_307_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_308_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_308_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_308_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_308_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_308_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_308_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_309_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_309_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_309_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_309_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_309_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_309_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_310_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_310_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_310_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_310_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_310_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_310_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_311_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_311_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_311_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_311_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_311_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_311_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_312_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_312_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_312_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_312_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_312_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_312_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_313_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_313_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_313_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_313_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_313_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_313_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_314_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_314_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_314_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_314_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_314_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_314_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_315_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_315_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_315_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_315_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_315_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_315_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_316_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_316_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_316_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_316_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_316_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_316_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_317_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_317_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_317_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_317_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_317_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_317_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_318_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_318_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_318_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_318_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_318_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_318_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_319_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_319_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_319_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_319_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_319_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_319_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_320_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_320_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_320_46 ();
 FILLER_ASAP7_75t_R FILLER_0_320_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_320_6515 ();
 DECAPx6_ASAP7_75t_R FILLER_0_320_6537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_320_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_320_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_321_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_321_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_321_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_321_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_321_6506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_321_6510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_321_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_321_6554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_322_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_322_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_322_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_322_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_322_6506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_322_6508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_322_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_322_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_323_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_323_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_323_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_323_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_323_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_323_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_324_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_324_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_324_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_324_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_324_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_324_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_325_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_325_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_325_46 ();
 FILLER_ASAP7_75t_R FILLER_0_325_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_325_6515 ();
 DECAPx6_ASAP7_75t_R FILLER_0_325_6537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_325_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_325_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_326_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_326_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_326_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_326_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_326_6502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_326_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_326_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_326_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_327_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_327_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_327_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_327_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_327_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_328_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_328_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_328_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_328_6513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_328_6535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_328_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_329_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_329_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_329_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_329_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_329_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_329_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_330_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_330_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_330_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_330_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_330_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_330_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_331_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_331_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_331_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_331_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_331_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_331_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_332_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_332_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_332_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_332_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_332_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_332_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_333_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_333_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_333_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_333_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_333_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_333_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_334_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_334_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_334_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_334_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_334_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_334_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_335_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_335_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_335_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_335_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_335_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_335_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_336_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_336_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_336_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_336_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_336_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_336_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_337_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_337_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_337_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_337_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_337_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_337_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_338_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_338_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_338_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_338_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_338_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_338_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_339_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_339_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_339_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_339_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_339_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_339_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_340_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_340_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_340_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_340_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_340_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_340_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_341_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_341_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_341_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_341_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_341_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_341_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_342_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_342_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_342_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_342_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_342_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_342_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_343_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_343_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_343_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_343_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_343_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_343_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_344_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_344_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_344_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_344_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_344_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_344_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_345_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_345_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_345_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_345_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_345_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_345_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_346_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_346_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_346_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_346_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_346_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_346_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_347_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_347_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_347_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_347_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_347_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_347_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_348_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_348_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_348_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_348_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_348_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_348_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_349_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_349_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_349_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_349_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_349_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_349_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_350_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_350_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_350_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_350_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_350_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_350_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_351_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_351_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_351_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_351_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_351_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_351_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_352_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_352_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_352_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_352_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_352_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_352_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_353_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_353_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_353_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_353_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_353_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_353_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_354_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_354_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_354_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_355_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_355_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_355_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_355_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_355_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_355_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_355_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_355_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_355_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_355_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_355_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_355_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_355_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_355_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_355_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_356_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_356_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_356_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_356_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_356_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_356_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_356_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_356_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_356_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_356_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_356_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_356_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_356_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_356_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_356_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_357_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_357_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_357_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_357_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_357_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_357_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_357_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_357_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_357_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_357_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_357_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_357_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_357_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_357_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_357_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_358_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_358_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_358_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_358_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_358_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_358_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_358_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_358_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_358_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_358_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_358_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_358_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_358_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_358_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_358_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_359_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_359_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_359_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_359_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_359_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_359_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_359_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_359_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_359_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_359_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_359_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_359_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_359_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_359_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_359_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_360_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_360_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_360_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_360_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_360_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_360_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_360_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_360_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_360_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_360_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_360_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_360_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_360_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_360_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_360_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_361_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_361_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_361_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_361_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_361_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_361_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_361_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_361_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_361_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_361_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_361_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_361_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_361_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_361_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_361_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_362_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_362_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_362_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_362_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_362_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_362_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_362_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_362_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_362_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_362_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_362_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_362_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_362_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_362_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_362_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_363_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_363_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_363_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_363_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_363_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_363_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_363_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_363_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_363_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_363_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_363_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_363_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_363_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_363_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_363_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_364_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_364_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_364_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_364_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_364_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_364_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_364_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_364_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_364_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_364_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_364_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_364_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_364_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_364_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_364_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1674 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_1696 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_1710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1746 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1768 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1790 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1812 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_1834 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_4982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5048 ();
 DECAPx4_ASAP7_75t_R FILLER_0_365_5070 ();
 FILLER_ASAP7_75t_R FILLER_0_365_5080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_365_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_365_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_365_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_366_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_366_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_366_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_366_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_366_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_366_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_367_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_367_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_367_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_367_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_367_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_367_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_368_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_368_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_368_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_368_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_368_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_368_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_369_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_369_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_369_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_369_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_369_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_369_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_370_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_370_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_370_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_370_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_370_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_370_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_371_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_371_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_371_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_371_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_371_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_371_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_372_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_372_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_372_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_372_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_372_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_372_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_373_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_373_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_373_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_373_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_373_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_373_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_374_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_374_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_374_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_374_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_374_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_374_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_375_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_375_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_375_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_375_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_375_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_375_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_376_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_376_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_376_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_376_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_376_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_376_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_377_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_377_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_377_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_377_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_377_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_377_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_378_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_378_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_378_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_378_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_378_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_378_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_379_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_379_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_379_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_379_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_379_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_379_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_380_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_380_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_380_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_380_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_380_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_380_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_381_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_381_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_381_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_381_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_381_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_381_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_382_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_382_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_382_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_382_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_382_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_382_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_383_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_383_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_383_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_383_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_383_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_383_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_384_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_384_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_384_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_384_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_384_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_384_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_385_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_385_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_385_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_385_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_385_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_385_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_386_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_386_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_386_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_386_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_386_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_386_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_387_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_387_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_387_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_387_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_387_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_387_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_388_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_388_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_388_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_388_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_388_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_388_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_389_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_389_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_389_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_389_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_389_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_389_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_390_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_390_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_390_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_390_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_390_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_390_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_391_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_391_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_391_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_391_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_391_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_391_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_392_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_392_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_392_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_392_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_392_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_392_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_393_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_393_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_393_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_393_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_393_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_393_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_394_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_394_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_394_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_394_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_394_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_394_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_395_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_395_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_395_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_395_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_395_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_395_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_396_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_396_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_396_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_396_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_396_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_396_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_397_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_397_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_397_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_397_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_397_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_397_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_398_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_398_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_398_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_398_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_398_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_398_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_399_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_399_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_399_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_399_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_399_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_399_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_400_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_400_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_400_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_400_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_400_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_400_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_401_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_401_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_401_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_401_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_401_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_401_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_402_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_402_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_402_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_402_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_402_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_402_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_403_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_403_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_403_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_403_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_403_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_403_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_404_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_404_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_404_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_404_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_404_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_404_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_405_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_405_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_405_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_405_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_405_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_405_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_406_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_406_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_406_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_406_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_406_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_406_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_407_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_407_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_407_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_407_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_407_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_407_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_408_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_408_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_408_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_408_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_408_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_408_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_409_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_409_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_409_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_409_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_409_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_409_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_410_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_410_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_410_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_410_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_410_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_410_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_411_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_411_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_411_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_411_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_411_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_411_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_412_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_412_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_412_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_412_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_412_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_412_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_413_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_413_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_413_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_413_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_413_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_413_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_414_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_414_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_414_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_414_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_414_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_414_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_415_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_415_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_415_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_415_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_415_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_415_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_416_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_416_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_416_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_416_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_416_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_416_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_417_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_417_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_417_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_417_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_417_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_417_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_418_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_418_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_418_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_418_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_418_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_418_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_419_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_419_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_419_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_419_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_419_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_419_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_420_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_420_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_420_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_420_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_420_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_420_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_421_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_421_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_421_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_421_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_421_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_421_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_422_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_422_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_422_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_422_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_422_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_422_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_423_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_423_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_423_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_423_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_423_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_423_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_424_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_424_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_424_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_424_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_424_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_424_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_424_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_424_6528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_424_6535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_424_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_425_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_425_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_425_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_425_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_425_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_425_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_425_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_425_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_425_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_425_6539 ();
 FILLER_ASAP7_75t_R FILLER_0_425_6545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_425_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_425_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_425_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_426_7 ();
 DECAPx1_ASAP7_75t_R FILLER_0_426_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_426_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_426_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_426_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_426_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_426_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_426_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_426_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_426_6530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_426_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_426_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_426_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_427_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_427_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_427_13 ();
 FILLER_ASAP7_75t_R FILLER_0_427_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_427_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_427_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_427_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_427_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_427_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_427_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_427_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_427_6536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_427_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_427_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_427_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_427_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_428_12 ();
 FILLER_ASAP7_75t_R FILLER_0_428_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_428_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_428_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_428_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_428_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_428_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_428_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_428_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_428_6537 ();
 DECAPx1_ASAP7_75t_R FILLER_0_428_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_428_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_429_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_429_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_429_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_429_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_429_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_429_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_429_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_429_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_429_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_429_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_429_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_429_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_430_2 ();
 FILLER_ASAP7_75t_R FILLER_0_430_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_430_10 ();
 DECAPx10_ASAP7_75t_R FILLER_0_430_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_430_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_430_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_430_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_430_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_430_6533 ();
 FILLER_ASAP7_75t_R FILLER_0_430_6539 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_430_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_430_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_430_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_430_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_431_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_431_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_431_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_431_59 ();
 FILLER_ASAP7_75t_R FILLER_0_431_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_431_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_431_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_431_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_431_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_431_6534 ();
 DECAPx4_ASAP7_75t_R FILLER_0_432_2 ();
 FILLER_ASAP7_75t_R FILLER_0_432_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_432_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_432_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_432_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_432_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_432_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_432_6546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_433_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_433_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_433_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_433_67 ();
 DECAPx6_ASAP7_75t_R FILLER_0_433_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_433_6506 ();
 DECAPx1_ASAP7_75t_R FILLER_0_433_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_433_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_434_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_434_13 ();
 FILLER_ASAP7_75t_R FILLER_0_434_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_434_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_434_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_434_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_434_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_434_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_434_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_434_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_434_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_434_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_434_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_434_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_434_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_435_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_435_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_435_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_435_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_435_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_435_67 ();
 DECAPx1_ASAP7_75t_R FILLER_0_435_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_435_6517 ();
 DECAPx2_ASAP7_75t_R FILLER_0_435_6531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_435_6537 ();
 DECAPx1_ASAP7_75t_R FILLER_0_435_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_435_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_436_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_436_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_436_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_436_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_436_54 ();
 DECAPx2_ASAP7_75t_R FILLER_0_436_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_436_6519 ();
 DECAPx1_ASAP7_75t_R FILLER_0_436_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_436_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_436_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_436_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_436_6548 ();
 DECAPx4_ASAP7_75t_R FILLER_0_437_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_437_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_437_18 ();
 FILLER_ASAP7_75t_R FILLER_0_437_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_437_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_437_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_437_59 ();
 FILLER_ASAP7_75t_R FILLER_0_437_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_437_67 ();
 DECAPx6_ASAP7_75t_R FILLER_0_437_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_437_6506 ();
 DECAPx4_ASAP7_75t_R FILLER_0_437_6531 ();
 FILLER_ASAP7_75t_R FILLER_0_437_6541 ();
 DECAPx1_ASAP7_75t_R FILLER_0_437_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_437_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_438_12 ();
 FILLER_ASAP7_75t_R FILLER_0_438_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_438_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_438_51 ();
 FILLER_ASAP7_75t_R FILLER_0_438_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_438_67 ();
 DECAPx4_ASAP7_75t_R FILLER_0_438_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_438_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_438_6532 ();
 DECAPx6_ASAP7_75t_R FILLER_0_438_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_438_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_439_7 ();
 FILLER_ASAP7_75t_R FILLER_0_439_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_439_15 ();
 DECAPx6_ASAP7_75t_R FILLER_0_439_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_439_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_439_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_439_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_439_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_439_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_439_6542 ();
 DECAPx6_ASAP7_75t_R FILLER_0_440_2 ();
 FILLER_ASAP7_75t_R FILLER_0_440_16 ();
 DECAPx2_ASAP7_75t_R FILLER_0_440_23 ();
 FILLER_ASAP7_75t_R FILLER_0_440_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_440_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_440_58 ();
 FILLER_ASAP7_75t_R FILLER_0_440_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_440_6494 ();
 DECAPx1_ASAP7_75t_R FILLER_0_440_6537 ();
 FILLER_ASAP7_75t_R FILLER_0_440_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_441_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_441_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_441_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_441_44 ();
 FILLER_ASAP7_75t_R FILLER_0_441_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_441_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_441_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_441_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_441_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_441_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_441_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_441_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_441_6557 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_442_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_442_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_442_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_442_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_442_64 ();
 DECAPx4_ASAP7_75t_R FILLER_0_442_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_442_6502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_442_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_442_6544 ();
 DECAPx1_ASAP7_75t_R FILLER_0_442_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_442_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_443_7 ();
 FILLER_ASAP7_75t_R FILLER_0_443_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_443_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_443_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_443_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_443_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_443_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_443_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_443_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_443_6547 ();
 DECAPx4_ASAP7_75t_R FILLER_0_444_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_444_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_444_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_444_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_444_33 ();
 DECAPx4_ASAP7_75t_R FILLER_0_444_55 ();
 FILLER_ASAP7_75t_R FILLER_0_444_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_444_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_444_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_444_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_444_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_444_6547 ();
 FILLER_ASAP7_75t_R FILLER_0_445_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_445_9 ();
 DECAPx10_ASAP7_75t_R FILLER_0_445_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_445_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_445_59 ();
 FILLER_ASAP7_75t_R FILLER_0_445_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_445_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_445_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_445_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_445_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_445_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_446_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_446_12 ();
 FILLER_ASAP7_75t_R FILLER_0_446_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_446_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_446_52 ();
 FILLER_ASAP7_75t_R FILLER_0_446_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_446_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_446_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_446_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_446_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_446_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_447_7 ();
 DECAPx1_ASAP7_75t_R FILLER_0_447_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_447_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_447_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_447_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_447_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_447_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_447_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_447_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_447_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_447_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_447_6540 ();
 DECAPx2_ASAP7_75t_R FILLER_0_447_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_447_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_448_12 ();
 FILLER_ASAP7_75t_R FILLER_0_448_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_448_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_448_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_448_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_448_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_448_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_448_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_448_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_448_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_448_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_448_6542 ();
 DECAPx2_ASAP7_75t_R FILLER_0_448_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_448_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_448_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_449_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_449_13 ();
 FILLER_ASAP7_75t_R FILLER_0_449_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_449_21 ();
 FILLER_ASAP7_75t_R FILLER_0_449_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_449_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_449_56 ();
 FILLER_ASAP7_75t_R FILLER_0_449_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_449_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_449_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_449_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_449_6526 ();
 DECAPx2_ASAP7_75t_R FILLER_0_449_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_449_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_449_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_449_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_449_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_450_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_450_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_450_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_450_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_450_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_450_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_450_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_450_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_450_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_450_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_450_6548 ();
 DECAPx1_ASAP7_75t_R FILLER_0_450_6554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_451_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_451_11 ();
 DECAPx2_ASAP7_75t_R FILLER_0_451_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_451_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_451_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_451_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_451_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_451_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_451_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_451_6535 ();
 FILLER_ASAP7_75t_R FILLER_0_451_6545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_451_6547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_452_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_452_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_452_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_452_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_452_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_452_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_452_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_452_6542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_453_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_453_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_453_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_453_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_453_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_453_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_453_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_453_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_453_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_453_6546 ();
 DECAPx6_ASAP7_75t_R FILLER_0_454_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_454_21 ();
 FILLER_ASAP7_75t_R FILLER_0_454_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_454_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_454_56 ();
 FILLER_ASAP7_75t_R FILLER_0_454_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_454_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_454_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_454_6533 ();
 DECAPx1_ASAP7_75t_R FILLER_0_454_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_454_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_455_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_455_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_455_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_455_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_455_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_455_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_455_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_455_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_455_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_456_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_456_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_456_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_456_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_456_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_456_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_456_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_456_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_456_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_456_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_456_6522 ();
 DECAPx1_ASAP7_75t_R FILLER_0_456_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_456_6532 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_456_6538 ();
 DECAPx6_ASAP7_75t_R FILLER_0_456_6544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_457_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_457_13 ();
 FILLER_ASAP7_75t_R FILLER_0_457_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_457_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_457_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_457_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_457_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_457_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_457_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_457_6552 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_458_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_458_13 ();
 DECAPx10_ASAP7_75t_R FILLER_0_458_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_458_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_458_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_458_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_458_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_458_6530 ();
 DECAPx6_ASAP7_75t_R FILLER_0_458_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_458_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_458_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_459_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_459_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_459_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_459_44 ();
 FILLER_ASAP7_75t_R FILLER_0_459_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_459_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_459_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_459_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_459_6539 ();
 DECAPx1_ASAP7_75t_R FILLER_0_459_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_459_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_460_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_460_11 ();
 DECAPx2_ASAP7_75t_R FILLER_0_460_17 ();
 FILLER_ASAP7_75t_R FILLER_0_460_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_460_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_460_52 ();
 FILLER_ASAP7_75t_R FILLER_0_460_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_460_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_460_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_460_6528 ();
 FILLER_ASAP7_75t_R FILLER_0_460_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_460_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_460_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_461_2 ();
 FILLER_ASAP7_75t_R FILLER_0_461_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_461_10 ();
 DECAPx1_ASAP7_75t_R FILLER_0_461_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_461_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_461_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_461_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_461_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_461_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_461_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_461_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_461_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_461_6538 ();
 DECAPx6_ASAP7_75t_R FILLER_0_462_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_462_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_462_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_462_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_462_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_462_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_462_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_462_6547 ();
 DECAPx2_ASAP7_75t_R FILLER_0_463_2 ();
 FILLER_ASAP7_75t_R FILLER_0_463_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_463_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_463_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_463_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_463_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_463_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_463_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_463_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_463_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_463_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_463_6530 ();
 DECAPx6_ASAP7_75t_R FILLER_0_463_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_463_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_463_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_464_12 ();
 FILLER_ASAP7_75t_R FILLER_0_464_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_464_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_464_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_464_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_464_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_464_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_464_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_464_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_464_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_465_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_465_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_465_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_465_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_465_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_465_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_465_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_465_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_465_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_465_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_465_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_465_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_465_6548 ();
 FILLER_ASAP7_75t_R FILLER_0_465_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_465_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_466_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_466_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_466_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_466_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_466_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_466_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_466_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_466_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_466_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_466_6542 ();
 DECAPx2_ASAP7_75t_R FILLER_0_467_2 ();
 FILLER_ASAP7_75t_R FILLER_0_467_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_467_10 ();
 DECAPx10_ASAP7_75t_R FILLER_0_467_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_467_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_467_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_467_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_467_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_467_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_467_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_467_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_467_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_467_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_467_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_467_6557 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_468_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_468_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_468_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_468_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_468_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_468_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_468_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_468_6528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_468_6539 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_468_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_468_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_468_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_468_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_469_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_469_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_469_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_469_33 ();
 DECAPx4_ASAP7_75t_R FILLER_0_469_55 ();
 FILLER_ASAP7_75t_R FILLER_0_469_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_469_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_469_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_469_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_469_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_469_6534 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_469_6540 ();
 DECAPx4_ASAP7_75t_R FILLER_0_469_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_469_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_470_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_470_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_470_51 ();
 FILLER_ASAP7_75t_R FILLER_0_470_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_470_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_470_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_470_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_470_6528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_470_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_470_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_471_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_471_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_471_46 ();
 FILLER_ASAP7_75t_R FILLER_0_471_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_471_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_471_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_471_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_472_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_472_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_472_46 ();
 FILLER_ASAP7_75t_R FILLER_0_472_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_472_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_472_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_472_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_473_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_473_24 ();
 DECAPx4_ASAP7_75t_R FILLER_0_473_46 ();
 FILLER_ASAP7_75t_R FILLER_0_473_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_473_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_473_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_473_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_473_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_474_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_474_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_474_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_474_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_474_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_474_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_475_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_475_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_475_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_475_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_475_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_475_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_476_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_476_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_476_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_476_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_476_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_476_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_477_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_477_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_477_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_477_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_477_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_477_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_478_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_478_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_478_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_478_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_478_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_478_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_479_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_479_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_479_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_479_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_479_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_479_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_480_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_480_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_480_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_480_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_480_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_480_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_481_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_481_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_481_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_481_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_481_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_481_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_482_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_482_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_482_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_482_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_482_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_482_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_483_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_483_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_483_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_483_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_483_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_483_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_484_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_484_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_484_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_484_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_484_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_484_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_485_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_485_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_485_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_485_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_485_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_485_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_486_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_486_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_486_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_486_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_486_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_486_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_487_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_487_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_487_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_487_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_487_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_487_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_488_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_488_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_488_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_488_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_488_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_488_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_489_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_489_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_489_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_489_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_489_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_489_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_490_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_490_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_490_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_490_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_490_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_490_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_491_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_491_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_491_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_491_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_491_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_491_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_492_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_492_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_492_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_492_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_492_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_492_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_493_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_493_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_493_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_493_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_493_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_493_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_494_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_494_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_494_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_494_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_494_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_494_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_495_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_495_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_495_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_495_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_495_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_495_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_496_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_496_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_496_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_496_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_496_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_496_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_497_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_497_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_497_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_497_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_497_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_497_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_498_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_498_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_498_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_498_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_498_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_498_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_499_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_499_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_499_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_499_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_499_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_499_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_500_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_500_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_500_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_500_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_500_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_500_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_501_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_501_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_501_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_501_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_501_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_501_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_502_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_502_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_502_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_502_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_502_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_502_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_503_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_503_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_503_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_503_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_503_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_503_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_504_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_504_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_504_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_504_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_504_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_504_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_505_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_505_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_505_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_505_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_505_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_505_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_506_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_506_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_506_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_506_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_506_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_506_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_507_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_507_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_507_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_507_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_507_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_507_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_508_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_508_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_508_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_508_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_508_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_508_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_509_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_509_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_509_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_509_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_509_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_509_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_510_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_510_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_510_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_510_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_510_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_510_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_511_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_511_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_511_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_511_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_511_6506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_511_6510 ();
 DECAPx6_ASAP7_75t_R FILLER_0_511_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_511_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_511_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_512_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_512_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_512_46 ();
 DECAPx2_ASAP7_75t_R FILLER_0_512_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_512_6498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_512_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_512_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_513_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_513_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_513_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_513_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_513_6506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_513_6510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_513_6519 ();
 DECAPx6_ASAP7_75t_R FILLER_0_513_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_513_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_513_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_514_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_514_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_514_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_514_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_514_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_514_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_515_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_515_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_515_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_515_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_515_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_515_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_516_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_516_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_516_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_516_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_516_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_516_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_516_6530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_516_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_517_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_517_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_517_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_517_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_517_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_517_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_517_6542 ();
 DECAPx2_ASAP7_75t_R FILLER_0_517_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_517_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_517_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_518_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_518_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_518_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_518_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_518_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_518_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_519_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_519_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_519_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_519_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_519_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_519_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_519_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_520_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_520_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_520_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_520_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_520_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_520_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_521_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_521_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_521_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_521_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_521_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_521_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_521_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_521_6537 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_521_6541 ();
 DECAPx4_ASAP7_75t_R FILLER_0_521_6548 ();
 DECAPx10_ASAP7_75t_R FILLER_0_522_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_522_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_522_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_522_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_522_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_522_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_523_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_523_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_523_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_523_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_523_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_523_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_523_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_523_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_524_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_524_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_524_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_524_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_524_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_524_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_525_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_525_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_525_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_525_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_525_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_525_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_526_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_526_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_526_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_526_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_526_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_526_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_527_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_527_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_527_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_527_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_527_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_527_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_528_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_528_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_528_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_528_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_528_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_528_6530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_528_6532 ();
 DECAPx6_ASAP7_75t_R FILLER_0_528_6539 ();
 DECAPx1_ASAP7_75t_R FILLER_0_528_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_528_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_529_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_529_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_529_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_529_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_529_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_529_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_529_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_530_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_530_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_530_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1674 ();
 DECAPx1_ASAP7_75t_R FILLER_0_530_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1818 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_1840 ();
 FILLER_ASAP7_75t_R FILLER_0_530_1846 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_530_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2488 ();
 DECAPx1_ASAP7_75t_R FILLER_0_530_2510 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_530_2514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2611 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2633 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2677 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2699 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2721 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2743 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_2765 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_530_2771 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_530_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_530_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3786 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_3808 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_530_3814 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3845 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3867 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3889 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3911 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3933 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3955 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3977 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_3999 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4021 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4043 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4065 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4087 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4109 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4131 ();
 DECAPx1_ASAP7_75t_R FILLER_0_530_4153 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_530_4157 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_530_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_4614 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_4622 ();
 FILLER_ASAP7_75t_R FILLER_0_530_4628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4704 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4726 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4748 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4770 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4792 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4814 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4836 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4858 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4880 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4902 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4924 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4946 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4968 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_4990 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5012 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5034 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5056 ();
 DECAPx1_ASAP7_75t_R FILLER_0_530_5078 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_530_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_530_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_530_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6470 ();
 FILLER_ASAP7_75t_R FILLER_0_530_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_530_6494 ();
 DECAPx10_ASAP7_75t_R FILLER_0_530_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_530_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_530_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_531_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_531_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_531_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_531_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_531_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_531_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_531_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_531_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_531_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_531_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_531_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_531_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_531_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_531_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_531_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_531_6519 ();
 DECAPx6_ASAP7_75t_R FILLER_0_531_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_531_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_531_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_532_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_532_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_532_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_532_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_532_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_532_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_532_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_532_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_532_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_532_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_532_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_532_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_532_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_532_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_532_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_533_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_533_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_533_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_533_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_533_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_533_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_533_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_533_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_533_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_533_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_533_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_533_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_533_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_533_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_533_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_534_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_534_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_534_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_534_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_534_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_534_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_534_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_534_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_534_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_534_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_534_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_534_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_534_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_534_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_534_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_535_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_535_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_535_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_535_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_535_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_535_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_535_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_535_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_535_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_535_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_535_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_535_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_535_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_535_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_535_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_536_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_536_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_536_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_536_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_536_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_536_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_536_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_536_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_536_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_536_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_536_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_536_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_536_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_536_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_536_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_537_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_537_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_537_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_537_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_537_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_537_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_537_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_537_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_537_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_537_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_537_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_537_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_537_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_537_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_537_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_538_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_538_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_538_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_538_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_538_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_538_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_538_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_538_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_538_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_538_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_538_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_538_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_538_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_538_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_538_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_539_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_539_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_539_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_539_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_539_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_539_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_539_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_539_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_539_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_539_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_539_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_539_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_539_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_539_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_539_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_540_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_540_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_540_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_540_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_540_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_540_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_540_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_540_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_540_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_540_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_540_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_540_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_540_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_540_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_540_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3126 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_3148 ();
 FILLER_ASAP7_75t_R FILLER_0_541_3162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_541_3164 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3195 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_3217 ();
 FILLER_ASAP7_75t_R FILLER_0_541_3231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_541_3233 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_3690 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_3698 ();
 FILLER_ASAP7_75t_R FILLER_0_541_3712 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_541_3714 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3745 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3767 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3789 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3811 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3833 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3855 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3877 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3899 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3921 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3943 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3965 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_3987 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4009 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4031 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4053 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4075 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4097 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4119 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_4141 ();
 FILLER_ASAP7_75t_R FILLER_0_541_4155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_541_4157 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_4160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_4174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_541_4180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4211 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4233 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4255 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4277 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4299 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4321 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4343 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4365 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4387 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4409 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4431 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4453 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4475 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4497 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4519 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4541 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4563 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4585 ();
 DECAPx4_ASAP7_75t_R FILLER_0_541_4607 ();
 FILLER_ASAP7_75t_R FILLER_0_541_4617 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_541_4619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_541_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_541_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_541_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_542_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_542_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_542_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_542_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_542_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_542_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_543_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_543_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_543_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_543_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_543_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_543_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_544_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_544_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_544_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_544_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_544_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_544_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_545_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_545_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_545_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_545_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_545_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_545_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_546_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_546_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_546_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_546_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_546_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_546_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_547_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_547_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_547_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_547_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_547_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_547_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_548_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_548_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_548_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_548_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_548_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_548_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_549_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_549_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_549_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_549_6513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_549_6535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_549_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_550_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_550_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_550_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_550_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_550_6535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_550_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_551_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_551_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_551_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_551_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_551_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_551_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_552_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_552_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_552_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_552_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_552_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_552_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_553_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_553_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_553_46 ();
 FILLER_ASAP7_75t_R FILLER_0_553_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_553_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_554_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_554_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_554_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_554_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_554_6506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_554_6531 ();
 DECAPx1_ASAP7_75t_R FILLER_0_554_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_554_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_555_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_555_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_555_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_555_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_555_6506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_555_6508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_555_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_555_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_556_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_556_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_556_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_556_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_556_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_556_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_557_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_557_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_557_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_557_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_557_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_557_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_558_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_558_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_558_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_558_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_558_6506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_558_6529 ();
 DECAPx2_ASAP7_75t_R FILLER_0_558_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_558_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_559_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_559_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_559_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_559_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_559_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_559_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_560_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_560_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_560_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_560_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_560_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_560_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_561_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_561_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_561_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_561_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_561_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_561_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_562_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_562_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_562_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_562_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_562_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_562_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_563_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_563_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_563_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_563_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_563_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_563_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_564_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_564_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_564_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_564_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_564_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_564_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_565_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_565_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_565_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_565_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_565_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_565_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_566_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_566_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_566_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_566_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_566_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_566_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_567_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_567_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_567_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_567_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_567_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_567_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_568_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_568_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_568_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_568_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_568_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_568_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_569_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_569_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_569_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_569_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_569_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_569_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_570_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_570_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_570_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_570_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_570_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_570_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_571_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_571_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_571_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_571_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_571_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_571_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_572_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_572_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_572_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_572_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_572_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_572_6528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_572_6535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_572_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_573_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_573_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_573_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_573_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_573_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_573_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_574_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_574_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_574_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_574_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_574_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_574_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_575_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_575_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_575_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_575_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_575_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_575_6536 ();
 DECAPx6_ASAP7_75t_R FILLER_0_575_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_575_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_576_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_576_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_576_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_576_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_576_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_576_6524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_576_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_576_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_577_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_577_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_577_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_577_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_577_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_577_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_577_6530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_577_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_578_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_578_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_578_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_578_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_578_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_578_6536 ();
 DECAPx6_ASAP7_75t_R FILLER_0_578_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_578_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_579_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_579_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_579_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_579_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_579_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_579_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_580_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_580_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_580_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_580_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_580_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_580_6524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_580_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_580_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_581_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_581_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_581_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_581_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_581_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_581_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_582_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_582_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_582_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_582_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_582_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_582_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_582_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_582_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_583_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_583_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_583_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_583_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_583_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_583_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_584_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_584_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_584_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_584_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_584_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_584_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_584_6534 ();
 DECAPx6_ASAP7_75t_R FILLER_0_584_6540 ();
 DECAPx1_ASAP7_75t_R FILLER_0_584_6554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_585_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_585_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_585_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_585_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_585_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_585_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_586_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_586_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_586_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_586_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_586_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_586_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_587_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_587_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_587_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_587_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_587_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_587_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_588_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_588_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_588_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_588_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_588_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_588_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_589_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_589_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_589_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_589_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_589_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_589_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_590_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_590_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_590_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_590_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_590_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_590_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_591_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_591_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_591_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_591_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_591_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_591_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_592_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_592_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_592_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_592_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_592_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_592_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_593_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_593_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_593_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_593_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_593_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_593_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_594_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_594_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_594_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_594_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_594_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_594_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_595_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_595_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_595_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_595_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_595_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_595_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_596_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_596_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_596_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_596_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_596_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_596_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_597_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_597_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_597_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_597_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_597_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_597_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_598_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_598_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_598_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_598_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_598_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_598_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_599_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_599_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_599_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_599_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_599_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_599_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_600_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_600_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_600_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_600_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_600_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_600_6528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_600_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_600_6556 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_601_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_601_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_601_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_601_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_601_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_601_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_601_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_601_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_601_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_601_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_601_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_601_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_602_2 ();
 FILLER_ASAP7_75t_R FILLER_0_602_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_602_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_602_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_602_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_602_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_602_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_602_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_602_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_602_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_602_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_602_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_603_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_603_6 ();
 DECAPx6_ASAP7_75t_R FILLER_0_603_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_603_26 ();
 FILLER_ASAP7_75t_R FILLER_0_603_35 ();
 DECAPx10_ASAP7_75t_R FILLER_0_603_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_603_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_603_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_603_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_603_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_603_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_603_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_604_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_604_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_604_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_604_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_604_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_604_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_604_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_604_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_604_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_605_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_605_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_605_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_605_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_605_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_605_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_605_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_605_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_605_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_605_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_605_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_605_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_605_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_605_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_605_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_606_2 ();
 FILLER_ASAP7_75t_R FILLER_0_606_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_606_19 ();
 FILLER_ASAP7_75t_R FILLER_0_606_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_606_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_606_59 ();
 FILLER_ASAP7_75t_R FILLER_0_606_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_606_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_606_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_606_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_606_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_606_6530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_606_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_606_6542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_606_6546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_606_6552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_607_12 ();
 FILLER_ASAP7_75t_R FILLER_0_607_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_607_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_607_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_607_56 ();
 FILLER_ASAP7_75t_R FILLER_0_607_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_607_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_607_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_607_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_607_6530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_607_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_607_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_608_7 ();
 FILLER_ASAP7_75t_R FILLER_0_608_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_608_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_608_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_608_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_608_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_608_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_608_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_608_6534 ();
 DECAPx2_ASAP7_75t_R FILLER_0_608_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_608_6546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_608_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_609_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_609_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_609_21 ();
 DECAPx2_ASAP7_75t_R FILLER_0_609_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_609_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_609_60 ();
 FILLER_ASAP7_75t_R FILLER_0_609_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_609_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_609_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_609_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_609_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_610_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_610_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_610_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_610_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_610_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_610_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_610_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_610_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_610_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_610_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_610_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_610_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_610_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_611_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_611_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_611_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_611_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_611_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_611_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_611_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_611_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_611_6536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_611_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_612_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_612_11 ();
 DECAPx1_ASAP7_75t_R FILLER_0_612_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_612_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_612_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_612_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_612_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_612_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_612_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_612_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_612_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_613_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_613_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_613_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_613_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_613_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_613_51 ();
 FILLER_ASAP7_75t_R FILLER_0_613_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_613_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_613_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_613_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_613_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_613_6542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_613_6544 ();
 FILLER_ASAP7_75t_R FILLER_0_613_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_613_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_614_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_614_11 ();
 DECAPx2_ASAP7_75t_R FILLER_0_614_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_614_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_614_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_614_51 ();
 FILLER_ASAP7_75t_R FILLER_0_614_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_614_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_614_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_614_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_614_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_614_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_615_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_615_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_615_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_615_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_615_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_615_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_615_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_615_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_615_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_615_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_615_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_615_6539 ();
 FILLER_ASAP7_75t_R FILLER_0_615_6545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_615_6547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_616_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_616_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_616_56 ();
 FILLER_ASAP7_75t_R FILLER_0_616_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_616_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_616_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_616_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_616_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_616_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_616_6556 ();
 DECAPx2_ASAP7_75t_R FILLER_0_617_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_617_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_617_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_617_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_617_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_617_51 ();
 FILLER_ASAP7_75t_R FILLER_0_617_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_617_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_617_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_617_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_617_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_617_6532 ();
 FILLER_ASAP7_75t_R FILLER_0_617_6538 ();
 DECAPx1_ASAP7_75t_R FILLER_0_617_6545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_617_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_617_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_617_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_618_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_618_4 ();
 DECAPx2_ASAP7_75t_R FILLER_0_618_10 ();
 DECAPx4_ASAP7_75t_R FILLER_0_618_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_618_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_618_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_618_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_618_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_618_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_618_6522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_618_6533 ();
 FILLER_ASAP7_75t_R FILLER_0_618_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_618_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_619_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_619_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_619_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_619_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_619_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_619_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_619_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_619_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_619_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_619_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_619_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_619_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_619_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_620_2 ();
 FILLER_ASAP7_75t_R FILLER_0_620_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_620_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_620_51 ();
 FILLER_ASAP7_75t_R FILLER_0_620_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_620_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_620_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_620_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_620_6528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_620_6534 ();
 DECAPx4_ASAP7_75t_R FILLER_0_620_6548 ();
 DECAPx6_ASAP7_75t_R FILLER_0_621_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_621_16 ();
 FILLER_ASAP7_75t_R FILLER_0_621_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_621_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_621_56 ();
 FILLER_ASAP7_75t_R FILLER_0_621_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_621_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_621_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_621_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_621_6530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_621_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_621_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_622_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_622_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_622_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_622_44 ();
 FILLER_ASAP7_75t_R FILLER_0_622_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_622_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_622_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_622_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_622_6547 ();
 DECAPx4_ASAP7_75t_R FILLER_0_623_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_623_17 ();
 FILLER_ASAP7_75t_R FILLER_0_623_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_623_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_623_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_623_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_623_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_623_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_623_6541 ();
 DECAPx1_ASAP7_75t_R FILLER_0_623_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_623_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_623_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_624_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_624_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_624_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_624_44 ();
 FILLER_ASAP7_75t_R FILLER_0_624_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_624_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_624_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_624_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_624_6531 ();
 DECAPx4_ASAP7_75t_R FILLER_0_624_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_624_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_625_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_625_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_625_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_625_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_625_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_625_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_625_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_625_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_625_6530 ();
 FILLER_ASAP7_75t_R FILLER_0_625_6541 ();
 DECAPx4_ASAP7_75t_R FILLER_0_625_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_626_2 ();
 FILLER_ASAP7_75t_R FILLER_0_626_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_626_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_626_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_626_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_626_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_626_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_626_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_626_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_626_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_626_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_626_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_627_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_627_4 ();
 DECAPx4_ASAP7_75t_R FILLER_0_627_10 ();
 FILLER_ASAP7_75t_R FILLER_0_627_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_627_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_627_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_627_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_627_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_627_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_627_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_627_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_627_6522 ();
 DECAPx2_ASAP7_75t_R FILLER_0_627_6528 ();
 FILLER_ASAP7_75t_R FILLER_0_627_6534 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_627_6536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_627_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_627_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_627_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_628_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_628_11 ();
 DECAPx4_ASAP7_75t_R FILLER_0_628_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_628_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_628_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_628_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_628_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_628_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_628_6544 ();
 FILLER_ASAP7_75t_R FILLER_0_628_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_628_6552 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_629_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_629_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_629_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_629_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_629_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_629_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_629_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_629_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_629_6533 ();
 DECAPx4_ASAP7_75t_R FILLER_0_629_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_629_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_629_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_630_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_630_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_630_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_630_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_630_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_630_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_630_6519 ();
 FILLER_ASAP7_75t_R FILLER_0_630_6541 ();
 DECAPx1_ASAP7_75t_R FILLER_0_630_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_630_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_631_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_631_11 ();
 DECAPx1_ASAP7_75t_R FILLER_0_631_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_631_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_631_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_631_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_631_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_631_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_631_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_631_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_631_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_631_6522 ();
 DECAPx4_ASAP7_75t_R FILLER_0_631_6538 ();
 DECAPx1_ASAP7_75t_R FILLER_0_631_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_631_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_632_2 ();
 FILLER_ASAP7_75t_R FILLER_0_632_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_632_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_632_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_632_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_632_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_632_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_632_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_632_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_632_6544 ();
 FILLER_ASAP7_75t_R FILLER_0_632_6556 ();
 FILLER_ASAP7_75t_R FILLER_0_633_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_633_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_633_41 ();
 DECAPx1_ASAP7_75t_R FILLER_0_633_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_633_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_633_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_633_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_633_6516 ();
 DECAPx2_ASAP7_75t_R FILLER_0_633_6522 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_633_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_633_6534 ();
 DECAPx4_ASAP7_75t_R FILLER_0_633_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_633_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_633_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_634_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_634_4 ();
 FILLER_ASAP7_75t_R FILLER_0_634_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_634_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_634_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_634_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_634_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_634_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_634_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_634_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_634_6539 ();
 FILLER_ASAP7_75t_R FILLER_0_635_2 ();
 FILLER_ASAP7_75t_R FILLER_0_635_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_635_11 ();
 DECAPx4_ASAP7_75t_R FILLER_0_635_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_635_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_635_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_635_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_635_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_635_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_635_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_635_6538 ();
 DECAPx1_ASAP7_75t_R FILLER_0_636_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_636_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_636_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_636_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_636_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_636_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_636_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_636_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_636_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_636_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_636_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_636_6537 ();
 DECAPx4_ASAP7_75t_R FILLER_0_636_6548 ();
 DECAPx6_ASAP7_75t_R FILLER_0_637_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_637_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_637_20 ();
 DECAPx2_ASAP7_75t_R FILLER_0_637_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_637_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_637_59 ();
 FILLER_ASAP7_75t_R FILLER_0_637_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_637_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_637_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_637_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_637_6518 ();
 DECAPx1_ASAP7_75t_R FILLER_0_637_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_637_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_637_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_637_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_637_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_637_6548 ();
 DECAPx4_ASAP7_75t_R FILLER_0_638_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_638_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_638_23 ();
 FILLER_ASAP7_75t_R FILLER_0_638_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_638_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_638_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_638_59 ();
 FILLER_ASAP7_75t_R FILLER_0_638_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_638_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_638_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_638_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_638_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_638_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_638_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_638_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_639_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_639_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_639_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_639_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_639_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_639_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_639_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_639_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_639_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_639_6544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_639_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_639_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_640_2 ();
 FILLER_ASAP7_75t_R FILLER_0_640_12 ();
 FILLER_ASAP7_75t_R FILLER_0_640_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_640_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_640_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_640_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_640_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_640_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_640_6518 ();
 DECAPx4_ASAP7_75t_R FILLER_0_640_6524 ();
 FILLER_ASAP7_75t_R FILLER_0_640_6539 ();
 DECAPx2_ASAP7_75t_R FILLER_0_640_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_640_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_641_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_641_21 ();
 DECAPx2_ASAP7_75t_R FILLER_0_641_27 ();
 FILLER_ASAP7_75t_R FILLER_0_641_33 ();
 DECAPx10_ASAP7_75t_R FILLER_0_641_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_641_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_641_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_641_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_641_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_641_6542 ();
 DECAPx6_ASAP7_75t_R FILLER_0_642_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_642_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_642_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_642_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_642_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_642_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_642_6538 ();
 FILLER_ASAP7_75t_R FILLER_0_642_6544 ();
 FILLER_ASAP7_75t_R FILLER_0_642_6551 ();
 DECAPx1_ASAP7_75t_R FILLER_0_643_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_643_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_643_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_643_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_643_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_643_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_643_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_643_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_643_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_643_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_643_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_643_6548 ();
 DECAPx1_ASAP7_75t_R FILLER_0_644_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_644_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_644_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_644_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_644_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_644_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_644_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_644_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_644_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_644_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_645_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_645_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_645_44 ();
 FILLER_ASAP7_75t_R FILLER_0_645_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_645_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_645_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_645_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_645_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_645_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_645_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_645_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_645_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_646_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_646_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_646_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_646_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_646_22 ();
 DECAPx6_ASAP7_75t_R FILLER_0_646_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_646_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_646_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_646_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_646_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_646_6528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_646_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_646_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_647_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_647_24 ();
 DECAPx4_ASAP7_75t_R FILLER_0_647_46 ();
 FILLER_ASAP7_75t_R FILLER_0_647_56 ();
 DECAPx1_ASAP7_75t_R FILLER_0_647_61 ();
 DECAPx10_ASAP7_75t_R FILLER_0_647_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_647_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_647_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_648_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_648_24 ();
 DECAPx4_ASAP7_75t_R FILLER_0_648_46 ();
 FILLER_ASAP7_75t_R FILLER_0_648_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_648_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_648_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_648_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_648_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_649_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_649_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_649_46 ();
 DECAPx1_ASAP7_75t_R FILLER_0_649_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_649_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_649_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_649_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_649_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_650_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_650_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_650_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_650_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_650_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_650_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_651_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_651_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_651_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_651_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_651_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_651_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_652_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_652_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_652_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_652_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_652_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_652_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_653_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_653_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_653_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_653_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_653_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_653_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_654_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_654_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_654_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_654_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_654_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_654_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_655_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_655_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_655_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_655_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_655_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_655_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_656_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_656_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_656_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_656_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_656_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_656_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_657_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_657_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_657_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_657_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_657_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_657_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_658_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_658_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_658_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_658_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_658_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_658_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_659_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_659_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_659_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_659_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_659_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_659_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_660_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_660_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_660_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_660_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_660_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_660_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_661_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_661_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_661_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_661_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_661_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_661_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_662_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_662_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_662_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_662_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_662_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_662_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_663_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_663_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_663_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_663_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_663_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_663_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_664_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_664_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_664_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_664_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_664_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_664_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_665_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_665_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_665_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_665_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_665_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_665_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_666_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_666_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_666_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_666_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_666_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_666_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_667_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_667_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_667_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_667_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_667_6523 ();
 DECAPx4_ASAP7_75t_R FILLER_0_667_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_667_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_667_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_668_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_668_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_668_46 ();
 FILLER_ASAP7_75t_R FILLER_0_668_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_668_6494 ();
 DECAPx6_ASAP7_75t_R FILLER_0_668_6537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_668_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_668_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_669_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_669_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_669_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_669_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_669_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_669_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_670_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_670_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_670_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_670_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_670_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_670_6516 ();
 DECAPx6_ASAP7_75t_R FILLER_0_670_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_670_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_671_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_671_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_671_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_671_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_671_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_671_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_672_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_672_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_672_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_672_6513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_672_6535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_672_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_673_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_673_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_673_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_673_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_673_6506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_673_6508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_673_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_673_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_674_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_674_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_674_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_674_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_674_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_674_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_675_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_675_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_675_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_675_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_675_6502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_675_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_675_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_675_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_676_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_676_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_676_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_676_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_676_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_676_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_677_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_677_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_677_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_677_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_677_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_677_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_678_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_678_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_678_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_678_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_678_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_678_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_679_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_679_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_679_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_679_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_679_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_679_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_680_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_680_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_680_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_680_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_680_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_680_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_681_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_681_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_681_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_681_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_681_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_681_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_682_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_682_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_682_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_682_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_682_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_682_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_683_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_683_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_683_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_683_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_683_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_683_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_684_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_684_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_684_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_684_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_684_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_684_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_685_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_685_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_685_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_685_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_685_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_685_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_686_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_686_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_686_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_686_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_686_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_686_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_687_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_687_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_687_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_687_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_687_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_687_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_688_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_688_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_688_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_688_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_688_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_688_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_688_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_688_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_688_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_689_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_689_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_689_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_689_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_689_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_689_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_690_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_690_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_690_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_690_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_690_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_690_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_691_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_691_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_691_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_691_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_691_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_691_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_691_6538 ();
 DECAPx6_ASAP7_75t_R FILLER_0_691_6544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_692_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_692_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_692_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_692_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_692_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_692_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_692_6530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_692_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_693_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_693_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_693_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_693_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_693_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_693_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_694_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_694_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_694_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_694_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_694_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_694_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_694_6542 ();
 DECAPx2_ASAP7_75t_R FILLER_0_694_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_694_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_694_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_695_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_695_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_695_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_695_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_695_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_695_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_695_6530 ();
 FILLER_ASAP7_75t_R FILLER_0_695_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_695_6538 ();
 DECAPx6_ASAP7_75t_R FILLER_0_695_6544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_696_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_696_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_696_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_696_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_696_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_696_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_697_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_697_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_697_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_697_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_697_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_697_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_698_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_698_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_698_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_698_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_698_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_698_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_699_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_699_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_699_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_699_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_699_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_699_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_700_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_700_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_700_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_700_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_700_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_700_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_700_6537 ();
 DECAPx6_ASAP7_75t_R FILLER_0_700_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_700_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_701_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_701_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_701_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_701_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_701_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_701_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_702_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_702_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_702_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_702_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_702_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_702_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_703_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_703_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_703_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_703_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_703_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_703_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_704_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_704_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_704_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_704_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_704_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_704_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_705_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_705_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_705_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_705_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_705_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_705_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_705_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_705_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_705_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4622 ();
 FILLER_ASAP7_75t_R FILLER_0_706_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_4984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5050 ();
 DECAPx4_ASAP7_75t_R FILLER_0_706_5072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5084 ();
 DECAPx1_ASAP7_75t_R FILLER_0_706_5106 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_706_5110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5141 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5163 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5251 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5295 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5317 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5339 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5361 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5383 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5405 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5427 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5449 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5471 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5493 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5515 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_5537 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_706_5543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_5568 ();
 FILLER_ASAP7_75t_R FILLER_0_706_5574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5606 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5672 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5694 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5716 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5738 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5760 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5782 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5804 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5826 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5848 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5870 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5892 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5914 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5936 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5958 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_5980 ();
 DECAPx1_ASAP7_75t_R FILLER_0_706_6002 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_706_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_706_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_706_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_706_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_706_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_706_6547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_707_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_707_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_707_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_707_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_707_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_707_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_707_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_707_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_707_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_707_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_707_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_707_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_707_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_707_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_707_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_707_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_707_6542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_708_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_708_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_708_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_708_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_708_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_708_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_708_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_708_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_708_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_708_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_708_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_708_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_708_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_708_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6008 ();
 DECAPx4_ASAP7_75t_R FILLER_0_708_6030 ();
 FILLER_ASAP7_75t_R FILLER_0_708_6040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_708_6512 ();
 DECAPx1_ASAP7_75t_R FILLER_0_708_6534 ();
 DECAPx1_ASAP7_75t_R FILLER_0_708_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_708_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_708_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_708_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_709_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_709_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_709_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_709_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_709_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_709_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_709_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_709_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_709_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_709_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_709_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_709_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_709_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_709_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_709_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_709_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_709_6546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_710_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_710_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_710_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_710_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_710_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_710_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_710_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_710_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_710_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_710_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_710_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_710_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_710_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_710_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_710_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_710_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_711_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_711_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_711_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_711_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_711_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_711_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_711_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_711_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_711_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_711_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_711_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_711_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_711_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_711_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_711_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_711_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_711_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_711_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_712_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_712_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_712_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_712_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_712_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_712_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_712_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_712_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_712_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_712_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_712_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_712_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_712_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_712_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_712_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_712_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_712_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_712_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_712_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_712_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_713_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_713_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_713_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_713_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_713_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_713_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_713_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_713_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_713_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_713_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_713_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_713_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_713_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_713_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_713_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_713_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_713_6546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_714_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_714_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_714_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_714_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_714_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_714_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_714_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_714_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_714_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_714_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_714_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_714_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_714_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_714_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_714_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_714_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_714_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_714_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_714_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_715_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_715_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_715_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_715_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_715_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_715_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_715_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_715_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_715_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_715_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_715_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_715_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_715_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_715_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_715_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_715_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_715_6528 ();
 FILLER_ASAP7_75t_R FILLER_0_715_6535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_715_6542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_716_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_716_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_716_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_716_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_716_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_716_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_716_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_716_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_716_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_716_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_716_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_716_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_716_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_716_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_716_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_716_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_716_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_716_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_716_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3126 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_3148 ();
 FILLER_ASAP7_75t_R FILLER_0_717_3162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_717_3164 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3195 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_3217 ();
 FILLER_ASAP7_75t_R FILLER_0_717_3231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_717_3233 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_717_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_717_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_717_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_717_6542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_718_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_718_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_718_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_718_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_718_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_718_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_718_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_718_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_718_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_718_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_719_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_719_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_719_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_719_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_719_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_719_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_719_6546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_720_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_720_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_720_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_720_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_720_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_720_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_720_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_720_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_720_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_721_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_721_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_721_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_721_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_721_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_721_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_721_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_721_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_722_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_722_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_722_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_722_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_722_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_722_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_722_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_722_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_722_6547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_723_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_723_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_723_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_723_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_723_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_723_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_723_6537 ();
 DECAPx1_ASAP7_75t_R FILLER_0_723_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_723_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_724_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_724_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_724_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_724_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_724_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_724_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_724_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_724_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_725_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_725_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_725_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_725_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_725_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_725_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_725_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_725_6547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_726_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_726_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_726_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_726_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_726_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_726_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_726_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_726_6547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_727_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_727_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_727_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_727_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_727_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_727_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_727_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_727_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_727_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_727_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_727_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_728_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_728_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_728_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_728_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_728_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_728_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_728_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_728_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_728_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_729_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_729_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_729_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_729_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_729_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_729_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_730_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_730_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_730_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_730_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_730_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_730_6536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_730_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_730_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_731_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_731_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_731_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_731_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_731_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_732_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_732_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_732_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_732_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_732_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_732_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_733_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_733_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_733_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_733_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_733_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_733_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_734_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_734_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_734_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_734_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_734_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_734_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_735_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_735_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_735_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_735_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_735_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_735_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_736_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_736_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_736_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_736_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_736_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_736_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_737_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_737_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_737_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_737_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_737_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_737_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_738_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_738_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_738_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_738_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_738_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_738_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_739_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_739_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_739_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_739_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_739_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_739_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_740_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_740_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_740_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_740_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_740_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_740_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_741_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_741_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_741_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_741_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_741_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_741_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_742_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_742_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_742_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_742_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_742_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_742_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_743_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_743_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_743_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_743_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_743_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_743_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_744_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_744_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_744_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_744_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_744_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_744_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_745_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_745_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_745_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_745_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_745_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_745_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_746_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_746_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_746_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_746_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_746_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_746_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_747_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_747_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_747_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_747_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_747_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_747_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_747_6530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_747_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_748_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_748_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_748_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_748_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_748_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_748_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_749_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_749_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_749_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_749_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_749_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_749_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_750_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_750_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_750_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_750_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_750_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_750_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_751_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_751_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_751_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_751_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_751_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_751_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_751_6538 ();
 DECAPx6_ASAP7_75t_R FILLER_0_751_6544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_752_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_752_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_752_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_752_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_752_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_752_6518 ();
 DECAPx10_ASAP7_75t_R FILLER_0_752_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_752_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_752_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_753_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_753_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_753_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_753_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_753_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_753_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_754_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_754_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_754_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_754_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_754_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_754_6528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_754_6535 ();
 DECAPx6_ASAP7_75t_R FILLER_0_754_6544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_755_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_755_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_755_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_755_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_755_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_755_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_755_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_755_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_756_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_756_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_756_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_756_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_756_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_756_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_756_6534 ();
 DECAPx2_ASAP7_75t_R FILLER_0_756_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_756_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_756_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_757_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_757_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_757_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_757_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_757_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_757_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_758_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_758_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_758_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_758_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_758_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_758_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_759_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_759_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_759_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_759_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_759_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_759_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_760_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_760_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_760_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_760_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_760_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_760_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_761_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_761_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_761_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_761_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_761_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_761_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_762_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_762_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_762_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_762_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_762_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_762_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_763_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_763_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_763_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_763_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_763_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_763_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_764_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_764_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_764_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_764_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_764_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_764_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_765_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_765_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_765_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_765_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_765_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_765_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_766_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_766_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_766_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_766_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_766_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_766_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_767_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_767_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_767_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_767_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_767_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_767_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_768_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_768_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_768_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_768_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_768_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_768_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_769_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_769_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_769_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_769_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_769_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_769_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_770_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_770_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_770_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_770_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_770_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_770_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_771_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_771_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_771_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_771_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_771_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_771_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_772_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_772_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_772_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_772_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_772_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_772_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_773_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_773_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_773_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_773_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_773_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_773_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_774_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_774_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_774_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_774_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_774_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_774_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_775_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_775_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_775_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_775_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_775_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_775_6536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_776_2 ();
 FILLER_ASAP7_75t_R FILLER_0_776_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_776_10 ();
 DECAPx10_ASAP7_75t_R FILLER_0_776_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_776_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_776_60 ();
 FILLER_ASAP7_75t_R FILLER_0_776_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_776_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_776_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_776_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_776_6540 ();
 DECAPx4_ASAP7_75t_R FILLER_0_776_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_776_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_777_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_777_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_777_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_777_44 ();
 FILLER_ASAP7_75t_R FILLER_0_777_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_777_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_777_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_777_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_777_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_777_6556 ();
 DECAPx2_ASAP7_75t_R FILLER_0_778_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_778_13 ();
 FILLER_ASAP7_75t_R FILLER_0_778_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_778_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_778_52 ();
 FILLER_ASAP7_75t_R FILLER_0_778_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_778_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_778_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_778_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_778_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_778_6544 ();
 FILLER_ASAP7_75t_R FILLER_0_778_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_778_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_779_2 ();
 FILLER_ASAP7_75t_R FILLER_0_779_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_779_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_779_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_779_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_779_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_779_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_779_6542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_779_6544 ();
 FILLER_ASAP7_75t_R FILLER_0_779_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_779_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_780_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_780_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_780_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_780_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_780_43 ();
 FILLER_ASAP7_75t_R FILLER_0_780_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_780_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_780_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_780_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_780_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_780_6551 ();
 DECAPx1_ASAP7_75t_R FILLER_0_781_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_781_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_781_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_781_44 ();
 FILLER_ASAP7_75t_R FILLER_0_781_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_781_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_781_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_781_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_781_6530 ();
 FILLER_ASAP7_75t_R FILLER_0_781_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_781_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_781_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_781_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_782_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_782_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_782_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_782_44 ();
 FILLER_ASAP7_75t_R FILLER_0_782_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_782_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_782_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_782_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_782_6532 ();
 DECAPx2_ASAP7_75t_R FILLER_0_782_6538 ();
 FILLER_ASAP7_75t_R FILLER_0_782_6544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_782_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_782_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_783_7 ();
 DECAPx1_ASAP7_75t_R FILLER_0_783_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_783_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_783_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_783_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_783_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_783_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_783_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_783_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_783_6535 ();
 DECAPx4_ASAP7_75t_R FILLER_0_783_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_783_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_784_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_784_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_784_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_784_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_784_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_784_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_784_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_784_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_784_6524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_784_6536 ();
 DECAPx6_ASAP7_75t_R FILLER_0_785_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_785_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_785_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_785_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_785_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_785_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_785_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_785_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_785_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_785_6551 ();
 DECAPx2_ASAP7_75t_R FILLER_0_786_2 ();
 FILLER_ASAP7_75t_R FILLER_0_786_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_786_10 ();
 FILLER_ASAP7_75t_R FILLER_0_786_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_786_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_786_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_786_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_786_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_786_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_786_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_786_6547 ();
 DECAPx4_ASAP7_75t_R FILLER_0_787_2 ();
 FILLER_ASAP7_75t_R FILLER_0_787_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_787_14 ();
 DECAPx4_ASAP7_75t_R FILLER_0_787_20 ();
 FILLER_ASAP7_75t_R FILLER_0_787_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_787_32 ();
 DECAPx10_ASAP7_75t_R FILLER_0_787_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_787_60 ();
 FILLER_ASAP7_75t_R FILLER_0_787_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_787_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_787_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_787_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_787_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_788_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_788_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_788_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_788_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_788_41 ();
 DECAPx1_ASAP7_75t_R FILLER_0_788_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_788_67 ();
 DECAPx6_ASAP7_75t_R FILLER_0_788_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_788_6506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_788_6508 ();
 DECAPx2_ASAP7_75t_R FILLER_0_788_6530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_788_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_788_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_788_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_788_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_789_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_789_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_789_43 ();
 FILLER_ASAP7_75t_R FILLER_0_789_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_789_67 ();
 FILLER_ASAP7_75t_R FILLER_0_789_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_789_6541 ();
 DECAPx4_ASAP7_75t_R FILLER_0_789_6548 ();
 DECAPx4_ASAP7_75t_R FILLER_0_790_7 ();
 FILLER_ASAP7_75t_R FILLER_0_790_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_790_19 ();
 DECAPx2_ASAP7_75t_R FILLER_0_790_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_790_36 ();
 DECAPx10_ASAP7_75t_R FILLER_0_790_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_790_64 ();
 DECAPx2_ASAP7_75t_R FILLER_0_790_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_790_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_790_6542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_791_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_791_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_791_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_791_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_791_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_791_59 ();
 FILLER_ASAP7_75t_R FILLER_0_791_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_791_67 ();
 DECAPx4_ASAP7_75t_R FILLER_0_791_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_791_6533 ();
 DECAPx1_ASAP7_75t_R FILLER_0_791_6547 ();
 FILLER_ASAP7_75t_R FILLER_0_791_6556 ();
 DECAPx2_ASAP7_75t_R FILLER_0_792_2 ();
 FILLER_ASAP7_75t_R FILLER_0_792_8 ();
 FILLER_ASAP7_75t_R FILLER_0_792_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_792_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_792_44 ();
 FILLER_ASAP7_75t_R FILLER_0_792_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_792_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_792_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_792_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_792_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_792_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_793_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_793_8 ();
 FILLER_ASAP7_75t_R FILLER_0_793_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_793_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_793_43 ();
 FILLER_ASAP7_75t_R FILLER_0_793_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_793_67 ();
 DECAPx6_ASAP7_75t_R FILLER_0_793_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_793_6506 ();
 DECAPx2_ASAP7_75t_R FILLER_0_793_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_793_6544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_793_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_793_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_794_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_794_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_794_15 ();
 DECAPx2_ASAP7_75t_R FILLER_0_794_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_794_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_794_59 ();
 FILLER_ASAP7_75t_R FILLER_0_794_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_794_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_794_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_794_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_794_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_794_6534 ();
 DECAPx1_ASAP7_75t_R FILLER_0_794_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_794_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_795_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_795_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_795_32 ();
 DECAPx10_ASAP7_75t_R FILLER_0_795_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_795_60 ();
 FILLER_ASAP7_75t_R FILLER_0_795_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_795_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_795_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_795_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_795_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_795_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_796_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_796_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_796_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_796_44 ();
 FILLER_ASAP7_75t_R FILLER_0_796_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_796_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_796_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_796_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_796_6542 ();
 DECAPx6_ASAP7_75t_R FILLER_0_797_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_797_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_797_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_797_33 ();
 DECAPx4_ASAP7_75t_R FILLER_0_797_55 ();
 FILLER_ASAP7_75t_R FILLER_0_797_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_797_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_797_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_797_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_797_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_797_6526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_797_6532 ();
 DECAPx2_ASAP7_75t_R FILLER_0_797_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_797_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_797_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_797_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_798_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_798_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_798_17 ();
 FILLER_ASAP7_75t_R FILLER_0_798_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_798_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_798_56 ();
 FILLER_ASAP7_75t_R FILLER_0_798_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_798_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_798_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_798_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_798_6532 ();
 FILLER_ASAP7_75t_R FILLER_0_798_6543 ();
 DECAPx2_ASAP7_75t_R FILLER_0_798_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_798_6556 ();
 DECAPx2_ASAP7_75t_R FILLER_0_799_7 ();
 FILLER_ASAP7_75t_R FILLER_0_799_13 ();
 DECAPx4_ASAP7_75t_R FILLER_0_799_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_799_30 ();
 DECAPx10_ASAP7_75t_R FILLER_0_799_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_799_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_799_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_799_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_799_6528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_799_6544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_799_6548 ();
 DECAPx1_ASAP7_75t_R FILLER_0_799_6554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_800_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_800_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_800_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_800_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_800_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_800_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_800_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_800_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_800_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_800_6530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_800_6536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_800_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_800_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_801_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_801_11 ();
 DECAPx1_ASAP7_75t_R FILLER_0_801_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_801_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_801_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_801_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_801_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_801_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_801_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_801_6537 ();
 DECAPx1_ASAP7_75t_R FILLER_0_801_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_801_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_801_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_801_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_802_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_802_8 ();
 DECAPx2_ASAP7_75t_R FILLER_0_802_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_802_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_802_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_802_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_802_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_802_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_802_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_802_6524 ();
 DECAPx6_ASAP7_75t_R FILLER_0_802_6535 ();
 DECAPx1_ASAP7_75t_R FILLER_0_802_6549 ();
 DECAPx2_ASAP7_75t_R FILLER_0_803_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_803_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_803_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_803_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_803_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_803_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_803_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_803_6539 ();
 DECAPx1_ASAP7_75t_R FILLER_0_803_6554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_804_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_804_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_804_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_804_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_804_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_804_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_804_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_804_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_804_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_804_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_804_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_804_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_804_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_804_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_804_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_805_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_805_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_805_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_805_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_805_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_805_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_805_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_805_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_805_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_805_6543 ();
 DECAPx1_ASAP7_75t_R FILLER_0_806_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_806_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_806_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_806_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_806_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_806_51 ();
 FILLER_ASAP7_75t_R FILLER_0_806_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_806_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_806_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_806_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_806_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_806_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_806_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_806_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_806_6554 ();
 DECAPx4_ASAP7_75t_R FILLER_0_807_2 ();
 FILLER_ASAP7_75t_R FILLER_0_807_12 ();
 FILLER_ASAP7_75t_R FILLER_0_807_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_807_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_807_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_807_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_807_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_807_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_807_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_808_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_808_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_808_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_808_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_808_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_808_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_808_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_808_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_808_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_808_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_809_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_809_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_809_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_809_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_809_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_809_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_809_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_809_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_809_6533 ();
 DECAPx1_ASAP7_75t_R FILLER_0_809_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_809_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_810_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_810_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_810_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_810_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_810_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_810_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_810_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_810_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_810_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_810_6539 ();
 FILLER_ASAP7_75t_R FILLER_0_810_6549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_810_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_810_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_811_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_811_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_811_43 ();
 FILLER_ASAP7_75t_R FILLER_0_811_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_811_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_811_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_811_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_811_6533 ();
 DECAPx1_ASAP7_75t_R FILLER_0_811_6539 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_811_6543 ();
 DECAPx1_ASAP7_75t_R FILLER_0_811_6554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_812_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_812_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_812_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_812_18 ();
 FILLER_ASAP7_75t_R FILLER_0_812_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_812_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_812_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_812_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_812_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_812_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_812_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_812_6542 ();
 DECAPx2_ASAP7_75t_R FILLER_0_813_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_813_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_813_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_813_51 ();
 FILLER_ASAP7_75t_R FILLER_0_813_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_813_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_813_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_813_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_813_6528 ();
 FILLER_ASAP7_75t_R FILLER_0_813_6535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_813_6537 ();
 DECAPx4_ASAP7_75t_R FILLER_0_813_6548 ();
 DECAPx4_ASAP7_75t_R FILLER_0_814_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_814_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_814_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_814_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_814_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_814_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_814_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_814_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_814_6539 ();
 FILLER_ASAP7_75t_R FILLER_0_814_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_814_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_815_2 ();
 FILLER_ASAP7_75t_R FILLER_0_815_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_815_14 ();
 FILLER_ASAP7_75t_R FILLER_0_815_20 ();
 DECAPx1_ASAP7_75t_R FILLER_0_815_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_815_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_815_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_815_59 ();
 FILLER_ASAP7_75t_R FILLER_0_815_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_815_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_815_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_815_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_815_6520 ();
 DECAPx2_ASAP7_75t_R FILLER_0_815_6526 ();
 DECAPx4_ASAP7_75t_R FILLER_0_815_6537 ();
 FILLER_ASAP7_75t_R FILLER_0_815_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_815_6554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_816_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_816_16 ();
 FILLER_ASAP7_75t_R FILLER_0_816_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_816_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_816_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_816_52 ();
 FILLER_ASAP7_75t_R FILLER_0_816_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_816_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_816_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_816_6524 ();
 DECAPx1_ASAP7_75t_R FILLER_0_816_6531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_816_6535 ();
 DECAPx4_ASAP7_75t_R FILLER_0_816_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_816_6556 ();
 FILLER_ASAP7_75t_R FILLER_0_817_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_817_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_817_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_817_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_817_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_817_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_817_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_817_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_817_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_817_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_817_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_818_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_818_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_818_35 ();
 DECAPx4_ASAP7_75t_R FILLER_0_818_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_818_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_818_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_818_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_818_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_818_6537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_819_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_819_8 ();
 DECAPx2_ASAP7_75t_R FILLER_0_819_19 ();
 FILLER_ASAP7_75t_R FILLER_0_819_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_819_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_819_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_819_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_819_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_819_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_819_6537 ();
 FILLER_ASAP7_75t_R FILLER_0_819_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_819_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_819_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_820_2 ();
 FILLER_ASAP7_75t_R FILLER_0_820_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_820_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_820_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_820_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_820_35 ();
 DECAPx4_ASAP7_75t_R FILLER_0_820_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_820_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_820_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_820_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_820_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_820_6538 ();
 DECAPx1_ASAP7_75t_R FILLER_0_820_6544 ();
 DECAPx4_ASAP7_75t_R FILLER_0_821_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_821_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_821_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_821_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_821_51 ();
 FILLER_ASAP7_75t_R FILLER_0_821_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_821_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_821_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_821_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_821_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_821_6540 ();
 DECAPx1_ASAP7_75t_R FILLER_0_821_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_821_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_821_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_822_2 ();
 FILLER_ASAP7_75t_R FILLER_0_822_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_822_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_822_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_822_47 ();
 DECAPx1_ASAP7_75t_R FILLER_0_822_61 ();
 DECAPx10_ASAP7_75t_R FILLER_0_822_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_822_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_822_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_822_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_822_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_822_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_823_2 ();
 FILLER_ASAP7_75t_R FILLER_0_823_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_823_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_823_37 ();
 FILLER_ASAP7_75t_R FILLER_0_823_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_823_61 ();
 DECAPx10_ASAP7_75t_R FILLER_0_823_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_823_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_823_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_824_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_824_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_824_46 ();
 FILLER_ASAP7_75t_R FILLER_0_824_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_824_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_824_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_824_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_825_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_825_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_825_46 ();
 FILLER_ASAP7_75t_R FILLER_0_825_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_825_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_825_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_825_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_826_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_826_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_826_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_826_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_826_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_826_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_827_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_827_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_827_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_827_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_827_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_827_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_828_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_828_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_828_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_828_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_828_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_828_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_829_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_829_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_829_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_829_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_829_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_829_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_830_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_830_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_830_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_830_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_830_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_830_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_831_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_831_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_831_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_831_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_831_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_831_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_832_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_832_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_832_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_832_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_832_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_832_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_833_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_833_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_833_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_833_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_833_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_833_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_834_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_834_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_834_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_834_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_834_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_834_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_835_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_835_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_835_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_835_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_835_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_835_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_836_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_836_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_836_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_836_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_836_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_836_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_837_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_837_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_837_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_837_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_837_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_837_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_838_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_838_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_838_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_838_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_838_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_838_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_839_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_839_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_839_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_839_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_839_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_839_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_840_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_840_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_840_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_840_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_840_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_840_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_841_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_841_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_841_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_841_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_841_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_841_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_842_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_842_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_842_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_842_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_842_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_842_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_843_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_843_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_843_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_843_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_843_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_843_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_844_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_844_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_844_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_844_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_844_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_844_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_845_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_845_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_845_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_845_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_845_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_845_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_846_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_846_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_846_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_846_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_846_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_846_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_847_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_847_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_847_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_847_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_847_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_847_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_848_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_848_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_848_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_848_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_848_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_848_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_849_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_849_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_849_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_849_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_849_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_849_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_850_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_850_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_850_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_850_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_850_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_850_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_851_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_851_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_851_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_851_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_851_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_851_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_852_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_852_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_852_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_852_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_852_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_852_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_853_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_853_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_853_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_853_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_853_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_853_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_854_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_854_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_854_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_854_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_854_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_854_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_855_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_855_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_855_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_855_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_855_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_855_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_856_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_856_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_856_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_856_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_856_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_856_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_857_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_857_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_857_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_857_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_857_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_857_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_858_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_858_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_858_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_858_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_858_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_858_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_859_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_859_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_859_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_859_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_859_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_859_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_860_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_860_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_860_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_860_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_860_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_860_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_861_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_861_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_861_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_861_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_861_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_861_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_862_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_862_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_862_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_862_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_862_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_862_6524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_862_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_863_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_863_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_863_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_863_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_863_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_863_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_864_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_864_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_864_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_864_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_864_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_864_6524 ();
 DECAPx6_ASAP7_75t_R FILLER_0_864_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_864_6544 ();
 DECAPx1_ASAP7_75t_R FILLER_0_864_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_864_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_865_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_865_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_865_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_865_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_865_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_865_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_865_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_865_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_866_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_866_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_866_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_866_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_866_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_866_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_867_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_867_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_867_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_867_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_867_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_867_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_868_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_868_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_868_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_868_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_868_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_868_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_869_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_869_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_869_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_869_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_869_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_869_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_870_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_870_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_870_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_870_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_870_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_870_6521 ();
 DECAPx6_ASAP7_75t_R FILLER_0_870_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_870_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_871_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_871_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_871_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_871_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_871_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_871_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_872_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_872_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_872_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_872_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_872_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_872_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_872_6526 ();
 DECAPx10_ASAP7_75t_R FILLER_0_872_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_872_6554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_873_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_873_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_873_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_873_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_873_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_873_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_874_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_874_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_874_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_874_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_874_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_874_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_875_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_875_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_875_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_875_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_875_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_875_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_876_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_876_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_876_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_876_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_876_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_876_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_876_6526 ();
 DECAPx10_ASAP7_75t_R FILLER_0_876_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_876_6554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_877_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_877_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_877_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_877_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_877_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_877_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_878_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_878_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_878_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_878_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_878_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_878_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_879_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_879_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_879_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_879_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_879_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_879_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_880_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_880_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_880_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_880_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_880_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_880_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_881_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_881_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_881_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_881_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_881_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_881_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_882_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_882_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_882_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_883_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_883_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_883_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_883_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_883_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_883_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_883_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_883_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_883_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_883_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_883_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_883_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_883_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_883_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_883_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_884_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_884_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_884_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_884_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_884_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_884_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_884_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_884_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_884_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_884_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_884_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_884_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_884_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_884_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_884_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_885_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_885_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_885_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_885_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_885_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_885_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_885_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_885_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_885_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_885_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_885_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_885_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_885_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_885_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_885_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_886_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_886_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_886_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_886_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_886_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_886_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_886_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_886_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_886_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_886_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_886_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_886_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_886_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_886_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_886_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_887_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_887_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_887_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_887_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_887_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_887_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_887_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_887_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_887_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_887_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_887_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_887_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_887_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_887_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_887_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_888_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_888_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_888_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_888_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_888_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_888_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_888_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_888_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_888_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_888_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_888_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_888_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_888_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_888_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_888_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_889_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_889_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_889_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_889_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_889_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_889_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_889_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_889_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_889_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_889_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_889_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_889_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_889_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_889_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_889_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_890_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_890_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_890_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_890_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_890_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_890_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_890_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_890_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_890_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_890_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_890_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_890_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_890_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_890_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_890_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_891_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_891_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_891_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_891_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_891_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_891_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_891_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_891_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_891_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_891_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_891_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_891_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_891_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_891_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_891_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_892_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_892_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_892_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_892_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_892_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_892_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_892_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_892_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_892_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_892_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_892_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_892_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_892_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_892_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_892_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_893_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_893_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_893_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_894_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_894_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_894_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_894_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_894_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_894_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_895_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_895_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_895_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_895_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_895_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_895_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_896_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_896_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_896_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_896_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_896_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_896_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_897_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_897_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_897_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_897_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_897_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_897_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_898_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_898_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_898_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_898_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_898_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_898_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_899_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_899_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_899_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_899_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_899_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_899_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_900_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_900_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_900_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_900_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_900_6506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_900_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_900_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_900_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_901_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_901_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_901_46 ();
 DECAPx2_ASAP7_75t_R FILLER_0_901_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_901_6498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_901_6521 ();
 DECAPx6_ASAP7_75t_R FILLER_0_901_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_901_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_902_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_902_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_902_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_902_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_902_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_902_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_903_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_903_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_903_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_903_6513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_903_6535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_903_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_904_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_904_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_904_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_904_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_904_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_904_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_905_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_905_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_905_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_905_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_905_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_905_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_906_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_906_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_906_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_906_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_906_6502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_906_6525 ();
 DECAPx4_ASAP7_75t_R FILLER_0_906_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_906_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_907_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_907_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_907_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_907_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_907_6502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_907_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_907_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_907_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_908_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_908_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_908_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_908_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_908_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_909_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_909_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_909_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_909_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_909_6502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_909_6504 ();
 DECAPx10_ASAP7_75t_R FILLER_0_909_6526 ();
 DECAPx4_ASAP7_75t_R FILLER_0_909_6548 ();
 DECAPx10_ASAP7_75t_R FILLER_0_910_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_910_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_910_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_910_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_910_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_910_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_911_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_911_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_911_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_911_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_911_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_911_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_912_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_912_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_912_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_912_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_912_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_912_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_913_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_913_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_913_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_913_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_913_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_913_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_914_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_914_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_914_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_914_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_914_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_914_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_915_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_915_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_915_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_915_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_915_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_915_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_916_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_916_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_916_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_916_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_916_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_916_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_917_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_917_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_917_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_917_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_917_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_917_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_918_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_918_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_918_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_918_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_918_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_918_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_919_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_919_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_919_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_919_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_919_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_919_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_920_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_920_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_920_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_920_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_920_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_920_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_921_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_921_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_921_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_921_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_921_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_921_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_921_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_921_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_921_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_921_6554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_922_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_922_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_922_46 ();
 FILLER_ASAP7_75t_R FILLER_0_922_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_922_6502 ();
 FILLER_ASAP7_75t_R FILLER_0_922_6508 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_922_6510 ();
 DECAPx6_ASAP7_75t_R FILLER_0_922_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_922_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_922_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_923_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_923_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_923_46 ();
 FILLER_ASAP7_75t_R FILLER_0_923_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_923_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_923_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_923_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_924_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_924_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_924_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_924_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_924_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_924_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_924_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_925_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_925_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_925_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_925_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_925_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_925_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_926_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_926_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_926_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_926_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_926_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_926_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_926_6542 ();
 DECAPx2_ASAP7_75t_R FILLER_0_926_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_926_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_926_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_927_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_927_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_927_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_927_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_927_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_927_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_928_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_928_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_928_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_928_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_928_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_928_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_929_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_929_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_929_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_929_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_929_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_929_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_929_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_930_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_930_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_930_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_930_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_930_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_930_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_931_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_931_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_931_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_931_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_931_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_931_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_931_6542 ();
 DECAPx2_ASAP7_75t_R FILLER_0_931_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_931_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_931_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_932_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_932_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_932_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_932_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_932_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_932_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_933_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_933_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_933_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_933_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_933_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_933_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_934_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_934_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_934_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_934_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_934_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_934_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_935_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_935_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_935_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_935_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_935_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_935_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_936_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_936_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_936_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_936_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_936_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_936_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_937_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_937_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_937_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_937_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_937_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_937_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_938_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_938_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_938_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_938_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_938_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_938_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_939_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_939_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_939_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_939_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_939_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_939_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_940_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_940_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_940_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_940_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_940_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_940_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_941_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_941_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_941_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_941_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_941_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_941_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_942_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_942_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_942_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_942_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_942_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_942_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_943_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_943_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_943_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_943_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_943_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_943_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_944_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_944_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_944_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_944_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_944_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_944_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_945_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_945_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_945_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_945_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_945_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_945_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_946_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_946_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_946_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_946_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_946_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_946_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_947_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_947_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_947_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_947_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_947_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_947_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_948_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_948_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_948_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_948_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_948_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_948_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_949_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_949_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_949_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_949_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_949_6506 ();
 DECAPx6_ASAP7_75t_R FILLER_0_949_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_949_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_950_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_950_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_950_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_950_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_950_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_950_6554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_951_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_951_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_951_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_951_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_951_6506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_951_6520 ();
 DECAPx6_ASAP7_75t_R FILLER_0_951_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_951_6556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_952_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_952_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_952_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_952_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_952_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_952_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_952_6537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_952_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_952_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_953_2 ();
 FILLER_ASAP7_75t_R FILLER_0_953_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_953_10 ();
 FILLER_ASAP7_75t_R FILLER_0_953_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_953_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_953_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_953_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_953_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_953_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_953_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_953_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_953_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_953_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_953_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_953_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_953_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_954_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_954_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_954_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_954_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_954_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_954_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_954_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_954_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_954_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_954_6540 ();
 DECAPx1_ASAP7_75t_R FILLER_0_954_6554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_955_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_955_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_955_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_955_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_955_43 ();
 FILLER_ASAP7_75t_R FILLER_0_955_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_955_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_955_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_955_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_955_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_955_6537 ();
 DECAPx4_ASAP7_75t_R FILLER_0_955_6548 ();
 FILLER_ASAP7_75t_R FILLER_0_956_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_956_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_956_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_956_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_956_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_956_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_956_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_956_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_956_6546 ();
 DECAPx2_ASAP7_75t_R FILLER_0_957_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_957_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_957_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_957_41 ();
 DECAPx1_ASAP7_75t_R FILLER_0_957_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_957_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_957_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_957_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_957_6520 ();
 DECAPx4_ASAP7_75t_R FILLER_0_957_6527 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_957_6537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_957_6543 ();
 FILLER_ASAP7_75t_R FILLER_0_957_6549 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_957_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_957_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_958_2 ();
 FILLER_ASAP7_75t_R FILLER_0_958_16 ();
 DECAPx2_ASAP7_75t_R FILLER_0_958_23 ();
 FILLER_ASAP7_75t_R FILLER_0_958_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_958_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_958_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_958_59 ();
 FILLER_ASAP7_75t_R FILLER_0_958_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_958_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_958_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_958_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_958_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_958_6530 ();
 FILLER_ASAP7_75t_R FILLER_0_958_6536 ();
 DECAPx6_ASAP7_75t_R FILLER_0_958_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_958_6557 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_959_7 ();
 DECAPx1_ASAP7_75t_R FILLER_0_959_13 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_959_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_959_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_959_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_959_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_959_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_959_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_959_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_959_6552 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_960_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_960_13 ();
 DECAPx10_ASAP7_75t_R FILLER_0_960_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_960_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_960_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_960_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_960_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_960_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_961_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_961_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_961_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_961_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_961_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_961_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_961_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_961_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_961_6548 ();
 FILLER_ASAP7_75t_R FILLER_0_961_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_961_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_962_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_962_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_962_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_962_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_962_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_962_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_962_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_962_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_962_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_962_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_963_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_963_9 ();
 FILLER_ASAP7_75t_R FILLER_0_963_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_963_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_963_44 ();
 FILLER_ASAP7_75t_R FILLER_0_963_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_963_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_963_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_963_6536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_963_6542 ();
 DECAPx2_ASAP7_75t_R FILLER_0_964_2 ();
 FILLER_ASAP7_75t_R FILLER_0_964_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_964_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_964_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_964_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_964_52 ();
 FILLER_ASAP7_75t_R FILLER_0_964_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_964_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_964_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_964_6524 ();
 DECAPx1_ASAP7_75t_R FILLER_0_964_6530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_964_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_964_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_964_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_964_6548 ();
 DECAPx6_ASAP7_75t_R FILLER_0_965_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_965_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_965_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_965_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_965_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_965_59 ();
 FILLER_ASAP7_75t_R FILLER_0_965_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_965_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_965_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_965_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_965_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_965_6540 ();
 DECAPx2_ASAP7_75t_R FILLER_0_965_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_965_6552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_966_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_966_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_966_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_966_36 ();
 DECAPx10_ASAP7_75t_R FILLER_0_966_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_966_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_966_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_966_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_966_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_966_6548 ();
 FILLER_ASAP7_75t_R FILLER_0_966_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_966_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_967_7 ();
 FILLER_ASAP7_75t_R FILLER_0_967_13 ();
 DECAPx10_ASAP7_75t_R FILLER_0_967_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_967_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_967_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_967_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_967_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_967_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_967_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_967_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_967_6551 ();
 DECAPx1_ASAP7_75t_R FILLER_0_968_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_968_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_968_12 ();
 FILLER_ASAP7_75t_R FILLER_0_968_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_968_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_968_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_968_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_968_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_968_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_968_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_968_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_968_6535 ();
 FILLER_ASAP7_75t_R FILLER_0_968_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_968_6552 ();
 FILLER_ASAP7_75t_R FILLER_0_969_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_969_4 ();
 FILLER_ASAP7_75t_R FILLER_0_969_10 ();
 DECAPx10_ASAP7_75t_R FILLER_0_969_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_969_44 ();
 FILLER_ASAP7_75t_R FILLER_0_969_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_969_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_969_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_969_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_969_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_969_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_970_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_970_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_970_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_970_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_970_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_970_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_970_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_970_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_970_6530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_970_6541 ();
 DECAPx4_ASAP7_75t_R FILLER_0_970_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_970_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_971_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_971_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_971_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_971_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_971_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_971_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_971_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_971_6546 ();
 DECAPx6_ASAP7_75t_R FILLER_0_972_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_972_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_972_32 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_972_36 ();
 DECAPx10_ASAP7_75t_R FILLER_0_972_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_972_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_972_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_972_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_972_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_972_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_972_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_973_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_973_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_973_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_973_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_973_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_973_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_973_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_973_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_973_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_974_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_974_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_974_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_974_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_974_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_974_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_974_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_974_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_974_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_975_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_975_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_975_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_975_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_975_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_975_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_975_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_975_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_975_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_975_6540 ();
 DECAPx2_ASAP7_75t_R FILLER_0_975_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_975_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_976_2 ();
 FILLER_ASAP7_75t_R FILLER_0_976_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_976_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_976_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_976_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_976_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_976_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_976_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_976_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_976_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_976_6544 ();
 FILLER_ASAP7_75t_R FILLER_0_976_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_976_6552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_977_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_977_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_977_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_977_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_977_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_977_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_977_6524 ();
 DECAPx6_ASAP7_75t_R FILLER_0_977_6531 ();
 FILLER_ASAP7_75t_R FILLER_0_977_6545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_977_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_978_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_978_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_978_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_978_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_978_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_978_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_978_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_978_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_978_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_978_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_978_6543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_979_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_979_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_979_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_979_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_979_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_979_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_979_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_979_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_979_6548 ();
 DECAPx1_ASAP7_75t_R FILLER_0_980_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_980_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_980_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_980_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_980_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_980_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_980_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_980_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_980_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_980_6531 ();
 DECAPx6_ASAP7_75t_R FILLER_0_980_6537 ();
 FILLER_ASAP7_75t_R FILLER_0_980_6556 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_981_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_981_8 ();
 FILLER_ASAP7_75t_R FILLER_0_981_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_981_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_981_52 ();
 FILLER_ASAP7_75t_R FILLER_0_981_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_981_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_981_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_981_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_981_6539 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_981_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_981_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_981_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_982_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_982_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_982_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_982_51 ();
 FILLER_ASAP7_75t_R FILLER_0_982_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_982_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_982_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_982_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_982_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_982_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_982_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_982_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_982_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_983_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_983_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_983_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_983_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_983_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_983_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_983_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_983_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_983_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_983_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_983_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_983_6530 ();
 FILLER_ASAP7_75t_R FILLER_0_983_6536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_983_6543 ();
 DECAPx1_ASAP7_75t_R FILLER_0_983_6554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_984_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_984_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_984_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_984_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_984_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_984_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_984_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_984_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_984_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_984_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_985_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_985_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_985_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_985_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_985_52 ();
 FILLER_ASAP7_75t_R FILLER_0_985_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_985_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_985_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_985_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_985_6547 ();
 FILLER_ASAP7_75t_R FILLER_0_986_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_986_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_986_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_986_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_986_43 ();
 FILLER_ASAP7_75t_R FILLER_0_986_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_986_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_986_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_986_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_986_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_986_6530 ();
 FILLER_ASAP7_75t_R FILLER_0_986_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_986_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_986_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_986_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_987_7 ();
 FILLER_ASAP7_75t_R FILLER_0_987_13 ();
 DECAPx1_ASAP7_75t_R FILLER_0_987_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_987_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_987_56 ();
 FILLER_ASAP7_75t_R FILLER_0_987_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_987_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_987_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_987_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_987_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_987_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_987_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_987_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_988_7 ();
 FILLER_ASAP7_75t_R FILLER_0_988_13 ();
 DECAPx2_ASAP7_75t_R FILLER_0_988_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_988_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_988_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_988_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_988_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_988_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_988_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_988_6522 ();
 DECAPx4_ASAP7_75t_R FILLER_0_988_6533 ();
 DECAPx4_ASAP7_75t_R FILLER_0_988_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_989_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_989_13 ();
 FILLER_ASAP7_75t_R FILLER_0_989_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_989_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_989_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_989_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_989_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_989_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_989_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_989_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_989_6556 ();
 DECAPx2_ASAP7_75t_R FILLER_0_990_12 ();
 FILLER_ASAP7_75t_R FILLER_0_990_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_990_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_990_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_990_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_990_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_990_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_990_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_990_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_990_6540 ();
 DECAPx2_ASAP7_75t_R FILLER_0_990_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_990_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_991_2 ();
 FILLER_ASAP7_75t_R FILLER_0_991_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_991_10 ();
 FILLER_ASAP7_75t_R FILLER_0_991_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_991_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_991_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_991_33 ();
 DECAPx4_ASAP7_75t_R FILLER_0_991_55 ();
 FILLER_ASAP7_75t_R FILLER_0_991_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_991_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_991_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_991_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_991_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_991_6534 ();
 DECAPx4_ASAP7_75t_R FILLER_0_991_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_991_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_991_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_992_7 ();
 DECAPx1_ASAP7_75t_R FILLER_0_992_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_992_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_992_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_992_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_992_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_992_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_992_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_992_6518 ();
 DECAPx4_ASAP7_75t_R FILLER_0_992_6524 ();
 FILLER_ASAP7_75t_R FILLER_0_992_6534 ();
 DECAPx2_ASAP7_75t_R FILLER_0_992_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_992_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_992_6554 ();
 DECAPx4_ASAP7_75t_R FILLER_0_993_12 ();
 FILLER_ASAP7_75t_R FILLER_0_993_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_993_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_993_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_993_52 ();
 FILLER_ASAP7_75t_R FILLER_0_993_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_993_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_993_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_993_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_993_6547 ();
 DECAPx6_ASAP7_75t_R FILLER_0_994_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_994_16 ();
 FILLER_ASAP7_75t_R FILLER_0_994_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_994_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_994_35 ();
 DECAPx4_ASAP7_75t_R FILLER_0_994_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_994_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_994_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_994_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_994_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_994_6535 ();
 DECAPx4_ASAP7_75t_R FILLER_0_994_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_994_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_995_7 ();
 FILLER_ASAP7_75t_R FILLER_0_995_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_995_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_995_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_995_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_995_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_995_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_995_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_995_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_995_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_995_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_995_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_995_6548 ();
 DECAPx1_ASAP7_75t_R FILLER_0_995_6554 ();
 DECAPx6_ASAP7_75t_R FILLER_0_996_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_996_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_996_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_996_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_996_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_996_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_996_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_996_6542 ();
 DECAPx6_ASAP7_75t_R FILLER_0_997_7 ();
 DECAPx1_ASAP7_75t_R FILLER_0_997_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_997_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_997_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_997_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_997_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_997_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_997_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_997_6530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_997_6536 ();
 DECAPx2_ASAP7_75t_R FILLER_0_997_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_997_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_997_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_998_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_998_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_998_22 ();
 DECAPx6_ASAP7_75t_R FILLER_0_998_44 ();
 DECAPx2_ASAP7_75t_R FILLER_0_998_58 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_998_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_998_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_998_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_998_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_998_6551 ();
 DECAPx4_ASAP7_75t_R FILLER_0_999_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_999_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_999_32 ();
 DECAPx2_ASAP7_75t_R FILLER_0_999_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_999_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_999_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_999_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_999_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_999_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_999_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_999_6548 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1000_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1000_24 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1000_46 ();
 FILLER_ASAP7_75t_R FILLER_0_1000_56 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1000_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1000_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1000_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1000_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1001_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1001_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1001_46 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1001_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1001_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1001_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1001_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1001_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1002_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1002_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1002_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1002_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1002_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1002_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1003_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1003_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1003_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1003_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1003_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1003_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1004_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1004_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1004_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1004_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1004_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1004_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1005_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1005_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1005_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1005_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1005_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1005_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1006_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1006_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1006_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1006_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1006_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1006_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1007_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1007_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1007_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1007_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1007_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1007_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1008_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1008_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1008_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1008_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1008_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1008_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1009_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1009_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1009_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1009_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1009_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1009_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1010_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1010_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1010_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1010_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1010_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1010_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1011_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1011_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1011_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1011_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1011_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1011_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1012_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1012_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1012_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1012_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1012_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1012_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1013_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1013_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1013_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1013_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1013_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1013_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1014_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1014_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1014_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1014_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1014_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1014_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1015_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1015_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1015_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1015_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1015_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1015_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1016_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1016_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1016_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1016_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_1016_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1016_6537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1016_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1016_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1017_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1017_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1017_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1017_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1017_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1017_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1018_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1018_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1018_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1018_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_1018_6502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1018_6525 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1018_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1018_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1019_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1019_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1019_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1019_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_1019_6502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1019_6525 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1019_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1019_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1020_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1020_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1020_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1020_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1020_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1020_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1021_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1021_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1021_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1021_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1021_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1021_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1022_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1022_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1022_46 ();
 FILLER_ASAP7_75t_R FILLER_0_1022_6513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1022_6515 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1022_6537 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1022_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1022_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1023_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1023_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1023_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1023_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1023_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1023_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1024_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1024_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1024_46 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1024_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_1024_6502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1024_6504 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1024_6526 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1024_6548 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1025_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1025_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1025_46 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1025_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_1025_6506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1025_6529 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1025_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1025_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1026_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1026_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1026_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1026_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1026_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1026_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1027_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1027_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1027_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1027_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1027_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1027_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1028_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1028_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1028_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1028_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1028_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1028_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1029_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1029_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1029_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1029_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1029_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1029_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1030_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1030_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1030_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1030_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1030_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1030_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1031_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1031_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1031_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1031_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1031_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1031_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1032_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1032_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1032_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1032_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1032_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1032_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1033_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1033_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1033_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1033_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1033_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1033_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1034_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1034_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1034_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1034_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1034_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1034_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1035_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1035_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1035_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1035_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1035_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1035_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1036_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1036_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1036_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1036_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1036_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1036_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1037_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1037_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1037_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1037_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1037_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1037_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1038_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1038_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1038_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1038_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1038_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1038_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1039_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1039_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1039_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1039_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1039_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1039_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1040_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1040_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1040_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1040_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1040_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1040_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1041_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1041_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1041_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1041_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1041_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1041_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1042_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1042_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1042_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1042_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1042_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1042_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1043_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1043_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1043_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1043_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1043_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1043_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1044_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1044_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1044_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1044_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1044_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1044_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1045_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1045_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1045_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1045_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1045_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1045_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1046_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1046_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1046_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1046_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1046_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1046_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1047_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1047_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1047_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1047_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1047_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1047_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1048_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1048_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1048_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1048_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1048_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1048_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1049_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1049_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1049_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1049_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1049_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1049_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1050_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1050_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1050_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1050_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1050_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1050_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1051_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1051_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1051_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1051_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1051_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1051_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1052_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1052_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1052_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1052_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1052_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1052_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1053_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1053_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1053_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1053_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1053_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1053_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1054_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1054_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1054_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1054_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1054_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1054_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1055_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1055_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1055_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1055_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1055_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1055_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1056_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1056_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1056_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1056_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1056_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1056_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1057_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1057_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1057_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1057_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1057_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1057_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3126 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_3148 ();
 FILLER_ASAP7_75t_R FILLER_0_1058_3162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1058_3164 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3195 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_3217 ();
 FILLER_ASAP7_75t_R FILLER_0_1058_3231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1058_3233 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1058_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1058_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1058_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1059_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1059_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1059_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1059_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1059_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1059_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1059_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1059_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1059_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1059_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1059_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1059_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1059_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1059_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1059_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1060_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1060_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1060_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1060_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1060_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1060_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1060_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1060_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1060_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1060_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1060_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1060_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1060_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1060_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1060_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1061_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1061_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1061_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1061_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1061_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1061_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1061_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1061_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1061_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1061_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1061_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1061_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1061_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1061_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1061_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1062_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1062_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1062_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1062_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1062_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1062_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1062_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1062_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1062_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1062_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1062_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1062_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1062_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1062_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1062_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1063_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1063_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1063_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1063_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1063_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1063_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1063_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1063_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1063_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1063_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1063_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1063_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1063_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1063_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1063_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1064_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1064_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1064_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1064_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1064_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1064_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1064_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1064_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1064_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1064_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1064_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1064_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1064_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1064_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1064_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1065_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1065_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1065_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1065_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1065_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1065_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1065_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1065_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1065_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1065_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1065_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1065_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1065_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1065_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1065_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1066_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1066_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1066_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1066_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1066_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1066_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1066_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1066_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1066_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1066_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1066_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1066_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1066_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1066_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1066_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1067_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1067_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1067_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1067_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1067_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1067_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1067_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1067_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1067_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1067_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1067_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1067_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1067_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1067_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1067_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1068_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1068_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1068_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1068_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1068_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1068_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1068_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1068_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1068_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1068_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1068_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1068_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1068_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1068_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1068_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1069_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1069_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1069_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1674 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1069_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1818 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_1840 ();
 FILLER_ASAP7_75t_R FILLER_0_1069_1846 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1069_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2488 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1069_2510 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1069_2514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2611 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2633 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2677 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2699 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2721 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2743 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_2765 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1069_2771 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1069_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1069_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3786 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_3808 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1069_3814 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3845 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3867 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3889 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3911 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3933 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3955 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3977 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_3999 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4021 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4043 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4065 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4087 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4109 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4131 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1069_4153 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1069_4157 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4468 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_4490 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1069_4496 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4519 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4541 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4563 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4585 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1069_4607 ();
 FILLER_ASAP7_75t_R FILLER_0_1069_4617 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1069_4619 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_4622 ();
 FILLER_ASAP7_75t_R FILLER_0_1069_4628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4704 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4726 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4748 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4770 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4792 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4814 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4836 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4858 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4880 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4902 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4924 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4946 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4968 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_4990 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5012 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5034 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5056 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1069_5078 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1069_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1069_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1069_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1069_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1069_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1070_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1070_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1070_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1070_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1070_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1070_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1071_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1071_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1071_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1071_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1071_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1071_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1072_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1072_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1072_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1072_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1072_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1072_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1073_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1073_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1073_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1073_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1073_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1073_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1074_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1074_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1074_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1074_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1074_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1074_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1075_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1075_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1075_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1075_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1075_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1075_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1076_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1076_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1076_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1076_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1076_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1076_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1077_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1077_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1077_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1077_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1077_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1077_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1078_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1078_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1078_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1078_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1078_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1078_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1079_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1079_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1079_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1079_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1079_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1079_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1080_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1080_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1080_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1080_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1080_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1080_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1081_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1081_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1081_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1081_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1081_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1081_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1082_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1082_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1082_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1082_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1082_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1082_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1083_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1083_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1083_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1083_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1083_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1083_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1084_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1084_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1084_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1084_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1084_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1084_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1085_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1085_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1085_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1085_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1085_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1085_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1086_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1086_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1086_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1086_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1086_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1086_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1087_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1087_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1087_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1087_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1087_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1087_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1088_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1088_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1088_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1088_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1088_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1088_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1089_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1089_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1089_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1089_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1089_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1089_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1090_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1090_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1090_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1090_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1090_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1090_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1091_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1091_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1091_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1091_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1091_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1091_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1092_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1092_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1092_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1092_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1092_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1092_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1093_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1093_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1093_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1093_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1093_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1093_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1094_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1094_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1094_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1094_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1094_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1094_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1095_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1095_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1095_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1095_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1095_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1095_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1096_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1096_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1096_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1096_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1096_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1096_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1097_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1097_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1097_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1097_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1097_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1097_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1098_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1098_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1098_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1098_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1098_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1098_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1099_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1099_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1099_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1099_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1099_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1099_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1100_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1100_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1100_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1100_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1100_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1100_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1101_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1101_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1101_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1101_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1101_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1101_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1102_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1102_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1102_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1102_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1102_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1102_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1103_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1103_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1103_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1103_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1103_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1103_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1104_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1104_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1104_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1104_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1104_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1104_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1105_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1105_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1105_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1105_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1105_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1105_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1106_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1106_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1106_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1106_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1106_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1106_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1107_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1107_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1107_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1107_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1107_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1107_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1108_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1108_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1108_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1108_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1108_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1108_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1109_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1109_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1109_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1109_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1109_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1109_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1110_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1110_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1110_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1110_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1110_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1110_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1111_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1111_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1111_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1111_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1111_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1111_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1112_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1112_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1112_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1112_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1112_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1112_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1113_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1113_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1113_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1113_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1113_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1113_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1114_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1114_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1114_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1114_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1114_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1114_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1115_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1115_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1115_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1115_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1115_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1115_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1116_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1116_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1116_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1116_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1116_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1116_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1117_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1117_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1117_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1117_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1117_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1117_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1118_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1118_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1118_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1118_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1118_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1118_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1119_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1119_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1119_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1119_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1119_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1119_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1120_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1120_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1120_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1120_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1120_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1120_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1121_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1121_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1121_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1121_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1121_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1121_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1122_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1122_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1122_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1122_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1122_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1122_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1123_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1123_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1123_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1123_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1123_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1123_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1124_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1124_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1124_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1124_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1124_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1124_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1125_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1125_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1125_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1125_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1125_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1125_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1126_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1126_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1126_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1126_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1126_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1126_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1127_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1127_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1127_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1127_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1127_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1127_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_1128_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1128_9 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1128_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1128_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1128_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1128_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1128_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1128_6528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1128_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_1128_6556 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1129_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1129_8 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1129_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1129_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1129_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1129_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1129_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1129_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1129_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1129_6522 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1129_6528 ();
 FILLER_ASAP7_75t_R FILLER_0_1129_6534 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1129_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_1129_6556 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1130_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1130_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1130_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1130_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1130_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1130_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1130_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1130_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1130_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1130_6542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1130_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1131_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1131_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1131_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1131_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1131_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1131_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1131_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1131_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1131_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1131_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1131_6530 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1131_6541 ();
 FILLER_ASAP7_75t_R FILLER_0_1131_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1131_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1132_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1132_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1132_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1132_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1132_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1132_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1132_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1132_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1132_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1132_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1132_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1133_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1133_8 ();
 FILLER_ASAP7_75t_R FILLER_0_1133_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1133_21 ();
 FILLER_ASAP7_75t_R FILLER_0_1133_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1133_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1133_56 ();
 FILLER_ASAP7_75t_R FILLER_0_1133_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1133_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1133_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1133_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1133_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1133_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1133_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1133_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1134_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1134_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1134_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1134_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1134_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1134_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1134_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_1134_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1134_6516 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1134_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1134_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1135_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1135_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1135_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1135_44 ();
 FILLER_ASAP7_75t_R FILLER_0_1135_66 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1135_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1135_6502 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1135_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1135_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1135_6544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1136_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1136_13 ();
 FILLER_ASAP7_75t_R FILLER_0_1136_19 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1136_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1136_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1136_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1136_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1136_67 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1136_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_1136_6502 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1136_6525 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1136_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_1136_6551 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1137_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1137_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1137_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1137_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1137_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1137_67 ();
 FILLER_ASAP7_75t_R FILLER_0_1137_6492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1137_6494 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1137_6516 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1137_6530 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1137_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1137_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1137_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1137_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1138_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1138_12 ();
 FILLER_ASAP7_75t_R FILLER_0_1138_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1138_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1138_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1138_67 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1138_6492 ();
 FILLER_ASAP7_75t_R FILLER_0_1138_6502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1138_6504 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1138_6531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1138_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1138_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1138_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1138_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1139_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1139_8 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1139_14 ();
 FILLER_ASAP7_75t_R FILLER_0_1139_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1139_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1139_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1139_59 ();
 FILLER_ASAP7_75t_R FILLER_0_1139_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1139_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1139_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1139_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1139_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1139_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1139_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_1140_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1140_9 ();
 FILLER_ASAP7_75t_R FILLER_0_1140_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1140_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1140_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1140_67 ();
 FILLER_ASAP7_75t_R FILLER_0_1140_6513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1140_6515 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1140_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_1141_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1141_4 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1141_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1141_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1141_59 ();
 FILLER_ASAP7_75t_R FILLER_0_1141_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1141_67 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1141_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1141_6517 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1141_6531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1141_6535 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1141_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1141_6547 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1142_7 ();
 FILLER_ASAP7_75t_R FILLER_0_1142_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1142_23 ();
 FILLER_ASAP7_75t_R FILLER_0_1142_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1142_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1142_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1142_59 ();
 FILLER_ASAP7_75t_R FILLER_0_1142_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1142_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1142_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1142_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1142_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1142_6526 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1142_6532 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1142_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1142_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1142_6552 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1143_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1143_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1143_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1143_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1143_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1143_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1143_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1143_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1143_6530 ();
 FILLER_ASAP7_75t_R FILLER_0_1143_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1143_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1143_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1143_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1144_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1144_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1144_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1144_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1144_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1144_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1144_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1144_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1144_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1144_6539 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1144_6550 ();
 FILLER_ASAP7_75t_R FILLER_0_1144_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1145_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1145_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1145_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1145_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1145_51 ();
 FILLER_ASAP7_75t_R FILLER_0_1145_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1145_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1145_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1145_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1145_6524 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1145_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_1145_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1145_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1146_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1146_8 ();
 FILLER_ASAP7_75t_R FILLER_0_1146_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1146_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1146_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1146_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1146_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1146_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1146_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1146_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1146_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_1146_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1146_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1146_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1146_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1147_7 ();
 FILLER_ASAP7_75t_R FILLER_0_1147_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1147_23 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1147_29 ();
 FILLER_ASAP7_75t_R FILLER_0_1147_35 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1147_42 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1147_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1147_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1147_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1147_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1147_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1147_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1148_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1148_11 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1148_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1148_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1148_51 ();
 FILLER_ASAP7_75t_R FILLER_0_1148_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1148_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1148_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1148_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1148_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1149_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1149_13 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1149_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1149_41 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1149_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1149_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1149_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1149_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1149_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1149_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1150_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1150_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1150_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1150_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1150_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1150_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1150_6538 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1150_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1150_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1151_7 ();
 FILLER_ASAP7_75t_R FILLER_0_1151_13 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1151_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1151_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1151_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1151_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1151_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1151_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1151_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1151_6543 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1151_6554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1152_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1152_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1152_17 ();
 FILLER_ASAP7_75t_R FILLER_0_1152_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1152_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1152_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1152_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1152_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1152_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1152_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1152_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1152_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_1153_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1153_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1153_41 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1153_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1153_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1153_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1153_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1153_6524 ();
 FILLER_ASAP7_75t_R FILLER_0_1153_6531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1153_6538 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1153_6544 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1154_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1154_16 ();
 FILLER_ASAP7_75t_R FILLER_0_1154_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1154_35 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1154_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1154_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1154_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1154_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1154_6528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1154_6534 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1154_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1154_6544 ();
 FILLER_ASAP7_75t_R FILLER_0_1154_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1154_6552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1155_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1155_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1155_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1155_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1155_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1155_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1155_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_1155_6546 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1156_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1156_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1156_14 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1156_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1156_26 ();
 FILLER_ASAP7_75t_R FILLER_0_1156_32 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1156_39 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1156_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1156_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1156_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1156_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1156_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1156_6530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1156_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_1156_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1157_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1157_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1157_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1157_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1157_33 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1157_55 ();
 FILLER_ASAP7_75t_R FILLER_0_1157_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1157_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1157_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1157_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1157_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1157_6542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1157_6546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1157_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1158_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1158_11 ();
 FILLER_ASAP7_75t_R FILLER_0_1158_17 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1158_24 ();
 FILLER_ASAP7_75t_R FILLER_0_1158_30 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1158_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1158_59 ();
 FILLER_ASAP7_75t_R FILLER_0_1158_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1158_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1158_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1158_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1158_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1158_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1158_6547 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1159_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1159_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1159_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1159_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1159_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1159_56 ();
 FILLER_ASAP7_75t_R FILLER_0_1159_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1159_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1159_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1159_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1159_6522 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1159_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1159_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1159_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1159_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1160_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1160_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1160_10 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1160_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1160_43 ();
 FILLER_ASAP7_75t_R FILLER_0_1160_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1160_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1160_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1160_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1160_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1160_6522 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1160_6528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1160_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_1160_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1161_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1161_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1161_14 ();
 FILLER_ASAP7_75t_R FILLER_0_1161_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1161_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1161_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1161_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1161_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1161_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1161_6522 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1161_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1161_6543 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1162_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1162_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1162_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1162_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1162_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1162_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1162_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1162_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1162_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1162_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1162_6552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1163_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1163_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1163_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1163_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1163_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1163_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1163_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1163_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1163_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1163_6522 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1163_6528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1163_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1163_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1164_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1164_11 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1164_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1164_32 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1164_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1164_60 ();
 FILLER_ASAP7_75t_R FILLER_0_1164_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1164_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1164_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1164_6533 ();
 FILLER_ASAP7_75t_R FILLER_0_1164_6543 ();
 FILLER_ASAP7_75t_R FILLER_0_1164_6550 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1164_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1165_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1165_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1165_14 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1165_20 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1165_24 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1165_30 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1165_34 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1165_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1165_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1165_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1165_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1165_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1165_6537 ();
 FILLER_ASAP7_75t_R FILLER_0_1165_6551 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1166_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1166_16 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1166_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1166_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1166_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1166_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1166_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1166_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1166_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1166_6530 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1166_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1166_6540 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1166_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1166_6557 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1167_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1167_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1167_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1167_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1167_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1167_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1167_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1167_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1167_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_1167_6545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1167_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1167_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1167_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1168_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1168_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1168_35 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1168_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1168_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1168_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1168_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1168_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1168_6542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1168_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1169_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1169_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1169_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1169_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1169_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1169_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1169_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1169_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1169_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1170_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1170_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1170_17 ();
 FILLER_ASAP7_75t_R FILLER_0_1170_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1170_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1170_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1170_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1170_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1170_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1170_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1170_6536 ();
 FILLER_ASAP7_75t_R FILLER_0_1170_6546 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1171_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1171_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1171_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1171_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1171_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1171_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1171_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1171_6539 ();
 FILLER_ASAP7_75t_R FILLER_0_1171_6545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1171_6547 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1172_7 ();
 FILLER_ASAP7_75t_R FILLER_0_1172_13 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1172_25 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1172_47 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1172_61 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1172_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1172_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1172_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1172_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1172_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1172_6547 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1173_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1173_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1173_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1173_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1173_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1173_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1173_6529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1173_6535 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1173_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_1173_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1174_7 ();
 FILLER_ASAP7_75t_R FILLER_0_1174_17 ();
 FILLER_ASAP7_75t_R FILLER_0_1174_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1174_31 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1174_53 ();
 FILLER_ASAP7_75t_R FILLER_0_1174_63 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1174_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1174_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1174_6541 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1174_6548 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1175_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1175_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1175_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1175_32 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1175_54 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1175_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1175_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1175_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1175_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1175_6536 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1175_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1175_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1176_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1176_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1176_46 ();
 FILLER_ASAP7_75t_R FILLER_0_1176_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1176_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1176_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1176_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1177_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1177_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1177_46 ();
 FILLER_ASAP7_75t_R FILLER_0_1177_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1177_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1177_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1177_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1178_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1178_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1178_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1178_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1178_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1178_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1179_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1179_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1179_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1179_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1179_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1179_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1180_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1180_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1180_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1180_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1180_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1180_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1181_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1181_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1181_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1181_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1181_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1181_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1182_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1182_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1182_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1182_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1182_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1182_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1183_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1183_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1183_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1183_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1183_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1183_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1184_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1184_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1184_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1184_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1184_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1184_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1185_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1185_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1185_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1185_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1185_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1185_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1186_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1186_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1186_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1186_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1186_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1186_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1187_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1187_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1187_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1187_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1187_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1187_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1188_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1188_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1188_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1188_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1188_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1188_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1189_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1189_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1189_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1189_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1189_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1189_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1190_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1190_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1190_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1190_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1190_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1190_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1191_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1191_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1191_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1191_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1191_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1191_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1192_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1192_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1192_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1192_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1192_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1192_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1193_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1193_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1193_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1193_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1193_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1193_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1194_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1194_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1194_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1194_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1194_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1194_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1195_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1195_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1195_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1195_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1195_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1195_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1196_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1196_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1196_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1196_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1196_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1196_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1197_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1197_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1197_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1197_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1197_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1197_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1198_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1198_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1198_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1198_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1198_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1198_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1199_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1199_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1199_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1199_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1199_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1199_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1200_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1200_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1200_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1200_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1200_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1200_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1201_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1201_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1201_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1201_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1201_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1201_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1202_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1202_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1202_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1202_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1202_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1202_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1203_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1203_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1203_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1203_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1203_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1203_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1204_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1204_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1204_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1204_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1204_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1204_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1205_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1205_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1205_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1205_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1205_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1205_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1206_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1206_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1206_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1206_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1206_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1206_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1207_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1207_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1207_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1207_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1207_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1207_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1208_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1208_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1208_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1208_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1208_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1208_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1209_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1209_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1209_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1209_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1209_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1209_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1210_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1210_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1210_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1210_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1210_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1210_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1211_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1211_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1211_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1211_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1211_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1211_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1212_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1212_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1212_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1212_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1212_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1212_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1213_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1213_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1213_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1213_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1213_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1213_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1214_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1214_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1214_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1214_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1214_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1214_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1215_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1215_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1215_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1215_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1215_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1215_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1216_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1216_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1216_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1216_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1216_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1216_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1217_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1217_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1217_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1217_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1217_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1217_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1218_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1218_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1218_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1218_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1218_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1218_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1219_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1219_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1219_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1219_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1219_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1219_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1220_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1220_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1220_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1220_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1220_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1220_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1221_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1221_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1221_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1221_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1221_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1221_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1222_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1222_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1222_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1222_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1222_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1222_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1223_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1223_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1223_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1223_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1223_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1223_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1224_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1224_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1224_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1224_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1224_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1224_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1225_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1225_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1225_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1225_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1225_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1225_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1226_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1226_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1226_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1226_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1226_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1226_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1227_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1227_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1227_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1227_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1227_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1227_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1228_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1228_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1228_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1228_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1228_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1228_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1229_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1229_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1229_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1229_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1229_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1229_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1230_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1230_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1230_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1230_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1230_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1230_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1231_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1231_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1231_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1231_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1231_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1231_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1232_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1232_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1232_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1232_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1232_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1232_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1233_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1233_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1233_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1233_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1233_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1233_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1674 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_1696 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_1710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1746 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1768 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1790 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1812 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_1834 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_4982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5048 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1234_5070 ();
 FILLER_ASAP7_75t_R FILLER_0_1234_5080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1234_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1234_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1234_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1235_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1235_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1235_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1235_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1235_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1235_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1235_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1235_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1235_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1235_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1235_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1235_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1235_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1235_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1235_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1236_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1236_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1236_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1236_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1236_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1236_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1236_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1236_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1236_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1236_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1236_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1236_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1236_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1236_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1236_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1237_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1237_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1237_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1237_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1237_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1237_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1237_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1237_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1237_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1237_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1237_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1237_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1237_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1237_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1237_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1238_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1238_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1238_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1238_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1238_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1238_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1238_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1238_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1238_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1238_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1238_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1238_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1238_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1238_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1238_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1239_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1239_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1239_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1239_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1239_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1239_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1239_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1239_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1239_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1239_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1239_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1239_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1239_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1239_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1239_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1240_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1240_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1240_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1240_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1240_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1240_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1240_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1240_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1240_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1240_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1240_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1240_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1240_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1240_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1240_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1241_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1241_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1241_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1241_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1241_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1241_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1241_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1241_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1241_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1241_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1241_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1241_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1241_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1241_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1241_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1242_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1242_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1242_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1242_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1242_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1242_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1242_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1242_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1242_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1242_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1242_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1242_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1242_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1242_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1242_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1243_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1243_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1243_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1243_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1243_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1243_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1243_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1243_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1243_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1243_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1243_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1243_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1243_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1243_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1243_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1244_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1244_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1244_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1244_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1244_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1244_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1244_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1244_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1244_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1244_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1244_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1244_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1244_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1244_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1244_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5128 ();
 FILLER_ASAP7_75t_R FILLER_0_1245_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_5536 ();
 FILLER_ASAP7_75t_R FILLER_0_1245_5542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1245_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1245_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1245_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1246_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1246_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1246_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1246_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1246_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1246_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1247_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1247_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1247_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1247_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1247_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1247_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1248_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1248_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1248_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1248_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1248_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1248_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1249_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1249_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1249_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1249_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1249_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1249_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1250_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1250_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1250_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1250_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1250_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1250_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1251_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1251_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1251_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1251_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1251_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1251_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1252_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1252_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1252_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1252_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1252_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1252_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1253_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1253_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1253_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1253_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1253_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1253_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1254_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1254_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1254_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1254_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1254_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1254_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1255_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1255_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1255_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1255_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1255_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1255_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1256_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1256_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1256_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1256_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1256_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1256_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1257_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1257_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1257_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1257_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1257_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1257_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1258_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1258_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1258_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1258_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1258_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1258_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1259_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1259_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1259_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1259_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1259_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1259_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1260_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1260_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1260_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1260_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1260_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1260_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1261_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1261_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1261_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1261_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1261_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1261_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1262_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1262_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1262_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1262_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1262_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1262_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1263_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1263_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1263_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1263_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1263_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1263_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1264_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1264_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1264_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1264_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1264_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1264_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1265_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1265_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1265_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1265_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1265_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1265_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1266_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1266_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1266_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1266_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1266_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1266_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1267_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1267_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1267_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1267_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1267_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1267_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1268_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1268_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1268_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1268_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1268_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1268_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1269_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1269_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1269_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1269_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1269_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1269_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1270_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1270_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1270_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1270_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1270_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1270_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1271_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1271_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1271_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1271_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1271_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1271_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1272_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1272_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1272_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1272_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1272_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1272_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1273_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1273_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1273_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1273_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1273_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1273_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1274_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1274_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1274_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1274_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1274_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1274_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1275_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1275_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1275_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1275_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1275_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1275_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1276_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1276_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1276_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1276_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1276_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1276_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1277_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1277_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1277_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1277_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1277_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1277_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1278_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1278_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1278_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1278_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1278_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1278_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1279_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1279_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1279_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1279_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1279_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1279_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1280_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1280_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1280_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1280_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1280_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1280_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1281_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1281_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1281_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1281_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1281_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1281_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1282_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1282_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1282_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1282_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1282_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1282_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1283_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1283_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1283_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1283_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1283_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1283_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1284_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1284_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1284_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1284_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1284_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1284_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1285_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1285_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1285_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1285_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1285_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1285_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1286_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1286_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1286_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1286_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1286_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1286_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1287_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1287_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1287_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1287_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1287_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1287_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1288_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1288_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1288_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1288_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1288_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1288_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1289_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1289_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1289_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1289_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1289_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1289_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1290_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1290_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1290_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1290_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1290_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1290_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1291_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1291_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1291_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1291_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1291_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1291_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1292_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1292_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1292_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1292_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1292_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1292_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1293_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1293_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1293_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1293_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1293_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1293_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1294_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1294_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1294_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1294_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1294_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1294_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1295_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1295_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1295_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1295_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1295_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1295_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1296_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1296_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1296_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1296_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1296_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1296_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1297_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1297_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1297_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1297_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1297_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1297_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1298_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1298_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1298_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1298_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1298_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1298_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1299_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1299_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1299_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1299_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1299_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1299_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1300_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1300_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1300_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1300_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1300_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1300_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1301_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1301_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1301_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1301_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1301_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1301_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1302_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1302_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1302_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1302_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1302_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1302_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1303_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1303_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1303_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1303_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1303_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1303_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1304_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1304_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1304_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1304_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1304_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1304_6528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1304_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_1304_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1305_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1305_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1305_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1305_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1305_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1305_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1305_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1305_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1305_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1305_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_1305_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_1305_6556 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1306_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1306_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1306_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1306_41 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1306_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1306_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1306_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1306_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1306_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1306_6539 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1306_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_1306_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1306_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1307_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1307_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1307_10 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1307_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1307_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1307_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1307_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1307_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1307_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1307_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1307_6528 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1307_6534 ();
 FILLER_ASAP7_75t_R FILLER_0_1307_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1307_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1307_6548 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1308_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1308_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1308_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1308_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1308_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1308_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1308_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1308_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1308_6528 ();
 FILLER_ASAP7_75t_R FILLER_0_1308_6534 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1308_6536 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1308_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_1308_6556 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1309_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1309_17 ();
 FILLER_ASAP7_75t_R FILLER_0_1309_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1309_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1309_56 ();
 FILLER_ASAP7_75t_R FILLER_0_1309_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1309_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1309_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1309_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1309_6522 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1309_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1309_6532 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1309_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1309_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1310_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1310_11 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1310_22 ();
 FILLER_ASAP7_75t_R FILLER_0_1310_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1310_35 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1310_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1310_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1310_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1310_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1310_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1310_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1310_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1310_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1310_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1310_6552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1311_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1311_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1311_45 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1311_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1311_6492 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1311_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1311_6518 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1311_6524 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1311_6530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1311_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1311_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1311_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1312_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1312_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1312_10 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1312_16 ();
 FILLER_ASAP7_75t_R FILLER_0_1312_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1312_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1312_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1312_52 ();
 FILLER_ASAP7_75t_R FILLER_0_1312_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1312_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1312_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1312_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1312_6543 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1313_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1313_8 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1313_14 ();
 FILLER_ASAP7_75t_R FILLER_0_1313_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1313_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1313_59 ();
 FILLER_ASAP7_75t_R FILLER_0_1313_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1313_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1313_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1313_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1313_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1313_6532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1313_6543 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1314_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1314_11 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1314_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1314_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1314_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1314_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1314_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1314_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1314_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1314_6552 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1315_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1315_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1315_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1315_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1315_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1315_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1315_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1315_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1315_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1315_6530 ();
 FILLER_ASAP7_75t_R FILLER_0_1315_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1315_6548 ();
 FILLER_ASAP7_75t_R FILLER_0_1316_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1316_4 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1316_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1316_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1316_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1316_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1316_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1316_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1316_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1316_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1316_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1316_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1317_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1317_6 ();
 FILLER_ASAP7_75t_R FILLER_0_1317_12 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1317_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1317_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1317_56 ();
 FILLER_ASAP7_75t_R FILLER_0_1317_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1317_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1317_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1317_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1317_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1317_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1317_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1318_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1318_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1318_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1318_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1318_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1318_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1318_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1318_6524 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1318_6531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1318_6535 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1318_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_1318_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1319_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1319_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1319_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1319_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1319_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1319_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1319_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1319_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1319_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1319_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1319_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1319_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1319_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1320_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1320_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1320_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1320_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1320_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1320_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1320_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1320_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1320_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1320_6537 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1320_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1321_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1321_13 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1321_33 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1321_55 ();
 FILLER_ASAP7_75t_R FILLER_0_1321_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1321_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1321_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1321_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1321_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1321_6542 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1322_7 ();
 FILLER_ASAP7_75t_R FILLER_0_1322_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1322_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1322_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1322_56 ();
 FILLER_ASAP7_75t_R FILLER_0_1322_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1322_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1322_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1322_6541 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1322_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1322_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1322_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1323_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1323_6 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1323_12 ();
 FILLER_ASAP7_75t_R FILLER_0_1323_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1323_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1323_60 ();
 FILLER_ASAP7_75t_R FILLER_0_1323_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1323_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1323_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1323_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1323_6552 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1324_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1324_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1324_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1324_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1324_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1324_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1324_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1324_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1324_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1324_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1324_6525 ();
 FILLER_ASAP7_75t_R FILLER_0_1324_6540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1324_6542 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1324_6548 ();
 FILLER_ASAP7_75t_R FILLER_0_1325_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1325_4 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1325_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1325_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1325_59 ();
 FILLER_ASAP7_75t_R FILLER_0_1325_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1325_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1325_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1325_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1325_6536 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1325_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1325_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1326_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1326_17 ();
 FILLER_ASAP7_75t_R FILLER_0_1326_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1326_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1326_31 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1326_53 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1326_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1326_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1326_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1326_6524 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1326_6531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1326_6545 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1326_6551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1326_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1327_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1327_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1327_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1327_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1327_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1327_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1327_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1327_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1327_6529 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1327_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1327_6552 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1328_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1328_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1328_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1328_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1328_56 ();
 FILLER_ASAP7_75t_R FILLER_0_1328_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1328_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1328_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1328_6536 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1328_6548 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1329_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1329_13 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1329_35 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1329_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1329_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1329_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1329_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1329_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1329_6539 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1329_6554 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1330_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1330_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1330_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1330_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1330_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1330_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1330_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1330_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1330_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1330_6522 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1330_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1330_6537 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1330_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1330_6557 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1331_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1331_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1331_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1331_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1331_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1331_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1331_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1331_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1331_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1331_6522 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1331_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1331_6532 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1331_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1331_6552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1332_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1332_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1332_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1332_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1332_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1332_51 ();
 FILLER_ASAP7_75t_R FILLER_0_1332_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1332_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1332_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1332_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1332_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1332_6522 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1332_6528 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1332_6548 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1333_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1333_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1333_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1333_18 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1333_24 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1333_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1333_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1333_56 ();
 FILLER_ASAP7_75t_R FILLER_0_1333_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1333_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1333_6514 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1333_6546 ();
 FILLER_ASAP7_75t_R FILLER_0_1333_6556 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1334_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1334_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1334_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1334_28 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1334_50 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1334_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1334_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1334_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1334_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1334_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_1334_6551 ();
 FILLER_ASAP7_75t_R FILLER_0_1335_2 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1335_9 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1335_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1335_37 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1335_59 ();
 FILLER_ASAP7_75t_R FILLER_0_1335_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1335_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1335_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1335_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1335_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1335_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1335_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_1335_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1335_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1336_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1336_13 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1336_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1336_41 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1336_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1336_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1336_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1336_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1336_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1336_6532 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1336_6538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1336_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1336_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1336_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1337_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1337_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1337_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1337_16 ();
 FILLER_ASAP7_75t_R FILLER_0_1337_22 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1337_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1337_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1337_52 ();
 FILLER_ASAP7_75t_R FILLER_0_1337_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1337_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1337_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1337_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1337_6530 ();
 FILLER_ASAP7_75t_R FILLER_0_1337_6541 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1337_6548 ();
 FILLER_ASAP7_75t_R FILLER_0_1338_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1338_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1338_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1338_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1338_52 ();
 FILLER_ASAP7_75t_R FILLER_0_1338_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1338_6492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1338_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1338_6520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1338_6522 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1338_6528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1338_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_1338_6551 ();
 FILLER_ASAP7_75t_R FILLER_0_1339_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1339_4 ();
 FILLER_ASAP7_75t_R FILLER_0_1339_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1339_12 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1339_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1339_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1339_34 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1339_56 ();
 FILLER_ASAP7_75t_R FILLER_0_1339_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1339_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1339_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1339_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1339_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_1339_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1339_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1339_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1340_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1340_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1340_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1340_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1340_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1340_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1340_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1340_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1340_6534 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1340_6540 ();
 FILLER_ASAP7_75t_R FILLER_0_1340_6546 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1341_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1341_12 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1341_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1341_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1341_30 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1341_52 ();
 FILLER_ASAP7_75t_R FILLER_0_1341_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1341_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1341_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1341_6524 ();
 FILLER_ASAP7_75t_R FILLER_0_1341_6531 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1341_6538 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1341_6544 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1342_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1342_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1342_40 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1342_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1342_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1342_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1342_6533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1342_6537 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1342_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1342_6547 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1342_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1342_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1343_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1343_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1343_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1343_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1343_32 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1343_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1343_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1343_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1343_6528 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1343_6534 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1343_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1343_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_1343_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1343_6557 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1344_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1344_6 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1344_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1344_44 ();
 FILLER_ASAP7_75t_R FILLER_0_1344_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1344_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1344_6514 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1344_6528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1344_6532 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1344_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1344_6557 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1345_2 ();
 FILLER_ASAP7_75t_R FILLER_0_1345_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1345_10 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1345_26 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1345_48 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1345_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1345_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1345_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1345_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1345_6538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1345_6549 ();
 FILLER_ASAP7_75t_R FILLER_0_1345_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1345_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_1346_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1346_4 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1346_10 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1346_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1346_38 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1346_60 ();
 FILLER_ASAP7_75t_R FILLER_0_1346_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1346_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1346_6514 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1346_6543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1346_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1347_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1347_17 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1347_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1347_30 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1347_36 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1347_58 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1347_6492 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1347_6514 ();
 FILLER_ASAP7_75t_R FILLER_0_1347_6524 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1347_6531 ();
 FILLER_ASAP7_75t_R FILLER_0_1347_6546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1347_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1347_6557 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1348_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1348_27 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1348_49 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1348_63 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1348_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1348_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1348_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1348_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1348_6542 ();
 FILLER_ASAP7_75t_R FILLER_0_1349_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1349_4 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1349_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1349_14 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1349_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1349_35 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1349_57 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1349_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1349_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1349_6514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1349_6528 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1349_6544 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1350_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1350_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1350_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1350_29 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1350_51 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1350_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1350_6514 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1350_6536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1350_6542 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1350_6553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1350_6557 ();
 FILLER_ASAP7_75t_R FILLER_0_1351_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1351_9 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1351_31 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1351_53 ();
 FILLER_ASAP7_75t_R FILLER_0_1351_59 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1351_61 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1351_6492 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1351_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1351_6533 ();
 FILLER_ASAP7_75t_R FILLER_0_1351_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1351_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1352_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1352_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1352_46 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1352_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1352_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1352_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1352_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1352_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1353_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1353_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1353_46 ();
 FILLER_ASAP7_75t_R FILLER_0_1353_60 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1353_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1353_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1353_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1354_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1354_24 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1354_46 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1354_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1354_64 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1354_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1354_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1354_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1355_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1355_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1355_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1355_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1355_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1355_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1356_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1356_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1356_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1356_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1356_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1356_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1357_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1357_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1357_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1357_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1357_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1357_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1358_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1358_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1358_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1358_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1358_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1358_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1359_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1359_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1359_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1359_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1359_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1359_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1360_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1360_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1360_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1360_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1360_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1360_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1361_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1361_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1361_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1361_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1361_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1361_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1362_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1362_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1362_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1362_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1362_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1362_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1363_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1363_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1363_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1363_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1363_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1363_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1364_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1364_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1364_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1364_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1364_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1364_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1365_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1365_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1365_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1365_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1365_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1365_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1366_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1366_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1366_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1366_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1366_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1366_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1367_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1367_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1367_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1367_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1367_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1367_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1368_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1368_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1368_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1368_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1368_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1368_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1369_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1369_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1369_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1369_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1369_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1369_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1370_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1370_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1370_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1370_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1370_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1370_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1371_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1371_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1371_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1371_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1371_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1371_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1372_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1372_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1372_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1372_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1372_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1372_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1373_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1373_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1373_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1373_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1373_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1373_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1374_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1374_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1374_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1374_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1374_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1374_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1375_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1375_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1375_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1375_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1375_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1375_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1376_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1376_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1376_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1376_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1376_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1376_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1377_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1377_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1377_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1377_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1377_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1377_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1378_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1378_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1378_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1378_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1378_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1378_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1379_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1379_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1379_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1379_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1379_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1379_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1380_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1380_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1380_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1380_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1380_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1380_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1381_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1381_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1381_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1381_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1381_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1381_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1382_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1382_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1382_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1382_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1382_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1382_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1383_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1383_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1383_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1383_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1383_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1383_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1384_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1384_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1384_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1384_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1384_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1384_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1385_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1385_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1385_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1385_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1385_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1385_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1386_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1386_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1386_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1386_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1386_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1386_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1387_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1387_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1387_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1387_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1387_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1387_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1388_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1388_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1388_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1388_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1388_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1388_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1389_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1389_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1389_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1389_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1389_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1389_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1390_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1390_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1390_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1390_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1390_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1390_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1391_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1391_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1391_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1391_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1391_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1391_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1392_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1392_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1392_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1392_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1392_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1392_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1393_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1393_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1393_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1393_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1393_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1393_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1394_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1394_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1394_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1394_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1394_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1394_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1395_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1395_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1395_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1395_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1395_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1395_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1396_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1396_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1396_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1396_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1396_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1396_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1397_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1397_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1397_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1397_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1397_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1397_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1398_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1398_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1398_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1398_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1398_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1398_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1399_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1399_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1399_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1399_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1399_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1399_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1400_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1400_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1400_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1400_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1400_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1400_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1401_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1401_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1401_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1401_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1401_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1401_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1402_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1402_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1402_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1402_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1402_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1402_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1403_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1403_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1403_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1403_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1403_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1403_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1404_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1404_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1404_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1404_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1404_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1404_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1405_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1405_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1405_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1405_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1405_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1405_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1406_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1406_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1406_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1406_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1406_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1406_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1407_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1407_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1407_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1407_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1407_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1407_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1408_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1408_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1408_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1408_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1408_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1408_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1409_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1409_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1409_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1409_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1409_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1409_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1410_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1410_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1410_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1411_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1411_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1411_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1411_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1411_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1411_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1411_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1411_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1411_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1411_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1411_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1411_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1411_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1411_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1411_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1412_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1412_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1412_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1412_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1412_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1412_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1412_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1412_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1412_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1412_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1412_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1412_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1412_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1412_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1412_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1413_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1413_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1413_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1413_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1413_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1413_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1413_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1413_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1413_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1413_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1413_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1413_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1413_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1413_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1413_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1414_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1414_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1414_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1414_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1414_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1414_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1414_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1414_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1414_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1414_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1414_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1414_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1414_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1414_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1414_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1415_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1415_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1415_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1415_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1415_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1415_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1415_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1415_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1415_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1415_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1415_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1415_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1415_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1415_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1415_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1416_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1416_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1416_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1416_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1416_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1416_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1416_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1416_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1416_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1416_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1416_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1416_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1416_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1416_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1416_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1417_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1417_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1417_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1417_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1417_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1417_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1417_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1417_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1417_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1417_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1417_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1417_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1417_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1417_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1417_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1418_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1418_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1418_1366 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1418_1380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2268 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1418_2290 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1418_2304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1418_3214 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1418_3228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4116 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1418_4138 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1418_4152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1418_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1418_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_5964 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1418_5986 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1418_6000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1418_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_882 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1419_904 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1419_918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1146 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1168 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1190 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1278 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1300 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1322 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1806 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1419_1828 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1419_1842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1960 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_1982 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2004 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2026 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2048 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2070 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2092 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2730 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1419_2752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1419_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2884 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2906 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2928 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2950 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2972 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_2994 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3016 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3038 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3060 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3082 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3104 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3126 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3148 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3654 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1419_3676 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1419_3690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3808 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3830 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3852 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3874 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3896 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3918 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3940 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3962 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_3984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4578 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1419_4600 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1419_4614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5216 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1419_5524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1419_5538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_5986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1419_6448 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1419_6462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1419_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_332 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1420_354 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_391 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_461 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_471 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_496 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_506 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_526 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_537 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_550 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_575 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_597 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_641 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_663 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_685 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_707 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_729 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_751 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_773 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_795 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_817 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_839 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_861 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_883 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_905 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_927 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_949 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_971 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_993 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1015 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1037 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1059 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1081 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1103 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1125 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1147 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_1169 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_1175 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_1200 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_1206 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_1215 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_1230 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_1239 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_1250 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_1256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_1258 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1420_1264 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_1278 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_1285 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1420_1304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_1318 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_1324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_1328 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_1334 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_1359 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_1365 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_1379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_1385 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1432 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1718 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1740 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1762 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1784 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1806 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1828 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1938 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_1960 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_1982 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_1984 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_1990 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_2006 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_2021 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2031 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2033 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2039 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_2056 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_2065 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2075 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_2086 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_2095 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2105 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2111 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2118 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2120 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_2126 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2130 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_2136 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2142 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2144 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2150 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_2161 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2167 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2169 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2175 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2197 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2219 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2241 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2263 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2285 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2309 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2752 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2774 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2790 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_2806 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_2821 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2827 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_2833 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2839 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_2846 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2850 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_2856 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2870 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1420_2886 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2900 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2911 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2918 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2920 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_2926 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_2930 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2936 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_2943 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_2949 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_2966 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2975 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_2997 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3019 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3041 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3063 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3085 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3107 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3129 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3151 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3173 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3195 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1420_3217 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_3231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3233 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3566 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_3588 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3598 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_3609 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3613 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_3619 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3623 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_3634 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_3643 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3653 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_3659 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3678 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_3689 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_3714 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_3721 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3728 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_3734 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_3744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_3763 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_3769 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3771 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3777 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_3783 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_3787 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3793 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3815 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3837 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3859 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3881 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3903 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3925 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3947 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3969 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_3991 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4013 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4035 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4057 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4079 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4123 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_4145 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_4155 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_4157 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4358 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_4380 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_4390 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_4392 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_4398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_4423 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_4429 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_4435 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_4437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_4443 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_4454 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_4460 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_4477 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_4488 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_4502 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1420_4513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_4527 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_4538 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_4552 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_4563 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_4569 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_4571 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4604 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4626 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4648 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4670 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4692 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4714 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4736 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4758 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4780 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4802 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4824 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4846 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4868 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4890 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4912 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4934 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4956 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_4978 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5000 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5022 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5044 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1420_5066 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_5080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5172 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_5194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5201 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_5238 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_5249 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_5256 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_5262 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1420_5269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_5288 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_5304 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_5318 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_5329 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_5354 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_5369 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_5373 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_5384 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5393 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5415 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5437 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5459 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5481 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5503 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5525 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5569 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5591 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5613 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5635 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5657 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5679 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5701 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5723 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5745 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5767 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5789 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5811 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5833 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5855 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5877 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5899 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5921 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5943 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_5965 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_5987 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_5999 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_6005 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1420_6008 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_6022 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_6024 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_6035 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_6041 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_6043 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_6049 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_6059 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_6066 ();
 FILLER_ASAP7_75t_R FILLER_0_1420_6072 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_6079 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_6090 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_6099 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_6120 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_6129 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1420_6145 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1420_6154 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_6168 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1420_6179 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6195 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6283 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6327 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6349 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6371 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6393 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6415 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6437 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6459 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6481 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6503 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1420_6525 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1420_6547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1420_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_332 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_354 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_362 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_368 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_376 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_382 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_394 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_410 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_421 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_433 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_439 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_452 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_458 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_475 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_487 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_493 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_500 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_509 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_516 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_552 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_563 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_577 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_584 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_606 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_672 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_694 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_716 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_738 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_760 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_782 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_804 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_826 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_848 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_870 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_892 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_914 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1124 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1421_1146 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_1160 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_1171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_1178 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_1184 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_1194 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_1196 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_1202 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_1213 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_1220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_1227 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_1233 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_1239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_1241 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_1257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_1263 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_1279 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_1285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_1287 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_1293 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_1299 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_1311 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_1318 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_1329 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1344 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_1366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_1376 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_1382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_1384 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1742 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1764 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1786 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1808 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1421_1830 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_1844 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_1938 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_1960 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_1966 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_1973 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_1989 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_1998 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2004 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_2010 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2016 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2022 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2028 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_2044 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2053 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_2059 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2065 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_2076 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_2083 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_2092 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2096 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2107 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_2113 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_2119 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2121 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2127 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_2133 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2137 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_2143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_2158 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_2172 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2338 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2558 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2580 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2602 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2624 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2646 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2668 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2712 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2734 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_2756 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2774 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_2796 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2798 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2804 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_2810 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2822 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_2828 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_2839 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2841 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_2847 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_2854 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2858 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1421_2864 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_2883 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_2895 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_2904 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_2915 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2922 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2933 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_2939 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_2941 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_2984 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3006 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3028 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3050 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3072 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3094 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3534 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_3556 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_3568 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_3584 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_3588 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_3599 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_3605 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_3611 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_3617 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_3621 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_3627 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3633 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_3640 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3646 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_3648 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_3664 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3674 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_3681 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3703 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_3710 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3719 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3726 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_3728 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3734 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3746 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3753 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3760 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_3762 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_3773 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_3779 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_3785 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3792 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3814 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3836 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3858 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3880 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3902 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3924 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3946 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3968 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_3990 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4012 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4034 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4056 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4078 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4122 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4144 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4166 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4188 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4210 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4276 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4298 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_4364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_4368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_4379 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_4395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_4399 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_4415 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_4426 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_4428 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1421_4439 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_4453 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_4459 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_4470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_4472 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_4478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_4488 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_4494 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_4500 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_4507 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_4542 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_4544 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_4550 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_4569 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_4573 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_4584 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5150 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5172 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5183 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_5204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5208 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_5224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5226 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_5232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5236 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_5242 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5246 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_5252 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5254 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_5265 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_5284 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5296 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_5312 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_5321 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_5331 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_5338 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_5345 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_5354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5366 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_5388 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5396 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5418 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5440 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5484 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5506 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1421_5528 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_5542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_5942 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_5964 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_5970 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_5972 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_5978 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_5984 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_5996 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_6006 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_6012 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_6014 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_6025 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_6031 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_6037 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_6044 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_6050 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_6056 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_6067 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_6081 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_6093 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_6099 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1421_6114 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_6124 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1421_6131 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_6135 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_6141 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1421_6148 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1421_6154 ();
 FILLER_ASAP7_75t_R FILLER_0_1421_6170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1421_6536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_332 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1422_354 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_388 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_407 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_415 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_421 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_441 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_456 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_464 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_480 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_497 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_521 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_534 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_545 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_553 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_559 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_575 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_816 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_860 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_882 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_904 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1124 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_1168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1170 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1181 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1187 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1193 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_1199 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_1241 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1253 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_1259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1283 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_1289 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_1301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1393 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1415 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1437 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1459 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1481 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1503 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1525 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1569 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1591 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1613 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1635 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1657 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1679 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1701 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1723 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1745 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1767 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1789 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1811 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1833 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1855 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1877 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1899 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1921 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_1943 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_1965 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1422_1991 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1422_2031 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_2046 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2050 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2061 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2067 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2073 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2080 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2082 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2088 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2090 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2096 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2098 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2104 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2110 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2116 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2118 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2124 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2126 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2137 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2139 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2155 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_2166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2170 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2196 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2218 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2240 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2284 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_2306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_2752 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2758 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2760 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2791 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2793 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_2799 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2805 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_2816 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2820 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_2841 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2845 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2861 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2867 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2873 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_2880 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2889 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2891 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2907 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2909 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1422_2915 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2925 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_2937 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_2951 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2953 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2969 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_2975 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_2996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3194 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1422_3216 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_3230 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3522 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1422_3544 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_3558 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3560 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_3571 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3575 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3596 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3607 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_3618 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_3630 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_3642 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_3654 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3663 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3679 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3690 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_3696 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3702 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3708 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_3714 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_3725 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_3732 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_3748 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3752 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_3758 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_3765 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_3781 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3942 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3964 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_3986 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4008 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4030 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4052 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4074 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4096 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4118 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1422_4140 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_4154 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4336 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_4358 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4375 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4392 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_4398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4400 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_4411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4413 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_4419 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4425 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_4436 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4438 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_4444 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4446 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_4452 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_4501 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4503 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_4519 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_4528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4530 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1422_4546 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4556 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_4567 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_4574 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_4580 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4594 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4638 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4704 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4726 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4748 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4770 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4792 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4814 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4836 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4858 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4880 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4902 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4924 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4946 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4968 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_4990 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5012 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5034 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5056 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_5078 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5128 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1422_5150 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5162 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5173 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5184 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_5196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5200 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5211 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1422_5223 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5253 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5259 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5265 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_5282 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5286 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5292 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5294 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1422_5300 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5332 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5343 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5355 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5362 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5368 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5375 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5397 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5419 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5441 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5463 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5485 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5507 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5529 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5551 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5573 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5595 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5617 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5639 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5661 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5683 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5705 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5727 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5749 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5771 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5793 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5815 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5837 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5859 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5881 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5903 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_5925 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1422_5947 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_5961 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_5963 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_6004 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_6048 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_6057 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_6059 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_6065 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_6071 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_6083 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_6089 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1422_6096 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_6102 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_6108 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_6130 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_6132 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_6148 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_6154 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1422_6168 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_6172 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6193 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6215 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6237 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6259 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6325 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6347 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6369 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6391 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6413 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6435 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6457 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6479 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6501 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1422_6523 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1422_6545 ();
 FILLER_ASAP7_75t_R FILLER_0_1422_6555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1422_6557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_332 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1423_354 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_360 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_382 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_432 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_443 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_450 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_464 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_471 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_510 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_516 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_541 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_547 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1423_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_730 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_774 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_796 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_818 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_840 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_862 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_884 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1423_906 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_926 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_948 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_970 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_992 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1014 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1036 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1058 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1080 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1102 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1124 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1423_1146 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_1160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_1162 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_1173 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_1175 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_1196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_1200 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_1206 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_1212 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_1228 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_1234 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_1236 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_1247 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_1254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1728 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1750 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1772 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1794 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1816 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1423_1838 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1850 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1872 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1894 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1916 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_1938 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_1960 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_1962 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_1988 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_1994 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_2000 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_2007 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_2038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_2044 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_2050 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_2057 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2198 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2220 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2242 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2264 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2286 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_2308 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2378 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2730 ();
 DECAPx4_ASAP7_75t_R FILLER_0_1423_2752 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_2774 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_2838 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_2844 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_2850 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_2852 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_2928 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_2934 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_2940 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_2946 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_2998 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3020 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3042 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3064 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3086 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3108 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3130 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3152 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3174 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3196 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1423_3218 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_3232 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3544 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_3606 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_3613 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_3620 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_3629 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_3661 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_3680 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_3684 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_3690 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_3753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_3764 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_3775 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_3791 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_3996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4040 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4062 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4128 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1423_4150 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_4156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4226 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4248 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4270 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4292 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4336 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1423_4358 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_4364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4392 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_4413 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4422 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_4468 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4476 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_4492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4496 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_4527 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4540 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_4566 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_4578 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4582 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_4593 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4595 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1423_4601 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_4615 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_4619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4732 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4776 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4798 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4820 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4842 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4864 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4886 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4908 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4930 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4952 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4974 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_4996 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5018 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5040 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1423_5062 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1423_5076 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5084 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5128 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1423_5150 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_5164 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5166 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5177 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5223 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_5259 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5329 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_5350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5352 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_5363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5385 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5391 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5397 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5419 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5441 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5463 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5485 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5507 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1423_5529 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5722 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5766 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5788 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5810 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5832 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5854 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5876 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5898 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5920 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_5942 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_5964 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_5966 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_6002 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_6038 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_6054 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_6080 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_6186 ();
 FILLER_ASAP7_75t_R FILLER_0_1423_6192 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6199 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6221 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6243 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6265 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6287 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6309 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6331 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6353 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6375 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6397 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6419 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6441 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1423_6463 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1423_6467 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1423_6536 ();
endmodule
