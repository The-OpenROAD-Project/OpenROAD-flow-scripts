VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_256x95
  FOREIGN fakeram45_256x95 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 115.140 BY 119.000 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.365 0.070 1.435 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.645 0.070 1.715 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.925 0.070 1.995 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.205 0.070 2.275 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.485 0.070 2.555 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.765 0.070 2.835 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.045 0.070 3.115 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.325 0.070 3.395 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.605 0.070 3.675 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.885 0.070 3.955 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.165 0.070 4.235 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.445 0.070 4.515 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.725 0.070 4.795 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.005 0.070 5.075 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.285 0.070 5.355 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.565 0.070 5.635 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.845 0.070 5.915 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.125 0.070 6.195 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.405 0.070 6.475 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.685 0.070 6.755 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.965 0.070 7.035 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.245 0.070 7.315 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.525 0.070 7.595 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.805 0.070 7.875 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.085 0.070 8.155 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.365 0.070 8.435 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.645 0.070 8.715 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.925 0.070 8.995 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.205 0.070 9.275 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.485 0.070 9.555 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.765 0.070 9.835 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.045 0.070 10.115 ;
    END
  END w_mask_in[31]
  PIN w_mask_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.325 0.070 10.395 ;
    END
  END w_mask_in[32]
  PIN w_mask_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.605 0.070 10.675 ;
    END
  END w_mask_in[33]
  PIN w_mask_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.885 0.070 10.955 ;
    END
  END w_mask_in[34]
  PIN w_mask_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.165 0.070 11.235 ;
    END
  END w_mask_in[35]
  PIN w_mask_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.445 0.070 11.515 ;
    END
  END w_mask_in[36]
  PIN w_mask_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.725 0.070 11.795 ;
    END
  END w_mask_in[37]
  PIN w_mask_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.005 0.070 12.075 ;
    END
  END w_mask_in[38]
  PIN w_mask_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.285 0.070 12.355 ;
    END
  END w_mask_in[39]
  PIN w_mask_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.565 0.070 12.635 ;
    END
  END w_mask_in[40]
  PIN w_mask_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.845 0.070 12.915 ;
    END
  END w_mask_in[41]
  PIN w_mask_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.125 0.070 13.195 ;
    END
  END w_mask_in[42]
  PIN w_mask_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.405 0.070 13.475 ;
    END
  END w_mask_in[43]
  PIN w_mask_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.685 0.070 13.755 ;
    END
  END w_mask_in[44]
  PIN w_mask_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.965 0.070 14.035 ;
    END
  END w_mask_in[45]
  PIN w_mask_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.245 0.070 14.315 ;
    END
  END w_mask_in[46]
  PIN w_mask_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.525 0.070 14.595 ;
    END
  END w_mask_in[47]
  PIN w_mask_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.805 0.070 14.875 ;
    END
  END w_mask_in[48]
  PIN w_mask_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.085 0.070 15.155 ;
    END
  END w_mask_in[49]
  PIN w_mask_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.365 0.070 15.435 ;
    END
  END w_mask_in[50]
  PIN w_mask_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.645 0.070 15.715 ;
    END
  END w_mask_in[51]
  PIN w_mask_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.925 0.070 15.995 ;
    END
  END w_mask_in[52]
  PIN w_mask_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.205 0.070 16.275 ;
    END
  END w_mask_in[53]
  PIN w_mask_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.485 0.070 16.555 ;
    END
  END w_mask_in[54]
  PIN w_mask_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.765 0.070 16.835 ;
    END
  END w_mask_in[55]
  PIN w_mask_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.045 0.070 17.115 ;
    END
  END w_mask_in[56]
  PIN w_mask_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.325 0.070 17.395 ;
    END
  END w_mask_in[57]
  PIN w_mask_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.605 0.070 17.675 ;
    END
  END w_mask_in[58]
  PIN w_mask_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.885 0.070 17.955 ;
    END
  END w_mask_in[59]
  PIN w_mask_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.165 0.070 18.235 ;
    END
  END w_mask_in[60]
  PIN w_mask_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.445 0.070 18.515 ;
    END
  END w_mask_in[61]
  PIN w_mask_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.725 0.070 18.795 ;
    END
  END w_mask_in[62]
  PIN w_mask_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.005 0.070 19.075 ;
    END
  END w_mask_in[63]
  PIN w_mask_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.285 0.070 19.355 ;
    END
  END w_mask_in[64]
  PIN w_mask_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.565 0.070 19.635 ;
    END
  END w_mask_in[65]
  PIN w_mask_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.845 0.070 19.915 ;
    END
  END w_mask_in[66]
  PIN w_mask_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.125 0.070 20.195 ;
    END
  END w_mask_in[67]
  PIN w_mask_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.405 0.070 20.475 ;
    END
  END w_mask_in[68]
  PIN w_mask_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.685 0.070 20.755 ;
    END
  END w_mask_in[69]
  PIN w_mask_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.965 0.070 21.035 ;
    END
  END w_mask_in[70]
  PIN w_mask_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.245 0.070 21.315 ;
    END
  END w_mask_in[71]
  PIN w_mask_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.525 0.070 21.595 ;
    END
  END w_mask_in[72]
  PIN w_mask_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.805 0.070 21.875 ;
    END
  END w_mask_in[73]
  PIN w_mask_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.085 0.070 22.155 ;
    END
  END w_mask_in[74]
  PIN w_mask_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.365 0.070 22.435 ;
    END
  END w_mask_in[75]
  PIN w_mask_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.645 0.070 22.715 ;
    END
  END w_mask_in[76]
  PIN w_mask_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.925 0.070 22.995 ;
    END
  END w_mask_in[77]
  PIN w_mask_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.205 0.070 23.275 ;
    END
  END w_mask_in[78]
  PIN w_mask_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.485 0.070 23.555 ;
    END
  END w_mask_in[79]
  PIN w_mask_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.765 0.070 23.835 ;
    END
  END w_mask_in[80]
  PIN w_mask_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.045 0.070 24.115 ;
    END
  END w_mask_in[81]
  PIN w_mask_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.325 0.070 24.395 ;
    END
  END w_mask_in[82]
  PIN w_mask_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.605 0.070 24.675 ;
    END
  END w_mask_in[83]
  PIN w_mask_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.885 0.070 24.955 ;
    END
  END w_mask_in[84]
  PIN w_mask_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.165 0.070 25.235 ;
    END
  END w_mask_in[85]
  PIN w_mask_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.445 0.070 25.515 ;
    END
  END w_mask_in[86]
  PIN w_mask_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.725 0.070 25.795 ;
    END
  END w_mask_in[87]
  PIN w_mask_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.005 0.070 26.075 ;
    END
  END w_mask_in[88]
  PIN w_mask_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.285 0.070 26.355 ;
    END
  END w_mask_in[89]
  PIN w_mask_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.565 0.070 26.635 ;
    END
  END w_mask_in[90]
  PIN w_mask_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.845 0.070 26.915 ;
    END
  END w_mask_in[91]
  PIN w_mask_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.125 0.070 27.195 ;
    END
  END w_mask_in[92]
  PIN w_mask_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.405 0.070 27.475 ;
    END
  END w_mask_in[93]
  PIN w_mask_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.685 0.070 27.755 ;
    END
  END w_mask_in[94]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.945 0.070 36.015 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.225 0.070 36.295 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.505 0.070 36.575 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.785 0.070 36.855 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.065 0.070 37.135 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.345 0.070 37.415 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.625 0.070 37.695 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.905 0.070 37.975 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.185 0.070 38.255 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.465 0.070 38.535 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.745 0.070 38.815 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.025 0.070 39.095 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.305 0.070 39.375 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.585 0.070 39.655 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.865 0.070 39.935 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.145 0.070 40.215 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.425 0.070 40.495 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.705 0.070 40.775 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.985 0.070 41.055 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.265 0.070 41.335 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.545 0.070 41.615 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.825 0.070 41.895 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.105 0.070 42.175 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.385 0.070 42.455 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.665 0.070 42.735 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.945 0.070 43.015 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.225 0.070 43.295 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.505 0.070 43.575 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.785 0.070 43.855 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.065 0.070 44.135 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.345 0.070 44.415 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.625 0.070 44.695 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.905 0.070 44.975 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.185 0.070 45.255 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.465 0.070 45.535 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.745 0.070 45.815 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.025 0.070 46.095 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.305 0.070 46.375 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.585 0.070 46.655 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.865 0.070 46.935 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.145 0.070 47.215 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.425 0.070 47.495 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.705 0.070 47.775 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.985 0.070 48.055 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.265 0.070 48.335 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.545 0.070 48.615 ;
    END
  END rd_out[45]
  PIN rd_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.825 0.070 48.895 ;
    END
  END rd_out[46]
  PIN rd_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.105 0.070 49.175 ;
    END
  END rd_out[47]
  PIN rd_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.385 0.070 49.455 ;
    END
  END rd_out[48]
  PIN rd_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.665 0.070 49.735 ;
    END
  END rd_out[49]
  PIN rd_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.945 0.070 50.015 ;
    END
  END rd_out[50]
  PIN rd_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.225 0.070 50.295 ;
    END
  END rd_out[51]
  PIN rd_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.505 0.070 50.575 ;
    END
  END rd_out[52]
  PIN rd_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.785 0.070 50.855 ;
    END
  END rd_out[53]
  PIN rd_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.065 0.070 51.135 ;
    END
  END rd_out[54]
  PIN rd_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.345 0.070 51.415 ;
    END
  END rd_out[55]
  PIN rd_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.625 0.070 51.695 ;
    END
  END rd_out[56]
  PIN rd_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.905 0.070 51.975 ;
    END
  END rd_out[57]
  PIN rd_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.185 0.070 52.255 ;
    END
  END rd_out[58]
  PIN rd_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.465 0.070 52.535 ;
    END
  END rd_out[59]
  PIN rd_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.745 0.070 52.815 ;
    END
  END rd_out[60]
  PIN rd_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.025 0.070 53.095 ;
    END
  END rd_out[61]
  PIN rd_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.305 0.070 53.375 ;
    END
  END rd_out[62]
  PIN rd_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.585 0.070 53.655 ;
    END
  END rd_out[63]
  PIN rd_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.865 0.070 53.935 ;
    END
  END rd_out[64]
  PIN rd_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.145 0.070 54.215 ;
    END
  END rd_out[65]
  PIN rd_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.425 0.070 54.495 ;
    END
  END rd_out[66]
  PIN rd_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.705 0.070 54.775 ;
    END
  END rd_out[67]
  PIN rd_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.985 0.070 55.055 ;
    END
  END rd_out[68]
  PIN rd_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.265 0.070 55.335 ;
    END
  END rd_out[69]
  PIN rd_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.545 0.070 55.615 ;
    END
  END rd_out[70]
  PIN rd_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.825 0.070 55.895 ;
    END
  END rd_out[71]
  PIN rd_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.105 0.070 56.175 ;
    END
  END rd_out[72]
  PIN rd_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.385 0.070 56.455 ;
    END
  END rd_out[73]
  PIN rd_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.665 0.070 56.735 ;
    END
  END rd_out[74]
  PIN rd_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.945 0.070 57.015 ;
    END
  END rd_out[75]
  PIN rd_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.225 0.070 57.295 ;
    END
  END rd_out[76]
  PIN rd_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.505 0.070 57.575 ;
    END
  END rd_out[77]
  PIN rd_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.785 0.070 57.855 ;
    END
  END rd_out[78]
  PIN rd_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.065 0.070 58.135 ;
    END
  END rd_out[79]
  PIN rd_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.345 0.070 58.415 ;
    END
  END rd_out[80]
  PIN rd_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.625 0.070 58.695 ;
    END
  END rd_out[81]
  PIN rd_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.905 0.070 58.975 ;
    END
  END rd_out[82]
  PIN rd_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.185 0.070 59.255 ;
    END
  END rd_out[83]
  PIN rd_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.465 0.070 59.535 ;
    END
  END rd_out[84]
  PIN rd_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.745 0.070 59.815 ;
    END
  END rd_out[85]
  PIN rd_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.025 0.070 60.095 ;
    END
  END rd_out[86]
  PIN rd_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.305 0.070 60.375 ;
    END
  END rd_out[87]
  PIN rd_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.585 0.070 60.655 ;
    END
  END rd_out[88]
  PIN rd_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.865 0.070 60.935 ;
    END
  END rd_out[89]
  PIN rd_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.145 0.070 61.215 ;
    END
  END rd_out[90]
  PIN rd_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.425 0.070 61.495 ;
    END
  END rd_out[91]
  PIN rd_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.705 0.070 61.775 ;
    END
  END rd_out[92]
  PIN rd_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 61.985 0.070 62.055 ;
    END
  END rd_out[93]
  PIN rd_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 62.265 0.070 62.335 ;
    END
  END rd_out[94]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.525 0.070 70.595 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 70.805 0.070 70.875 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.085 0.070 71.155 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.365 0.070 71.435 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.645 0.070 71.715 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 71.925 0.070 71.995 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.205 0.070 72.275 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.485 0.070 72.555 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 72.765 0.070 72.835 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.045 0.070 73.115 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.325 0.070 73.395 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.605 0.070 73.675 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 73.885 0.070 73.955 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.165 0.070 74.235 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.445 0.070 74.515 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 74.725 0.070 74.795 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.005 0.070 75.075 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.285 0.070 75.355 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.565 0.070 75.635 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 75.845 0.070 75.915 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.125 0.070 76.195 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.405 0.070 76.475 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.685 0.070 76.755 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 76.965 0.070 77.035 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.245 0.070 77.315 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.525 0.070 77.595 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 77.805 0.070 77.875 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.085 0.070 78.155 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.365 0.070 78.435 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.645 0.070 78.715 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 78.925 0.070 78.995 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.205 0.070 79.275 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.485 0.070 79.555 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 79.765 0.070 79.835 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.045 0.070 80.115 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.325 0.070 80.395 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.605 0.070 80.675 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 80.885 0.070 80.955 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.165 0.070 81.235 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.445 0.070 81.515 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 81.725 0.070 81.795 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.005 0.070 82.075 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.285 0.070 82.355 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.565 0.070 82.635 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 82.845 0.070 82.915 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.125 0.070 83.195 ;
    END
  END wd_in[45]
  PIN wd_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.405 0.070 83.475 ;
    END
  END wd_in[46]
  PIN wd_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.685 0.070 83.755 ;
    END
  END wd_in[47]
  PIN wd_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 83.965 0.070 84.035 ;
    END
  END wd_in[48]
  PIN wd_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.245 0.070 84.315 ;
    END
  END wd_in[49]
  PIN wd_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.525 0.070 84.595 ;
    END
  END wd_in[50]
  PIN wd_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 84.805 0.070 84.875 ;
    END
  END wd_in[51]
  PIN wd_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.085 0.070 85.155 ;
    END
  END wd_in[52]
  PIN wd_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.365 0.070 85.435 ;
    END
  END wd_in[53]
  PIN wd_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.645 0.070 85.715 ;
    END
  END wd_in[54]
  PIN wd_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 85.925 0.070 85.995 ;
    END
  END wd_in[55]
  PIN wd_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.205 0.070 86.275 ;
    END
  END wd_in[56]
  PIN wd_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.485 0.070 86.555 ;
    END
  END wd_in[57]
  PIN wd_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 86.765 0.070 86.835 ;
    END
  END wd_in[58]
  PIN wd_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.045 0.070 87.115 ;
    END
  END wd_in[59]
  PIN wd_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.325 0.070 87.395 ;
    END
  END wd_in[60]
  PIN wd_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.605 0.070 87.675 ;
    END
  END wd_in[61]
  PIN wd_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 87.885 0.070 87.955 ;
    END
  END wd_in[62]
  PIN wd_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.165 0.070 88.235 ;
    END
  END wd_in[63]
  PIN wd_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.445 0.070 88.515 ;
    END
  END wd_in[64]
  PIN wd_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 88.725 0.070 88.795 ;
    END
  END wd_in[65]
  PIN wd_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.005 0.070 89.075 ;
    END
  END wd_in[66]
  PIN wd_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.285 0.070 89.355 ;
    END
  END wd_in[67]
  PIN wd_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.565 0.070 89.635 ;
    END
  END wd_in[68]
  PIN wd_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 89.845 0.070 89.915 ;
    END
  END wd_in[69]
  PIN wd_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.125 0.070 90.195 ;
    END
  END wd_in[70]
  PIN wd_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.405 0.070 90.475 ;
    END
  END wd_in[71]
  PIN wd_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.685 0.070 90.755 ;
    END
  END wd_in[72]
  PIN wd_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 90.965 0.070 91.035 ;
    END
  END wd_in[73]
  PIN wd_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.245 0.070 91.315 ;
    END
  END wd_in[74]
  PIN wd_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.525 0.070 91.595 ;
    END
  END wd_in[75]
  PIN wd_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 91.805 0.070 91.875 ;
    END
  END wd_in[76]
  PIN wd_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.085 0.070 92.155 ;
    END
  END wd_in[77]
  PIN wd_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.365 0.070 92.435 ;
    END
  END wd_in[78]
  PIN wd_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.645 0.070 92.715 ;
    END
  END wd_in[79]
  PIN wd_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 92.925 0.070 92.995 ;
    END
  END wd_in[80]
  PIN wd_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.205 0.070 93.275 ;
    END
  END wd_in[81]
  PIN wd_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.485 0.070 93.555 ;
    END
  END wd_in[82]
  PIN wd_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 93.765 0.070 93.835 ;
    END
  END wd_in[83]
  PIN wd_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.045 0.070 94.115 ;
    END
  END wd_in[84]
  PIN wd_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.325 0.070 94.395 ;
    END
  END wd_in[85]
  PIN wd_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.605 0.070 94.675 ;
    END
  END wd_in[86]
  PIN wd_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 94.885 0.070 94.955 ;
    END
  END wd_in[87]
  PIN wd_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.165 0.070 95.235 ;
    END
  END wd_in[88]
  PIN wd_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.445 0.070 95.515 ;
    END
  END wd_in[89]
  PIN wd_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 95.725 0.070 95.795 ;
    END
  END wd_in[90]
  PIN wd_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.005 0.070 96.075 ;
    END
  END wd_in[91]
  PIN wd_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.285 0.070 96.355 ;
    END
  END wd_in[92]
  PIN wd_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.565 0.070 96.635 ;
    END
  END wd_in[93]
  PIN wd_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 96.845 0.070 96.915 ;
    END
  END wd_in[94]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.105 0.070 105.175 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.385 0.070 105.455 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.665 0.070 105.735 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 105.945 0.070 106.015 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.225 0.070 106.295 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.505 0.070 106.575 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 106.785 0.070 106.855 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 107.065 0.070 107.135 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.325 0.070 115.395 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.605 0.070 115.675 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 115.885 0.070 115.955 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 117.600 ;
      RECT 3.500 1.400 3.780 117.600 ;
      RECT 5.740 1.400 6.020 117.600 ;
      RECT 7.980 1.400 8.260 117.600 ;
      RECT 10.220 1.400 10.500 117.600 ;
      RECT 12.460 1.400 12.740 117.600 ;
      RECT 14.700 1.400 14.980 117.600 ;
      RECT 16.940 1.400 17.220 117.600 ;
      RECT 19.180 1.400 19.460 117.600 ;
      RECT 21.420 1.400 21.700 117.600 ;
      RECT 23.660 1.400 23.940 117.600 ;
      RECT 25.900 1.400 26.180 117.600 ;
      RECT 28.140 1.400 28.420 117.600 ;
      RECT 30.380 1.400 30.660 117.600 ;
      RECT 32.620 1.400 32.900 117.600 ;
      RECT 34.860 1.400 35.140 117.600 ;
      RECT 37.100 1.400 37.380 117.600 ;
      RECT 39.340 1.400 39.620 117.600 ;
      RECT 41.580 1.400 41.860 117.600 ;
      RECT 43.820 1.400 44.100 117.600 ;
      RECT 46.060 1.400 46.340 117.600 ;
      RECT 48.300 1.400 48.580 117.600 ;
      RECT 50.540 1.400 50.820 117.600 ;
      RECT 52.780 1.400 53.060 117.600 ;
      RECT 55.020 1.400 55.300 117.600 ;
      RECT 57.260 1.400 57.540 117.600 ;
      RECT 59.500 1.400 59.780 117.600 ;
      RECT 61.740 1.400 62.020 117.600 ;
      RECT 63.980 1.400 64.260 117.600 ;
      RECT 66.220 1.400 66.500 117.600 ;
      RECT 68.460 1.400 68.740 117.600 ;
      RECT 70.700 1.400 70.980 117.600 ;
      RECT 72.940 1.400 73.220 117.600 ;
      RECT 75.180 1.400 75.460 117.600 ;
      RECT 77.420 1.400 77.700 117.600 ;
      RECT 79.660 1.400 79.940 117.600 ;
      RECT 81.900 1.400 82.180 117.600 ;
      RECT 84.140 1.400 84.420 117.600 ;
      RECT 86.380 1.400 86.660 117.600 ;
      RECT 88.620 1.400 88.900 117.600 ;
      RECT 90.860 1.400 91.140 117.600 ;
      RECT 93.100 1.400 93.380 117.600 ;
      RECT 95.340 1.400 95.620 117.600 ;
      RECT 97.580 1.400 97.860 117.600 ;
      RECT 99.820 1.400 100.100 117.600 ;
      RECT 102.060 1.400 102.340 117.600 ;
      RECT 104.300 1.400 104.580 117.600 ;
      RECT 106.540 1.400 106.820 117.600 ;
      RECT 108.780 1.400 109.060 117.600 ;
      RECT 111.020 1.400 111.300 117.600 ;
      RECT 113.260 1.400 113.540 117.600 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 117.600 ;
      RECT 4.620 1.400 4.900 117.600 ;
      RECT 6.860 1.400 7.140 117.600 ;
      RECT 9.100 1.400 9.380 117.600 ;
      RECT 11.340 1.400 11.620 117.600 ;
      RECT 13.580 1.400 13.860 117.600 ;
      RECT 15.820 1.400 16.100 117.600 ;
      RECT 18.060 1.400 18.340 117.600 ;
      RECT 20.300 1.400 20.580 117.600 ;
      RECT 22.540 1.400 22.820 117.600 ;
      RECT 24.780 1.400 25.060 117.600 ;
      RECT 27.020 1.400 27.300 117.600 ;
      RECT 29.260 1.400 29.540 117.600 ;
      RECT 31.500 1.400 31.780 117.600 ;
      RECT 33.740 1.400 34.020 117.600 ;
      RECT 35.980 1.400 36.260 117.600 ;
      RECT 38.220 1.400 38.500 117.600 ;
      RECT 40.460 1.400 40.740 117.600 ;
      RECT 42.700 1.400 42.980 117.600 ;
      RECT 44.940 1.400 45.220 117.600 ;
      RECT 47.180 1.400 47.460 117.600 ;
      RECT 49.420 1.400 49.700 117.600 ;
      RECT 51.660 1.400 51.940 117.600 ;
      RECT 53.900 1.400 54.180 117.600 ;
      RECT 56.140 1.400 56.420 117.600 ;
      RECT 58.380 1.400 58.660 117.600 ;
      RECT 60.620 1.400 60.900 117.600 ;
      RECT 62.860 1.400 63.140 117.600 ;
      RECT 65.100 1.400 65.380 117.600 ;
      RECT 67.340 1.400 67.620 117.600 ;
      RECT 69.580 1.400 69.860 117.600 ;
      RECT 71.820 1.400 72.100 117.600 ;
      RECT 74.060 1.400 74.340 117.600 ;
      RECT 76.300 1.400 76.580 117.600 ;
      RECT 78.540 1.400 78.820 117.600 ;
      RECT 80.780 1.400 81.060 117.600 ;
      RECT 83.020 1.400 83.300 117.600 ;
      RECT 85.260 1.400 85.540 117.600 ;
      RECT 87.500 1.400 87.780 117.600 ;
      RECT 89.740 1.400 90.020 117.600 ;
      RECT 91.980 1.400 92.260 117.600 ;
      RECT 94.220 1.400 94.500 117.600 ;
      RECT 96.460 1.400 96.740 117.600 ;
      RECT 98.700 1.400 98.980 117.600 ;
      RECT 100.940 1.400 101.220 117.600 ;
      RECT 103.180 1.400 103.460 117.600 ;
      RECT 105.420 1.400 105.700 117.600 ;
      RECT 107.660 1.400 107.940 117.600 ;
      RECT 109.900 1.400 110.180 117.600 ;
      RECT 112.140 1.400 112.420 117.600 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 115.140 119.000 ;
    LAYER metal2 ;
    RECT 0 0 115.140 119.000 ;
    LAYER metal3 ;
    RECT 0.070 0 115.140 119.000 ;
    RECT 0 0.000 0.070 1.365 ;
    RECT 0 1.435 0.070 1.645 ;
    RECT 0 1.715 0.070 1.925 ;
    RECT 0 1.995 0.070 2.205 ;
    RECT 0 2.275 0.070 2.485 ;
    RECT 0 2.555 0.070 2.765 ;
    RECT 0 2.835 0.070 3.045 ;
    RECT 0 3.115 0.070 3.325 ;
    RECT 0 3.395 0.070 3.605 ;
    RECT 0 3.675 0.070 3.885 ;
    RECT 0 3.955 0.070 4.165 ;
    RECT 0 4.235 0.070 4.445 ;
    RECT 0 4.515 0.070 4.725 ;
    RECT 0 4.795 0.070 5.005 ;
    RECT 0 5.075 0.070 5.285 ;
    RECT 0 5.355 0.070 5.565 ;
    RECT 0 5.635 0.070 5.845 ;
    RECT 0 5.915 0.070 6.125 ;
    RECT 0 6.195 0.070 6.405 ;
    RECT 0 6.475 0.070 6.685 ;
    RECT 0 6.755 0.070 6.965 ;
    RECT 0 7.035 0.070 7.245 ;
    RECT 0 7.315 0.070 7.525 ;
    RECT 0 7.595 0.070 7.805 ;
    RECT 0 7.875 0.070 8.085 ;
    RECT 0 8.155 0.070 8.365 ;
    RECT 0 8.435 0.070 8.645 ;
    RECT 0 8.715 0.070 8.925 ;
    RECT 0 8.995 0.070 9.205 ;
    RECT 0 9.275 0.070 9.485 ;
    RECT 0 9.555 0.070 9.765 ;
    RECT 0 9.835 0.070 10.045 ;
    RECT 0 10.115 0.070 10.325 ;
    RECT 0 10.395 0.070 10.605 ;
    RECT 0 10.675 0.070 10.885 ;
    RECT 0 10.955 0.070 11.165 ;
    RECT 0 11.235 0.070 11.445 ;
    RECT 0 11.515 0.070 11.725 ;
    RECT 0 11.795 0.070 12.005 ;
    RECT 0 12.075 0.070 12.285 ;
    RECT 0 12.355 0.070 12.565 ;
    RECT 0 12.635 0.070 12.845 ;
    RECT 0 12.915 0.070 13.125 ;
    RECT 0 13.195 0.070 13.405 ;
    RECT 0 13.475 0.070 13.685 ;
    RECT 0 13.755 0.070 13.965 ;
    RECT 0 14.035 0.070 14.245 ;
    RECT 0 14.315 0.070 14.525 ;
    RECT 0 14.595 0.070 14.805 ;
    RECT 0 14.875 0.070 15.085 ;
    RECT 0 15.155 0.070 15.365 ;
    RECT 0 15.435 0.070 15.645 ;
    RECT 0 15.715 0.070 15.925 ;
    RECT 0 15.995 0.070 16.205 ;
    RECT 0 16.275 0.070 16.485 ;
    RECT 0 16.555 0.070 16.765 ;
    RECT 0 16.835 0.070 17.045 ;
    RECT 0 17.115 0.070 17.325 ;
    RECT 0 17.395 0.070 17.605 ;
    RECT 0 17.675 0.070 17.885 ;
    RECT 0 17.955 0.070 18.165 ;
    RECT 0 18.235 0.070 18.445 ;
    RECT 0 18.515 0.070 18.725 ;
    RECT 0 18.795 0.070 19.005 ;
    RECT 0 19.075 0.070 19.285 ;
    RECT 0 19.355 0.070 19.565 ;
    RECT 0 19.635 0.070 19.845 ;
    RECT 0 19.915 0.070 20.125 ;
    RECT 0 20.195 0.070 20.405 ;
    RECT 0 20.475 0.070 20.685 ;
    RECT 0 20.755 0.070 20.965 ;
    RECT 0 21.035 0.070 21.245 ;
    RECT 0 21.315 0.070 21.525 ;
    RECT 0 21.595 0.070 21.805 ;
    RECT 0 21.875 0.070 22.085 ;
    RECT 0 22.155 0.070 22.365 ;
    RECT 0 22.435 0.070 22.645 ;
    RECT 0 22.715 0.070 22.925 ;
    RECT 0 22.995 0.070 23.205 ;
    RECT 0 23.275 0.070 23.485 ;
    RECT 0 23.555 0.070 23.765 ;
    RECT 0 23.835 0.070 24.045 ;
    RECT 0 24.115 0.070 24.325 ;
    RECT 0 24.395 0.070 24.605 ;
    RECT 0 24.675 0.070 24.885 ;
    RECT 0 24.955 0.070 25.165 ;
    RECT 0 25.235 0.070 25.445 ;
    RECT 0 25.515 0.070 25.725 ;
    RECT 0 25.795 0.070 26.005 ;
    RECT 0 26.075 0.070 26.285 ;
    RECT 0 26.355 0.070 26.565 ;
    RECT 0 26.635 0.070 26.845 ;
    RECT 0 26.915 0.070 27.125 ;
    RECT 0 27.195 0.070 27.405 ;
    RECT 0 27.475 0.070 27.685 ;
    RECT 0 27.755 0.070 35.945 ;
    RECT 0 36.015 0.070 36.225 ;
    RECT 0 36.295 0.070 36.505 ;
    RECT 0 36.575 0.070 36.785 ;
    RECT 0 36.855 0.070 37.065 ;
    RECT 0 37.135 0.070 37.345 ;
    RECT 0 37.415 0.070 37.625 ;
    RECT 0 37.695 0.070 37.905 ;
    RECT 0 37.975 0.070 38.185 ;
    RECT 0 38.255 0.070 38.465 ;
    RECT 0 38.535 0.070 38.745 ;
    RECT 0 38.815 0.070 39.025 ;
    RECT 0 39.095 0.070 39.305 ;
    RECT 0 39.375 0.070 39.585 ;
    RECT 0 39.655 0.070 39.865 ;
    RECT 0 39.935 0.070 40.145 ;
    RECT 0 40.215 0.070 40.425 ;
    RECT 0 40.495 0.070 40.705 ;
    RECT 0 40.775 0.070 40.985 ;
    RECT 0 41.055 0.070 41.265 ;
    RECT 0 41.335 0.070 41.545 ;
    RECT 0 41.615 0.070 41.825 ;
    RECT 0 41.895 0.070 42.105 ;
    RECT 0 42.175 0.070 42.385 ;
    RECT 0 42.455 0.070 42.665 ;
    RECT 0 42.735 0.070 42.945 ;
    RECT 0 43.015 0.070 43.225 ;
    RECT 0 43.295 0.070 43.505 ;
    RECT 0 43.575 0.070 43.785 ;
    RECT 0 43.855 0.070 44.065 ;
    RECT 0 44.135 0.070 44.345 ;
    RECT 0 44.415 0.070 44.625 ;
    RECT 0 44.695 0.070 44.905 ;
    RECT 0 44.975 0.070 45.185 ;
    RECT 0 45.255 0.070 45.465 ;
    RECT 0 45.535 0.070 45.745 ;
    RECT 0 45.815 0.070 46.025 ;
    RECT 0 46.095 0.070 46.305 ;
    RECT 0 46.375 0.070 46.585 ;
    RECT 0 46.655 0.070 46.865 ;
    RECT 0 46.935 0.070 47.145 ;
    RECT 0 47.215 0.070 47.425 ;
    RECT 0 47.495 0.070 47.705 ;
    RECT 0 47.775 0.070 47.985 ;
    RECT 0 48.055 0.070 48.265 ;
    RECT 0 48.335 0.070 48.545 ;
    RECT 0 48.615 0.070 48.825 ;
    RECT 0 48.895 0.070 49.105 ;
    RECT 0 49.175 0.070 49.385 ;
    RECT 0 49.455 0.070 49.665 ;
    RECT 0 49.735 0.070 49.945 ;
    RECT 0 50.015 0.070 50.225 ;
    RECT 0 50.295 0.070 50.505 ;
    RECT 0 50.575 0.070 50.785 ;
    RECT 0 50.855 0.070 51.065 ;
    RECT 0 51.135 0.070 51.345 ;
    RECT 0 51.415 0.070 51.625 ;
    RECT 0 51.695 0.070 51.905 ;
    RECT 0 51.975 0.070 52.185 ;
    RECT 0 52.255 0.070 52.465 ;
    RECT 0 52.535 0.070 52.745 ;
    RECT 0 52.815 0.070 53.025 ;
    RECT 0 53.095 0.070 53.305 ;
    RECT 0 53.375 0.070 53.585 ;
    RECT 0 53.655 0.070 53.865 ;
    RECT 0 53.935 0.070 54.145 ;
    RECT 0 54.215 0.070 54.425 ;
    RECT 0 54.495 0.070 54.705 ;
    RECT 0 54.775 0.070 54.985 ;
    RECT 0 55.055 0.070 55.265 ;
    RECT 0 55.335 0.070 55.545 ;
    RECT 0 55.615 0.070 55.825 ;
    RECT 0 55.895 0.070 56.105 ;
    RECT 0 56.175 0.070 56.385 ;
    RECT 0 56.455 0.070 56.665 ;
    RECT 0 56.735 0.070 56.945 ;
    RECT 0 57.015 0.070 57.225 ;
    RECT 0 57.295 0.070 57.505 ;
    RECT 0 57.575 0.070 57.785 ;
    RECT 0 57.855 0.070 58.065 ;
    RECT 0 58.135 0.070 58.345 ;
    RECT 0 58.415 0.070 58.625 ;
    RECT 0 58.695 0.070 58.905 ;
    RECT 0 58.975 0.070 59.185 ;
    RECT 0 59.255 0.070 59.465 ;
    RECT 0 59.535 0.070 59.745 ;
    RECT 0 59.815 0.070 60.025 ;
    RECT 0 60.095 0.070 60.305 ;
    RECT 0 60.375 0.070 60.585 ;
    RECT 0 60.655 0.070 60.865 ;
    RECT 0 60.935 0.070 61.145 ;
    RECT 0 61.215 0.070 61.425 ;
    RECT 0 61.495 0.070 61.705 ;
    RECT 0 61.775 0.070 61.985 ;
    RECT 0 62.055 0.070 62.265 ;
    RECT 0 62.335 0.070 70.525 ;
    RECT 0 70.595 0.070 70.805 ;
    RECT 0 70.875 0.070 71.085 ;
    RECT 0 71.155 0.070 71.365 ;
    RECT 0 71.435 0.070 71.645 ;
    RECT 0 71.715 0.070 71.925 ;
    RECT 0 71.995 0.070 72.205 ;
    RECT 0 72.275 0.070 72.485 ;
    RECT 0 72.555 0.070 72.765 ;
    RECT 0 72.835 0.070 73.045 ;
    RECT 0 73.115 0.070 73.325 ;
    RECT 0 73.395 0.070 73.605 ;
    RECT 0 73.675 0.070 73.885 ;
    RECT 0 73.955 0.070 74.165 ;
    RECT 0 74.235 0.070 74.445 ;
    RECT 0 74.515 0.070 74.725 ;
    RECT 0 74.795 0.070 75.005 ;
    RECT 0 75.075 0.070 75.285 ;
    RECT 0 75.355 0.070 75.565 ;
    RECT 0 75.635 0.070 75.845 ;
    RECT 0 75.915 0.070 76.125 ;
    RECT 0 76.195 0.070 76.405 ;
    RECT 0 76.475 0.070 76.685 ;
    RECT 0 76.755 0.070 76.965 ;
    RECT 0 77.035 0.070 77.245 ;
    RECT 0 77.315 0.070 77.525 ;
    RECT 0 77.595 0.070 77.805 ;
    RECT 0 77.875 0.070 78.085 ;
    RECT 0 78.155 0.070 78.365 ;
    RECT 0 78.435 0.070 78.645 ;
    RECT 0 78.715 0.070 78.925 ;
    RECT 0 78.995 0.070 79.205 ;
    RECT 0 79.275 0.070 79.485 ;
    RECT 0 79.555 0.070 79.765 ;
    RECT 0 79.835 0.070 80.045 ;
    RECT 0 80.115 0.070 80.325 ;
    RECT 0 80.395 0.070 80.605 ;
    RECT 0 80.675 0.070 80.885 ;
    RECT 0 80.955 0.070 81.165 ;
    RECT 0 81.235 0.070 81.445 ;
    RECT 0 81.515 0.070 81.725 ;
    RECT 0 81.795 0.070 82.005 ;
    RECT 0 82.075 0.070 82.285 ;
    RECT 0 82.355 0.070 82.565 ;
    RECT 0 82.635 0.070 82.845 ;
    RECT 0 82.915 0.070 83.125 ;
    RECT 0 83.195 0.070 83.405 ;
    RECT 0 83.475 0.070 83.685 ;
    RECT 0 83.755 0.070 83.965 ;
    RECT 0 84.035 0.070 84.245 ;
    RECT 0 84.315 0.070 84.525 ;
    RECT 0 84.595 0.070 84.805 ;
    RECT 0 84.875 0.070 85.085 ;
    RECT 0 85.155 0.070 85.365 ;
    RECT 0 85.435 0.070 85.645 ;
    RECT 0 85.715 0.070 85.925 ;
    RECT 0 85.995 0.070 86.205 ;
    RECT 0 86.275 0.070 86.485 ;
    RECT 0 86.555 0.070 86.765 ;
    RECT 0 86.835 0.070 87.045 ;
    RECT 0 87.115 0.070 87.325 ;
    RECT 0 87.395 0.070 87.605 ;
    RECT 0 87.675 0.070 87.885 ;
    RECT 0 87.955 0.070 88.165 ;
    RECT 0 88.235 0.070 88.445 ;
    RECT 0 88.515 0.070 88.725 ;
    RECT 0 88.795 0.070 89.005 ;
    RECT 0 89.075 0.070 89.285 ;
    RECT 0 89.355 0.070 89.565 ;
    RECT 0 89.635 0.070 89.845 ;
    RECT 0 89.915 0.070 90.125 ;
    RECT 0 90.195 0.070 90.405 ;
    RECT 0 90.475 0.070 90.685 ;
    RECT 0 90.755 0.070 90.965 ;
    RECT 0 91.035 0.070 91.245 ;
    RECT 0 91.315 0.070 91.525 ;
    RECT 0 91.595 0.070 91.805 ;
    RECT 0 91.875 0.070 92.085 ;
    RECT 0 92.155 0.070 92.365 ;
    RECT 0 92.435 0.070 92.645 ;
    RECT 0 92.715 0.070 92.925 ;
    RECT 0 92.995 0.070 93.205 ;
    RECT 0 93.275 0.070 93.485 ;
    RECT 0 93.555 0.070 93.765 ;
    RECT 0 93.835 0.070 94.045 ;
    RECT 0 94.115 0.070 94.325 ;
    RECT 0 94.395 0.070 94.605 ;
    RECT 0 94.675 0.070 94.885 ;
    RECT 0 94.955 0.070 95.165 ;
    RECT 0 95.235 0.070 95.445 ;
    RECT 0 95.515 0.070 95.725 ;
    RECT 0 95.795 0.070 96.005 ;
    RECT 0 96.075 0.070 96.285 ;
    RECT 0 96.355 0.070 96.565 ;
    RECT 0 96.635 0.070 96.845 ;
    RECT 0 96.915 0.070 105.105 ;
    RECT 0 105.175 0.070 105.385 ;
    RECT 0 105.455 0.070 105.665 ;
    RECT 0 105.735 0.070 105.945 ;
    RECT 0 106.015 0.070 106.225 ;
    RECT 0 106.295 0.070 106.505 ;
    RECT 0 106.575 0.070 106.785 ;
    RECT 0 106.855 0.070 107.065 ;
    RECT 0 107.135 0.070 115.325 ;
    RECT 0 115.395 0.070 115.605 ;
    RECT 0 115.675 0.070 115.885 ;
    RECT 0 115.955 0.070 119.000 ;
    LAYER metal4 ;
    RECT 0 0 115.140 1.400 ;
    RECT 0 117.600 115.140 119.000 ;
    RECT 0.000 1.400 1.260 117.600 ;
    RECT 1.540 1.400 2.380 117.600 ;
    RECT 2.660 1.400 3.500 117.600 ;
    RECT 3.780 1.400 4.620 117.600 ;
    RECT 4.900 1.400 5.740 117.600 ;
    RECT 6.020 1.400 6.860 117.600 ;
    RECT 7.140 1.400 7.980 117.600 ;
    RECT 8.260 1.400 9.100 117.600 ;
    RECT 9.380 1.400 10.220 117.600 ;
    RECT 10.500 1.400 11.340 117.600 ;
    RECT 11.620 1.400 12.460 117.600 ;
    RECT 12.740 1.400 13.580 117.600 ;
    RECT 13.860 1.400 14.700 117.600 ;
    RECT 14.980 1.400 15.820 117.600 ;
    RECT 16.100 1.400 16.940 117.600 ;
    RECT 17.220 1.400 18.060 117.600 ;
    RECT 18.340 1.400 19.180 117.600 ;
    RECT 19.460 1.400 20.300 117.600 ;
    RECT 20.580 1.400 21.420 117.600 ;
    RECT 21.700 1.400 22.540 117.600 ;
    RECT 22.820 1.400 23.660 117.600 ;
    RECT 23.940 1.400 24.780 117.600 ;
    RECT 25.060 1.400 25.900 117.600 ;
    RECT 26.180 1.400 27.020 117.600 ;
    RECT 27.300 1.400 28.140 117.600 ;
    RECT 28.420 1.400 29.260 117.600 ;
    RECT 29.540 1.400 30.380 117.600 ;
    RECT 30.660 1.400 31.500 117.600 ;
    RECT 31.780 1.400 32.620 117.600 ;
    RECT 32.900 1.400 33.740 117.600 ;
    RECT 34.020 1.400 34.860 117.600 ;
    RECT 35.140 1.400 35.980 117.600 ;
    RECT 36.260 1.400 37.100 117.600 ;
    RECT 37.380 1.400 38.220 117.600 ;
    RECT 38.500 1.400 39.340 117.600 ;
    RECT 39.620 1.400 40.460 117.600 ;
    RECT 40.740 1.400 41.580 117.600 ;
    RECT 41.860 1.400 42.700 117.600 ;
    RECT 42.980 1.400 43.820 117.600 ;
    RECT 44.100 1.400 44.940 117.600 ;
    RECT 45.220 1.400 46.060 117.600 ;
    RECT 46.340 1.400 47.180 117.600 ;
    RECT 47.460 1.400 48.300 117.600 ;
    RECT 48.580 1.400 49.420 117.600 ;
    RECT 49.700 1.400 50.540 117.600 ;
    RECT 50.820 1.400 51.660 117.600 ;
    RECT 51.940 1.400 52.780 117.600 ;
    RECT 53.060 1.400 53.900 117.600 ;
    RECT 54.180 1.400 55.020 117.600 ;
    RECT 55.300 1.400 56.140 117.600 ;
    RECT 56.420 1.400 57.260 117.600 ;
    RECT 57.540 1.400 58.380 117.600 ;
    RECT 58.660 1.400 59.500 117.600 ;
    RECT 59.780 1.400 60.620 117.600 ;
    RECT 60.900 1.400 61.740 117.600 ;
    RECT 62.020 1.400 62.860 117.600 ;
    RECT 63.140 1.400 63.980 117.600 ;
    RECT 64.260 1.400 65.100 117.600 ;
    RECT 65.380 1.400 66.220 117.600 ;
    RECT 66.500 1.400 67.340 117.600 ;
    RECT 67.620 1.400 68.460 117.600 ;
    RECT 68.740 1.400 69.580 117.600 ;
    RECT 69.860 1.400 70.700 117.600 ;
    RECT 70.980 1.400 71.820 117.600 ;
    RECT 72.100 1.400 72.940 117.600 ;
    RECT 73.220 1.400 74.060 117.600 ;
    RECT 74.340 1.400 75.180 117.600 ;
    RECT 75.460 1.400 76.300 117.600 ;
    RECT 76.580 1.400 77.420 117.600 ;
    RECT 77.700 1.400 78.540 117.600 ;
    RECT 78.820 1.400 79.660 117.600 ;
    RECT 79.940 1.400 80.780 117.600 ;
    RECT 81.060 1.400 81.900 117.600 ;
    RECT 82.180 1.400 83.020 117.600 ;
    RECT 83.300 1.400 84.140 117.600 ;
    RECT 84.420 1.400 85.260 117.600 ;
    RECT 85.540 1.400 86.380 117.600 ;
    RECT 86.660 1.400 87.500 117.600 ;
    RECT 87.780 1.400 88.620 117.600 ;
    RECT 88.900 1.400 89.740 117.600 ;
    RECT 90.020 1.400 90.860 117.600 ;
    RECT 91.140 1.400 91.980 117.600 ;
    RECT 92.260 1.400 93.100 117.600 ;
    RECT 93.380 1.400 94.220 117.600 ;
    RECT 94.500 1.400 95.340 117.600 ;
    RECT 95.620 1.400 96.460 117.600 ;
    RECT 96.740 1.400 97.580 117.600 ;
    RECT 97.860 1.400 98.700 117.600 ;
    RECT 98.980 1.400 99.820 117.600 ;
    RECT 100.100 1.400 100.940 117.600 ;
    RECT 101.220 1.400 102.060 117.600 ;
    RECT 102.340 1.400 103.180 117.600 ;
    RECT 103.460 1.400 104.300 117.600 ;
    RECT 104.580 1.400 105.420 117.600 ;
    RECT 105.700 1.400 106.540 117.600 ;
    RECT 106.820 1.400 107.660 117.600 ;
    RECT 107.940 1.400 108.780 117.600 ;
    RECT 109.060 1.400 109.900 117.600 ;
    RECT 110.180 1.400 111.020 117.600 ;
    RECT 111.300 1.400 112.140 117.600 ;
    RECT 112.420 1.400 113.260 117.600 ;
    RECT 113.540 1.400 115.140 117.600 ;
    LAYER OVERLAP ;
    RECT 0 0 115.140 119.000 ;
  END
END fakeram45_256x95

END LIBRARY
