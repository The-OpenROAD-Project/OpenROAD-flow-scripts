module MockArray(
  input        clock,
  input        reset,
  input  [7:0] io_insHorizontal_0_0,
  input  [7:0] io_insHorizontal_1_0,
  output [7:0] io_outsHorizontal_0_0,
  output [7:0] io_outsHorizontal_1_0,
  input  [7:0] io_insVertical_0_0,
  input  [7:0] io_insVertical_0_1,
  input  [7:0] io_insVertical_0_2,
  input  [7:0] io_insVertical_0_3,
  input  [7:0] io_insVertical_0_4,
  input  [7:0] io_insVertical_0_5,
  input  [7:0] io_insVertical_0_6,
  input  [7:0] io_insVertical_0_7,
  input  [7:0] io_insVertical_0_8,
  input  [7:0] io_insVertical_0_9,
  input  [7:0] io_insVertical_0_10,
  input  [7:0] io_insVertical_0_11,
  input  [7:0] io_insVertical_0_12,
  input  [7:0] io_insVertical_0_13,
  input  [7:0] io_insVertical_0_14,
  input  [7:0] io_insVertical_0_15,
  input  [7:0] io_insVertical_0_16,
  input  [7:0] io_insVertical_0_17,
  input  [7:0] io_insVertical_0_18,
  input  [7:0] io_insVertical_0_19,
  input  [7:0] io_insVertical_0_20,
  input  [7:0] io_insVertical_0_21,
  input  [7:0] io_insVertical_0_22,
  input  [7:0] io_insVertical_0_23,
  input  [7:0] io_insVertical_0_24,
  input  [7:0] io_insVertical_0_25,
  input  [7:0] io_insVertical_0_26,
  input  [7:0] io_insVertical_0_27,
  input  [7:0] io_insVertical_0_28,
  input  [7:0] io_insVertical_0_29,
  input  [7:0] io_insVertical_0_30,
  input  [7:0] io_insVertical_0_31,
  input  [7:0] io_insVertical_1_0,
  input  [7:0] io_insVertical_1_1,
  input  [7:0] io_insVertical_1_2,
  input  [7:0] io_insVertical_1_3,
  input  [7:0] io_insVertical_1_4,
  input  [7:0] io_insVertical_1_5,
  input  [7:0] io_insVertical_1_6,
  input  [7:0] io_insVertical_1_7,
  input  [7:0] io_insVertical_1_8,
  input  [7:0] io_insVertical_1_9,
  input  [7:0] io_insVertical_1_10,
  input  [7:0] io_insVertical_1_11,
  input  [7:0] io_insVertical_1_12,
  input  [7:0] io_insVertical_1_13,
  input  [7:0] io_insVertical_1_14,
  input  [7:0] io_insVertical_1_15,
  input  [7:0] io_insVertical_1_16,
  input  [7:0] io_insVertical_1_17,
  input  [7:0] io_insVertical_1_18,
  input  [7:0] io_insVertical_1_19,
  input  [7:0] io_insVertical_1_20,
  input  [7:0] io_insVertical_1_21,
  input  [7:0] io_insVertical_1_22,
  input  [7:0] io_insVertical_1_23,
  input  [7:0] io_insVertical_1_24,
  input  [7:0] io_insVertical_1_25,
  input  [7:0] io_insVertical_1_26,
  input  [7:0] io_insVertical_1_27,
  input  [7:0] io_insVertical_1_28,
  input  [7:0] io_insVertical_1_29,
  input  [7:0] io_insVertical_1_30,
  input  [7:0] io_insVertical_1_31,
  output [7:0] io_outsVertical_0_0,
  output [7:0] io_outsVertical_0_1,
  output [7:0] io_outsVertical_0_2,
  output [7:0] io_outsVertical_0_3,
  output [7:0] io_outsVertical_0_4,
  output [7:0] io_outsVertical_0_5,
  output [7:0] io_outsVertical_0_6,
  output [7:0] io_outsVertical_0_7,
  output [7:0] io_outsVertical_0_8,
  output [7:0] io_outsVertical_0_9,
  output [7:0] io_outsVertical_0_10,
  output [7:0] io_outsVertical_0_11,
  output [7:0] io_outsVertical_0_12,
  output [7:0] io_outsVertical_0_13,
  output [7:0] io_outsVertical_0_14,
  output [7:0] io_outsVertical_0_15,
  output [7:0] io_outsVertical_0_16,
  output [7:0] io_outsVertical_0_17,
  output [7:0] io_outsVertical_0_18,
  output [7:0] io_outsVertical_0_19,
  output [7:0] io_outsVertical_0_20,
  output [7:0] io_outsVertical_0_21,
  output [7:0] io_outsVertical_0_22,
  output [7:0] io_outsVertical_0_23,
  output [7:0] io_outsVertical_0_24,
  output [7:0] io_outsVertical_0_25,
  output [7:0] io_outsVertical_0_26,
  output [7:0] io_outsVertical_0_27,
  output [7:0] io_outsVertical_0_28,
  output [7:0] io_outsVertical_0_29,
  output [7:0] io_outsVertical_0_30,
  output [7:0] io_outsVertical_0_31,
  output [7:0] io_outsVertical_1_0,
  output [7:0] io_outsVertical_1_1,
  output [7:0] io_outsVertical_1_2,
  output [7:0] io_outsVertical_1_3,
  output [7:0] io_outsVertical_1_4,
  output [7:0] io_outsVertical_1_5,
  output [7:0] io_outsVertical_1_6,
  output [7:0] io_outsVertical_1_7,
  output [7:0] io_outsVertical_1_8,
  output [7:0] io_outsVertical_1_9,
  output [7:0] io_outsVertical_1_10,
  output [7:0] io_outsVertical_1_11,
  output [7:0] io_outsVertical_1_12,
  output [7:0] io_outsVertical_1_13,
  output [7:0] io_outsVertical_1_14,
  output [7:0] io_outsVertical_1_15,
  output [7:0] io_outsVertical_1_16,
  output [7:0] io_outsVertical_1_17,
  output [7:0] io_outsVertical_1_18,
  output [7:0] io_outsVertical_1_19,
  output [7:0] io_outsVertical_1_20,
  output [7:0] io_outsVertical_1_21,
  output [7:0] io_outsVertical_1_22,
  output [7:0] io_outsVertical_1_23,
  output [7:0] io_outsVertical_1_24,
  output [7:0] io_outsVertical_1_25,
  output [7:0] io_outsVertical_1_26,
  output [7:0] io_outsVertical_1_27,
  output [7:0] io_outsVertical_1_28,
  output [7:0] io_outsVertical_1_29,
  output [7:0] io_outsVertical_1_30,
  output [7:0] io_outsVertical_1_31,
  output       io_lsbs_0,
  output       io_lsbs_1,
  output       io_lsbs_2,
  output       io_lsbs_3,
  output       io_lsbs_4,
  output       io_lsbs_5,
  output       io_lsbs_6,
  output       io_lsbs_7,
  output       io_lsbs_8,
  output       io_lsbs_9,
  output       io_lsbs_10,
  output       io_lsbs_11,
  output       io_lsbs_12,
  output       io_lsbs_13,
  output       io_lsbs_14,
  output       io_lsbs_15,
  output       io_lsbs_16,
  output       io_lsbs_17,
  output       io_lsbs_18,
  output       io_lsbs_19,
  output       io_lsbs_20,
  output       io_lsbs_21,
  output       io_lsbs_22,
  output       io_lsbs_23,
  output       io_lsbs_24,
  output       io_lsbs_25,
  output       io_lsbs_26,
  output       io_lsbs_27,
  output       io_lsbs_28,
  output       io_lsbs_29,
  output       io_lsbs_30,
  output       io_lsbs_31
);
  wire  ces_0_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_0_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_1_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_1_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_2_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_2_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_3_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_3_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_4_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_4_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_5_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_5_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_6_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_6_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_7_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_7_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_8_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_8_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_9_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_9_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_10_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_10_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_11_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_11_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_12_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_12_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_13_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_13_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_14_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_14_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_15_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_15_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_16_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_16_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_17_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_17_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_18_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_18_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_19_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_19_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_20_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_20_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_21_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_21_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_22_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_22_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_23_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_23_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_24_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_24_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_25_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_25_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_26_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_26_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_27_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_27_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_28_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_28_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_29_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_29_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_30_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_30_0_io_outs_3; // @[MockArray.scala 36:52]
  wire  ces_31_0_clock; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_ins_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_ins_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_ins_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_ins_3; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_outs_0; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_outs_1; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_outs_2; // @[MockArray.scala 36:52]
  wire [7:0] ces_31_0_io_outs_3; // @[MockArray.scala 36:52]
  Element ces_0_0 ( // @[MockArray.scala 36:52]
    .clock(ces_0_0_clock),
    .io_ins_0(ces_0_0_io_ins_0),
    .io_ins_1(ces_0_0_io_ins_1),
    .io_ins_2(ces_0_0_io_ins_2),
    .io_ins_3(ces_0_0_io_ins_3),
    .io_outs_0(ces_0_0_io_outs_0),
    .io_outs_1(ces_0_0_io_outs_1),
    .io_outs_2(ces_0_0_io_outs_2),
    .io_outs_3(ces_0_0_io_outs_3)
  );
  Element ces_1_0 ( // @[MockArray.scala 36:52]
    .clock(ces_1_0_clock),
    .io_ins_0(ces_1_0_io_ins_0),
    .io_ins_1(ces_1_0_io_ins_1),
    .io_ins_2(ces_1_0_io_ins_2),
    .io_ins_3(ces_1_0_io_ins_3),
    .io_outs_0(ces_1_0_io_outs_0),
    .io_outs_1(ces_1_0_io_outs_1),
    .io_outs_2(ces_1_0_io_outs_2),
    .io_outs_3(ces_1_0_io_outs_3)
  );
  Element ces_2_0 ( // @[MockArray.scala 36:52]
    .clock(ces_2_0_clock),
    .io_ins_0(ces_2_0_io_ins_0),
    .io_ins_1(ces_2_0_io_ins_1),
    .io_ins_2(ces_2_0_io_ins_2),
    .io_ins_3(ces_2_0_io_ins_3),
    .io_outs_0(ces_2_0_io_outs_0),
    .io_outs_1(ces_2_0_io_outs_1),
    .io_outs_2(ces_2_0_io_outs_2),
    .io_outs_3(ces_2_0_io_outs_3)
  );
  Element ces_3_0 ( // @[MockArray.scala 36:52]
    .clock(ces_3_0_clock),
    .io_ins_0(ces_3_0_io_ins_0),
    .io_ins_1(ces_3_0_io_ins_1),
    .io_ins_2(ces_3_0_io_ins_2),
    .io_ins_3(ces_3_0_io_ins_3),
    .io_outs_0(ces_3_0_io_outs_0),
    .io_outs_1(ces_3_0_io_outs_1),
    .io_outs_2(ces_3_0_io_outs_2),
    .io_outs_3(ces_3_0_io_outs_3)
  );
  Element ces_4_0 ( // @[MockArray.scala 36:52]
    .clock(ces_4_0_clock),
    .io_ins_0(ces_4_0_io_ins_0),
    .io_ins_1(ces_4_0_io_ins_1),
    .io_ins_2(ces_4_0_io_ins_2),
    .io_ins_3(ces_4_0_io_ins_3),
    .io_outs_0(ces_4_0_io_outs_0),
    .io_outs_1(ces_4_0_io_outs_1),
    .io_outs_2(ces_4_0_io_outs_2),
    .io_outs_3(ces_4_0_io_outs_3)
  );
  Element ces_5_0 ( // @[MockArray.scala 36:52]
    .clock(ces_5_0_clock),
    .io_ins_0(ces_5_0_io_ins_0),
    .io_ins_1(ces_5_0_io_ins_1),
    .io_ins_2(ces_5_0_io_ins_2),
    .io_ins_3(ces_5_0_io_ins_3),
    .io_outs_0(ces_5_0_io_outs_0),
    .io_outs_1(ces_5_0_io_outs_1),
    .io_outs_2(ces_5_0_io_outs_2),
    .io_outs_3(ces_5_0_io_outs_3)
  );
  Element ces_6_0 ( // @[MockArray.scala 36:52]
    .clock(ces_6_0_clock),
    .io_ins_0(ces_6_0_io_ins_0),
    .io_ins_1(ces_6_0_io_ins_1),
    .io_ins_2(ces_6_0_io_ins_2),
    .io_ins_3(ces_6_0_io_ins_3),
    .io_outs_0(ces_6_0_io_outs_0),
    .io_outs_1(ces_6_0_io_outs_1),
    .io_outs_2(ces_6_0_io_outs_2),
    .io_outs_3(ces_6_0_io_outs_3)
  );
  Element ces_7_0 ( // @[MockArray.scala 36:52]
    .clock(ces_7_0_clock),
    .io_ins_0(ces_7_0_io_ins_0),
    .io_ins_1(ces_7_0_io_ins_1),
    .io_ins_2(ces_7_0_io_ins_2),
    .io_ins_3(ces_7_0_io_ins_3),
    .io_outs_0(ces_7_0_io_outs_0),
    .io_outs_1(ces_7_0_io_outs_1),
    .io_outs_2(ces_7_0_io_outs_2),
    .io_outs_3(ces_7_0_io_outs_3)
  );
  Element ces_8_0 ( // @[MockArray.scala 36:52]
    .clock(ces_8_0_clock),
    .io_ins_0(ces_8_0_io_ins_0),
    .io_ins_1(ces_8_0_io_ins_1),
    .io_ins_2(ces_8_0_io_ins_2),
    .io_ins_3(ces_8_0_io_ins_3),
    .io_outs_0(ces_8_0_io_outs_0),
    .io_outs_1(ces_8_0_io_outs_1),
    .io_outs_2(ces_8_0_io_outs_2),
    .io_outs_3(ces_8_0_io_outs_3)
  );
  Element ces_9_0 ( // @[MockArray.scala 36:52]
    .clock(ces_9_0_clock),
    .io_ins_0(ces_9_0_io_ins_0),
    .io_ins_1(ces_9_0_io_ins_1),
    .io_ins_2(ces_9_0_io_ins_2),
    .io_ins_3(ces_9_0_io_ins_3),
    .io_outs_0(ces_9_0_io_outs_0),
    .io_outs_1(ces_9_0_io_outs_1),
    .io_outs_2(ces_9_0_io_outs_2),
    .io_outs_3(ces_9_0_io_outs_3)
  );
  Element ces_10_0 ( // @[MockArray.scala 36:52]
    .clock(ces_10_0_clock),
    .io_ins_0(ces_10_0_io_ins_0),
    .io_ins_1(ces_10_0_io_ins_1),
    .io_ins_2(ces_10_0_io_ins_2),
    .io_ins_3(ces_10_0_io_ins_3),
    .io_outs_0(ces_10_0_io_outs_0),
    .io_outs_1(ces_10_0_io_outs_1),
    .io_outs_2(ces_10_0_io_outs_2),
    .io_outs_3(ces_10_0_io_outs_3)
  );
  Element ces_11_0 ( // @[MockArray.scala 36:52]
    .clock(ces_11_0_clock),
    .io_ins_0(ces_11_0_io_ins_0),
    .io_ins_1(ces_11_0_io_ins_1),
    .io_ins_2(ces_11_0_io_ins_2),
    .io_ins_3(ces_11_0_io_ins_3),
    .io_outs_0(ces_11_0_io_outs_0),
    .io_outs_1(ces_11_0_io_outs_1),
    .io_outs_2(ces_11_0_io_outs_2),
    .io_outs_3(ces_11_0_io_outs_3)
  );
  Element ces_12_0 ( // @[MockArray.scala 36:52]
    .clock(ces_12_0_clock),
    .io_ins_0(ces_12_0_io_ins_0),
    .io_ins_1(ces_12_0_io_ins_1),
    .io_ins_2(ces_12_0_io_ins_2),
    .io_ins_3(ces_12_0_io_ins_3),
    .io_outs_0(ces_12_0_io_outs_0),
    .io_outs_1(ces_12_0_io_outs_1),
    .io_outs_2(ces_12_0_io_outs_2),
    .io_outs_3(ces_12_0_io_outs_3)
  );
  Element ces_13_0 ( // @[MockArray.scala 36:52]
    .clock(ces_13_0_clock),
    .io_ins_0(ces_13_0_io_ins_0),
    .io_ins_1(ces_13_0_io_ins_1),
    .io_ins_2(ces_13_0_io_ins_2),
    .io_ins_3(ces_13_0_io_ins_3),
    .io_outs_0(ces_13_0_io_outs_0),
    .io_outs_1(ces_13_0_io_outs_1),
    .io_outs_2(ces_13_0_io_outs_2),
    .io_outs_3(ces_13_0_io_outs_3)
  );
  Element ces_14_0 ( // @[MockArray.scala 36:52]
    .clock(ces_14_0_clock),
    .io_ins_0(ces_14_0_io_ins_0),
    .io_ins_1(ces_14_0_io_ins_1),
    .io_ins_2(ces_14_0_io_ins_2),
    .io_ins_3(ces_14_0_io_ins_3),
    .io_outs_0(ces_14_0_io_outs_0),
    .io_outs_1(ces_14_0_io_outs_1),
    .io_outs_2(ces_14_0_io_outs_2),
    .io_outs_3(ces_14_0_io_outs_3)
  );
  Element ces_15_0 ( // @[MockArray.scala 36:52]
    .clock(ces_15_0_clock),
    .io_ins_0(ces_15_0_io_ins_0),
    .io_ins_1(ces_15_0_io_ins_1),
    .io_ins_2(ces_15_0_io_ins_2),
    .io_ins_3(ces_15_0_io_ins_3),
    .io_outs_0(ces_15_0_io_outs_0),
    .io_outs_1(ces_15_0_io_outs_1),
    .io_outs_2(ces_15_0_io_outs_2),
    .io_outs_3(ces_15_0_io_outs_3)
  );
  Element ces_16_0 ( // @[MockArray.scala 36:52]
    .clock(ces_16_0_clock),
    .io_ins_0(ces_16_0_io_ins_0),
    .io_ins_1(ces_16_0_io_ins_1),
    .io_ins_2(ces_16_0_io_ins_2),
    .io_ins_3(ces_16_0_io_ins_3),
    .io_outs_0(ces_16_0_io_outs_0),
    .io_outs_1(ces_16_0_io_outs_1),
    .io_outs_2(ces_16_0_io_outs_2),
    .io_outs_3(ces_16_0_io_outs_3)
  );
  Element ces_17_0 ( // @[MockArray.scala 36:52]
    .clock(ces_17_0_clock),
    .io_ins_0(ces_17_0_io_ins_0),
    .io_ins_1(ces_17_0_io_ins_1),
    .io_ins_2(ces_17_0_io_ins_2),
    .io_ins_3(ces_17_0_io_ins_3),
    .io_outs_0(ces_17_0_io_outs_0),
    .io_outs_1(ces_17_0_io_outs_1),
    .io_outs_2(ces_17_0_io_outs_2),
    .io_outs_3(ces_17_0_io_outs_3)
  );
  Element ces_18_0 ( // @[MockArray.scala 36:52]
    .clock(ces_18_0_clock),
    .io_ins_0(ces_18_0_io_ins_0),
    .io_ins_1(ces_18_0_io_ins_1),
    .io_ins_2(ces_18_0_io_ins_2),
    .io_ins_3(ces_18_0_io_ins_3),
    .io_outs_0(ces_18_0_io_outs_0),
    .io_outs_1(ces_18_0_io_outs_1),
    .io_outs_2(ces_18_0_io_outs_2),
    .io_outs_3(ces_18_0_io_outs_3)
  );
  Element ces_19_0 ( // @[MockArray.scala 36:52]
    .clock(ces_19_0_clock),
    .io_ins_0(ces_19_0_io_ins_0),
    .io_ins_1(ces_19_0_io_ins_1),
    .io_ins_2(ces_19_0_io_ins_2),
    .io_ins_3(ces_19_0_io_ins_3),
    .io_outs_0(ces_19_0_io_outs_0),
    .io_outs_1(ces_19_0_io_outs_1),
    .io_outs_2(ces_19_0_io_outs_2),
    .io_outs_3(ces_19_0_io_outs_3)
  );
  Element ces_20_0 ( // @[MockArray.scala 36:52]
    .clock(ces_20_0_clock),
    .io_ins_0(ces_20_0_io_ins_0),
    .io_ins_1(ces_20_0_io_ins_1),
    .io_ins_2(ces_20_0_io_ins_2),
    .io_ins_3(ces_20_0_io_ins_3),
    .io_outs_0(ces_20_0_io_outs_0),
    .io_outs_1(ces_20_0_io_outs_1),
    .io_outs_2(ces_20_0_io_outs_2),
    .io_outs_3(ces_20_0_io_outs_3)
  );
  Element ces_21_0 ( // @[MockArray.scala 36:52]
    .clock(ces_21_0_clock),
    .io_ins_0(ces_21_0_io_ins_0),
    .io_ins_1(ces_21_0_io_ins_1),
    .io_ins_2(ces_21_0_io_ins_2),
    .io_ins_3(ces_21_0_io_ins_3),
    .io_outs_0(ces_21_0_io_outs_0),
    .io_outs_1(ces_21_0_io_outs_1),
    .io_outs_2(ces_21_0_io_outs_2),
    .io_outs_3(ces_21_0_io_outs_3)
  );
  Element ces_22_0 ( // @[MockArray.scala 36:52]
    .clock(ces_22_0_clock),
    .io_ins_0(ces_22_0_io_ins_0),
    .io_ins_1(ces_22_0_io_ins_1),
    .io_ins_2(ces_22_0_io_ins_2),
    .io_ins_3(ces_22_0_io_ins_3),
    .io_outs_0(ces_22_0_io_outs_0),
    .io_outs_1(ces_22_0_io_outs_1),
    .io_outs_2(ces_22_0_io_outs_2),
    .io_outs_3(ces_22_0_io_outs_3)
  );
  Element ces_23_0 ( // @[MockArray.scala 36:52]
    .clock(ces_23_0_clock),
    .io_ins_0(ces_23_0_io_ins_0),
    .io_ins_1(ces_23_0_io_ins_1),
    .io_ins_2(ces_23_0_io_ins_2),
    .io_ins_3(ces_23_0_io_ins_3),
    .io_outs_0(ces_23_0_io_outs_0),
    .io_outs_1(ces_23_0_io_outs_1),
    .io_outs_2(ces_23_0_io_outs_2),
    .io_outs_3(ces_23_0_io_outs_3)
  );
  Element ces_24_0 ( // @[MockArray.scala 36:52]
    .clock(ces_24_0_clock),
    .io_ins_0(ces_24_0_io_ins_0),
    .io_ins_1(ces_24_0_io_ins_1),
    .io_ins_2(ces_24_0_io_ins_2),
    .io_ins_3(ces_24_0_io_ins_3),
    .io_outs_0(ces_24_0_io_outs_0),
    .io_outs_1(ces_24_0_io_outs_1),
    .io_outs_2(ces_24_0_io_outs_2),
    .io_outs_3(ces_24_0_io_outs_3)
  );
  Element ces_25_0 ( // @[MockArray.scala 36:52]
    .clock(ces_25_0_clock),
    .io_ins_0(ces_25_0_io_ins_0),
    .io_ins_1(ces_25_0_io_ins_1),
    .io_ins_2(ces_25_0_io_ins_2),
    .io_ins_3(ces_25_0_io_ins_3),
    .io_outs_0(ces_25_0_io_outs_0),
    .io_outs_1(ces_25_0_io_outs_1),
    .io_outs_2(ces_25_0_io_outs_2),
    .io_outs_3(ces_25_0_io_outs_3)
  );
  Element ces_26_0 ( // @[MockArray.scala 36:52]
    .clock(ces_26_0_clock),
    .io_ins_0(ces_26_0_io_ins_0),
    .io_ins_1(ces_26_0_io_ins_1),
    .io_ins_2(ces_26_0_io_ins_2),
    .io_ins_3(ces_26_0_io_ins_3),
    .io_outs_0(ces_26_0_io_outs_0),
    .io_outs_1(ces_26_0_io_outs_1),
    .io_outs_2(ces_26_0_io_outs_2),
    .io_outs_3(ces_26_0_io_outs_3)
  );
  Element ces_27_0 ( // @[MockArray.scala 36:52]
    .clock(ces_27_0_clock),
    .io_ins_0(ces_27_0_io_ins_0),
    .io_ins_1(ces_27_0_io_ins_1),
    .io_ins_2(ces_27_0_io_ins_2),
    .io_ins_3(ces_27_0_io_ins_3),
    .io_outs_0(ces_27_0_io_outs_0),
    .io_outs_1(ces_27_0_io_outs_1),
    .io_outs_2(ces_27_0_io_outs_2),
    .io_outs_3(ces_27_0_io_outs_3)
  );
  Element ces_28_0 ( // @[MockArray.scala 36:52]
    .clock(ces_28_0_clock),
    .io_ins_0(ces_28_0_io_ins_0),
    .io_ins_1(ces_28_0_io_ins_1),
    .io_ins_2(ces_28_0_io_ins_2),
    .io_ins_3(ces_28_0_io_ins_3),
    .io_outs_0(ces_28_0_io_outs_0),
    .io_outs_1(ces_28_0_io_outs_1),
    .io_outs_2(ces_28_0_io_outs_2),
    .io_outs_3(ces_28_0_io_outs_3)
  );
  Element ces_29_0 ( // @[MockArray.scala 36:52]
    .clock(ces_29_0_clock),
    .io_ins_0(ces_29_0_io_ins_0),
    .io_ins_1(ces_29_0_io_ins_1),
    .io_ins_2(ces_29_0_io_ins_2),
    .io_ins_3(ces_29_0_io_ins_3),
    .io_outs_0(ces_29_0_io_outs_0),
    .io_outs_1(ces_29_0_io_outs_1),
    .io_outs_2(ces_29_0_io_outs_2),
    .io_outs_3(ces_29_0_io_outs_3)
  );
  Element ces_30_0 ( // @[MockArray.scala 36:52]
    .clock(ces_30_0_clock),
    .io_ins_0(ces_30_0_io_ins_0),
    .io_ins_1(ces_30_0_io_ins_1),
    .io_ins_2(ces_30_0_io_ins_2),
    .io_ins_3(ces_30_0_io_ins_3),
    .io_outs_0(ces_30_0_io_outs_0),
    .io_outs_1(ces_30_0_io_outs_1),
    .io_outs_2(ces_30_0_io_outs_2),
    .io_outs_3(ces_30_0_io_outs_3)
  );
  Element ces_31_0 ( // @[MockArray.scala 36:52]
    .clock(ces_31_0_clock),
    .io_ins_0(ces_31_0_io_ins_0),
    .io_ins_1(ces_31_0_io_ins_1),
    .io_ins_2(ces_31_0_io_ins_2),
    .io_ins_3(ces_31_0_io_ins_3),
    .io_outs_0(ces_31_0_io_outs_0),
    .io_outs_1(ces_31_0_io_outs_1),
    .io_outs_2(ces_31_0_io_outs_2),
    .io_outs_3(ces_31_0_io_outs_3)
  );
  assign io_outsHorizontal_0_0 = ces_0_0_io_outs_0; // @[MockArray.scala 49:89]
  assign io_outsHorizontal_1_0 = ces_31_0_io_outs_2; // @[MockArray.scala 51:89]
  assign io_outsVertical_0_0 = ces_0_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_1 = ces_1_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_2 = ces_2_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_3 = ces_3_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_4 = ces_4_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_5 = ces_5_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_6 = ces_6_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_7 = ces_7_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_8 = ces_8_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_9 = ces_9_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_10 = ces_10_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_11 = ces_11_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_12 = ces_12_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_13 = ces_13_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_14 = ces_14_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_15 = ces_15_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_16 = ces_16_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_17 = ces_17_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_18 = ces_18_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_19 = ces_19_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_20 = ces_20_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_21 = ces_21_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_22 = ces_22_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_23 = ces_23_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_24 = ces_24_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_25 = ces_25_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_26 = ces_26_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_27 = ces_27_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_28 = ces_28_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_29 = ces_29_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_30 = ces_30_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_0_31 = ces_31_0_io_outs_1; // @[MockArray.scala 50:89]
  assign io_outsVertical_1_0 = ces_0_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_1 = ces_1_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_2 = ces_2_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_3 = ces_3_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_4 = ces_4_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_5 = ces_5_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_6 = ces_6_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_7 = ces_7_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_8 = ces_8_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_9 = ces_9_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_10 = ces_10_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_11 = ces_11_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_12 = ces_12_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_13 = ces_13_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_14 = ces_14_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_15 = ces_15_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_16 = ces_16_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_17 = ces_17_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_18 = ces_18_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_19 = ces_19_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_20 = ces_20_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_21 = ces_21_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_22 = ces_22_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_23 = ces_23_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_24 = ces_24_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_25 = ces_25_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_26 = ces_26_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_27 = ces_27_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_28 = ces_28_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_29 = ces_29_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_30 = ces_30_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_outsVertical_1_31 = ces_31_0_io_outs_3; // @[MockArray.scala 52:89]
  assign io_lsbs_0 = ces_0_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_1 = ces_1_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_2 = ces_2_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_3 = ces_3_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_4 = ces_4_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_5 = ces_5_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_6 = ces_6_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_7 = ces_7_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_8 = ces_8_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_9 = ces_9_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_10 = ces_10_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_11 = ces_11_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_12 = ces_12_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_13 = ces_13_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_14 = ces_14_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_15 = ces_15_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_16 = ces_16_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_17 = ces_17_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_18 = ces_18_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_19 = ces_19_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_20 = ces_20_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_21 = ces_21_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_22 = ces_22_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_23 = ces_23_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_24 = ces_24_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_25 = ces_25_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_26 = ces_26_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_27 = ces_27_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_28 = ces_28_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_29 = ces_29_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_30 = ces_30_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign io_lsbs_31 = ces_31_0_io_outs_0[0]; // @[MockArray.scala 38:44]
  assign ces_0_0_clock = clock;
  assign ces_0_0_io_ins_0 = io_insHorizontal_0_0; // @[MockArray.scala 44:87]
  assign ces_0_0_io_ins_1 = io_insVertical_0_0; // @[MockArray.scala 45:87]
  assign ces_0_0_io_ins_2 = ces_1_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_0_0_io_ins_3 = io_insVertical_1_0; // @[MockArray.scala 47:87]
  assign ces_1_0_clock = clock;
  assign ces_1_0_io_ins_0 = ces_0_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_1_0_io_ins_1 = io_insVertical_0_1; // @[MockArray.scala 45:87]
  assign ces_1_0_io_ins_2 = ces_2_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_1_0_io_ins_3 = io_insVertical_1_1; // @[MockArray.scala 47:87]
  assign ces_2_0_clock = clock;
  assign ces_2_0_io_ins_0 = ces_1_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_2_0_io_ins_1 = io_insVertical_0_2; // @[MockArray.scala 45:87]
  assign ces_2_0_io_ins_2 = ces_3_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_2_0_io_ins_3 = io_insVertical_1_2; // @[MockArray.scala 47:87]
  assign ces_3_0_clock = clock;
  assign ces_3_0_io_ins_0 = ces_2_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_3_0_io_ins_1 = io_insVertical_0_3; // @[MockArray.scala 45:87]
  assign ces_3_0_io_ins_2 = ces_4_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_3_0_io_ins_3 = io_insVertical_1_3; // @[MockArray.scala 47:87]
  assign ces_4_0_clock = clock;
  assign ces_4_0_io_ins_0 = ces_3_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_4_0_io_ins_1 = io_insVertical_0_4; // @[MockArray.scala 45:87]
  assign ces_4_0_io_ins_2 = ces_5_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_4_0_io_ins_3 = io_insVertical_1_4; // @[MockArray.scala 47:87]
  assign ces_5_0_clock = clock;
  assign ces_5_0_io_ins_0 = ces_4_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_5_0_io_ins_1 = io_insVertical_0_5; // @[MockArray.scala 45:87]
  assign ces_5_0_io_ins_2 = ces_6_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_5_0_io_ins_3 = io_insVertical_1_5; // @[MockArray.scala 47:87]
  assign ces_6_0_clock = clock;
  assign ces_6_0_io_ins_0 = ces_5_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_6_0_io_ins_1 = io_insVertical_0_6; // @[MockArray.scala 45:87]
  assign ces_6_0_io_ins_2 = ces_7_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_6_0_io_ins_3 = io_insVertical_1_6; // @[MockArray.scala 47:87]
  assign ces_7_0_clock = clock;
  assign ces_7_0_io_ins_0 = ces_6_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_7_0_io_ins_1 = io_insVertical_0_7; // @[MockArray.scala 45:87]
  assign ces_7_0_io_ins_2 = ces_8_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_7_0_io_ins_3 = io_insVertical_1_7; // @[MockArray.scala 47:87]
  assign ces_8_0_clock = clock;
  assign ces_8_0_io_ins_0 = ces_7_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_8_0_io_ins_1 = io_insVertical_0_8; // @[MockArray.scala 45:87]
  assign ces_8_0_io_ins_2 = ces_9_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_8_0_io_ins_3 = io_insVertical_1_8; // @[MockArray.scala 47:87]
  assign ces_9_0_clock = clock;
  assign ces_9_0_io_ins_0 = ces_8_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_9_0_io_ins_1 = io_insVertical_0_9; // @[MockArray.scala 45:87]
  assign ces_9_0_io_ins_2 = ces_10_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_9_0_io_ins_3 = io_insVertical_1_9; // @[MockArray.scala 47:87]
  assign ces_10_0_clock = clock;
  assign ces_10_0_io_ins_0 = ces_9_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_10_0_io_ins_1 = io_insVertical_0_10; // @[MockArray.scala 45:87]
  assign ces_10_0_io_ins_2 = ces_11_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_10_0_io_ins_3 = io_insVertical_1_10; // @[MockArray.scala 47:87]
  assign ces_11_0_clock = clock;
  assign ces_11_0_io_ins_0 = ces_10_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_11_0_io_ins_1 = io_insVertical_0_11; // @[MockArray.scala 45:87]
  assign ces_11_0_io_ins_2 = ces_12_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_11_0_io_ins_3 = io_insVertical_1_11; // @[MockArray.scala 47:87]
  assign ces_12_0_clock = clock;
  assign ces_12_0_io_ins_0 = ces_11_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_12_0_io_ins_1 = io_insVertical_0_12; // @[MockArray.scala 45:87]
  assign ces_12_0_io_ins_2 = ces_13_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_12_0_io_ins_3 = io_insVertical_1_12; // @[MockArray.scala 47:87]
  assign ces_13_0_clock = clock;
  assign ces_13_0_io_ins_0 = ces_12_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_13_0_io_ins_1 = io_insVertical_0_13; // @[MockArray.scala 45:87]
  assign ces_13_0_io_ins_2 = ces_14_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_13_0_io_ins_3 = io_insVertical_1_13; // @[MockArray.scala 47:87]
  assign ces_14_0_clock = clock;
  assign ces_14_0_io_ins_0 = ces_13_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_14_0_io_ins_1 = io_insVertical_0_14; // @[MockArray.scala 45:87]
  assign ces_14_0_io_ins_2 = ces_15_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_14_0_io_ins_3 = io_insVertical_1_14; // @[MockArray.scala 47:87]
  assign ces_15_0_clock = clock;
  assign ces_15_0_io_ins_0 = ces_14_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_15_0_io_ins_1 = io_insVertical_0_15; // @[MockArray.scala 45:87]
  assign ces_15_0_io_ins_2 = ces_16_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_15_0_io_ins_3 = io_insVertical_1_15; // @[MockArray.scala 47:87]
  assign ces_16_0_clock = clock;
  assign ces_16_0_io_ins_0 = ces_15_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_16_0_io_ins_1 = io_insVertical_0_16; // @[MockArray.scala 45:87]
  assign ces_16_0_io_ins_2 = ces_17_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_16_0_io_ins_3 = io_insVertical_1_16; // @[MockArray.scala 47:87]
  assign ces_17_0_clock = clock;
  assign ces_17_0_io_ins_0 = ces_16_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_17_0_io_ins_1 = io_insVertical_0_17; // @[MockArray.scala 45:87]
  assign ces_17_0_io_ins_2 = ces_18_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_17_0_io_ins_3 = io_insVertical_1_17; // @[MockArray.scala 47:87]
  assign ces_18_0_clock = clock;
  assign ces_18_0_io_ins_0 = ces_17_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_18_0_io_ins_1 = io_insVertical_0_18; // @[MockArray.scala 45:87]
  assign ces_18_0_io_ins_2 = ces_19_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_18_0_io_ins_3 = io_insVertical_1_18; // @[MockArray.scala 47:87]
  assign ces_19_0_clock = clock;
  assign ces_19_0_io_ins_0 = ces_18_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_19_0_io_ins_1 = io_insVertical_0_19; // @[MockArray.scala 45:87]
  assign ces_19_0_io_ins_2 = ces_20_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_19_0_io_ins_3 = io_insVertical_1_19; // @[MockArray.scala 47:87]
  assign ces_20_0_clock = clock;
  assign ces_20_0_io_ins_0 = ces_19_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_20_0_io_ins_1 = io_insVertical_0_20; // @[MockArray.scala 45:87]
  assign ces_20_0_io_ins_2 = ces_21_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_20_0_io_ins_3 = io_insVertical_1_20; // @[MockArray.scala 47:87]
  assign ces_21_0_clock = clock;
  assign ces_21_0_io_ins_0 = ces_20_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_21_0_io_ins_1 = io_insVertical_0_21; // @[MockArray.scala 45:87]
  assign ces_21_0_io_ins_2 = ces_22_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_21_0_io_ins_3 = io_insVertical_1_21; // @[MockArray.scala 47:87]
  assign ces_22_0_clock = clock;
  assign ces_22_0_io_ins_0 = ces_21_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_22_0_io_ins_1 = io_insVertical_0_22; // @[MockArray.scala 45:87]
  assign ces_22_0_io_ins_2 = ces_23_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_22_0_io_ins_3 = io_insVertical_1_22; // @[MockArray.scala 47:87]
  assign ces_23_0_clock = clock;
  assign ces_23_0_io_ins_0 = ces_22_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_23_0_io_ins_1 = io_insVertical_0_23; // @[MockArray.scala 45:87]
  assign ces_23_0_io_ins_2 = ces_24_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_23_0_io_ins_3 = io_insVertical_1_23; // @[MockArray.scala 47:87]
  assign ces_24_0_clock = clock;
  assign ces_24_0_io_ins_0 = ces_23_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_24_0_io_ins_1 = io_insVertical_0_24; // @[MockArray.scala 45:87]
  assign ces_24_0_io_ins_2 = ces_25_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_24_0_io_ins_3 = io_insVertical_1_24; // @[MockArray.scala 47:87]
  assign ces_25_0_clock = clock;
  assign ces_25_0_io_ins_0 = ces_24_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_25_0_io_ins_1 = io_insVertical_0_25; // @[MockArray.scala 45:87]
  assign ces_25_0_io_ins_2 = ces_26_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_25_0_io_ins_3 = io_insVertical_1_25; // @[MockArray.scala 47:87]
  assign ces_26_0_clock = clock;
  assign ces_26_0_io_ins_0 = ces_25_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_26_0_io_ins_1 = io_insVertical_0_26; // @[MockArray.scala 45:87]
  assign ces_26_0_io_ins_2 = ces_27_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_26_0_io_ins_3 = io_insVertical_1_26; // @[MockArray.scala 47:87]
  assign ces_27_0_clock = clock;
  assign ces_27_0_io_ins_0 = ces_26_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_27_0_io_ins_1 = io_insVertical_0_27; // @[MockArray.scala 45:87]
  assign ces_27_0_io_ins_2 = ces_28_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_27_0_io_ins_3 = io_insVertical_1_27; // @[MockArray.scala 47:87]
  assign ces_28_0_clock = clock;
  assign ces_28_0_io_ins_0 = ces_27_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_28_0_io_ins_1 = io_insVertical_0_28; // @[MockArray.scala 45:87]
  assign ces_28_0_io_ins_2 = ces_29_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_28_0_io_ins_3 = io_insVertical_1_28; // @[MockArray.scala 47:87]
  assign ces_29_0_clock = clock;
  assign ces_29_0_io_ins_0 = ces_28_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_29_0_io_ins_1 = io_insVertical_0_29; // @[MockArray.scala 45:87]
  assign ces_29_0_io_ins_2 = ces_30_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_29_0_io_ins_3 = io_insVertical_1_29; // @[MockArray.scala 47:87]
  assign ces_30_0_clock = clock;
  assign ces_30_0_io_ins_0 = ces_29_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_30_0_io_ins_1 = io_insVertical_0_30; // @[MockArray.scala 45:87]
  assign ces_30_0_io_ins_2 = ces_31_0_io_outs_0; // @[MockArray.scala 56:19]
  assign ces_30_0_io_ins_3 = io_insVertical_1_30; // @[MockArray.scala 47:87]
  assign ces_31_0_clock = clock;
  assign ces_31_0_io_ins_0 = ces_30_0_io_outs_2; // @[MockArray.scala 57:19]
  assign ces_31_0_io_ins_1 = io_insVertical_0_31; // @[MockArray.scala 45:87]
  assign ces_31_0_io_ins_2 = io_insHorizontal_1_0; // @[MockArray.scala 46:87]
  assign ces_31_0_io_ins_3 = io_insVertical_1_31; // @[MockArray.scala 47:87]
endmodule
