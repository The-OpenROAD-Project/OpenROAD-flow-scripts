../../../platforms/nangate45/lef/fakeram45_32x64.lef