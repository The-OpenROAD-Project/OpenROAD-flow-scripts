VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_64x7
  FOREIGN fakeram45_64x7 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 10.640 BY 36.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.400 0.070 1.470 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.380 0.070 2.450 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.360 0.070 3.430 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.340 0.070 4.410 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.320 0.070 5.390 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.300 0.070 6.370 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.280 0.070 7.350 ;
    END
  END w_mask_in[6]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.260 0.070 8.330 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.240 0.070 9.310 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.220 0.070 10.290 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.200 0.070 11.270 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.180 0.070 12.250 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.160 0.070 13.230 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.140 0.070 14.210 ;
    END
  END rd_out[6]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.120 0.070 15.190 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.100 0.070 16.170 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.080 0.070 17.150 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.060 0.070 18.130 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.040 0.070 19.110 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.020 0.070 20.090 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.000 0.070 21.070 ;
    END
  END wd_in[6]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.980 0.070 22.050 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.960 0.070 23.030 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.940 0.070 24.010 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.920 0.070 24.990 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.900 0.070 25.970 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.880 0.070 26.950 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.860 0.070 27.930 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.840 0.070 28.910 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.820 0.070 29.890 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 35.000 ;
      RECT 3.500 1.400 3.780 35.000 ;
      RECT 5.740 1.400 6.020 35.000 ;
      RECT 7.980 1.400 8.260 35.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 35.000 ;
      RECT 4.620 1.400 4.900 35.000 ;
      RECT 6.860 1.400 7.140 35.000 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 10.640 36.400 ;
    LAYER metal2 ;
    RECT 0 0 10.640 36.400 ;
    LAYER metal3 ;
    RECT 0.070 0 10.640 36.400 ;
    RECT 0 0.000 0.070 1.400 ;
    RECT 0 1.470 0.070 2.380 ;
    RECT 0 2.450 0.070 3.360 ;
    RECT 0 3.430 0.070 4.340 ;
    RECT 0 4.410 0.070 5.320 ;
    RECT 0 5.390 0.070 6.300 ;
    RECT 0 6.370 0.070 7.280 ;
    RECT 0 7.350 0.070 8.260 ;
    RECT 0 8.330 0.070 9.240 ;
    RECT 0 9.310 0.070 10.220 ;
    RECT 0 10.290 0.070 11.200 ;
    RECT 0 11.270 0.070 12.180 ;
    RECT 0 12.250 0.070 13.160 ;
    RECT 0 13.230 0.070 14.140 ;
    RECT 0 14.210 0.070 15.120 ;
    RECT 0 15.190 0.070 16.100 ;
    RECT 0 16.170 0.070 17.080 ;
    RECT 0 17.150 0.070 18.060 ;
    RECT 0 18.130 0.070 19.040 ;
    RECT 0 19.110 0.070 20.020 ;
    RECT 0 20.090 0.070 21.000 ;
    RECT 0 21.070 0.070 21.980 ;
    RECT 0 22.050 0.070 22.960 ;
    RECT 0 23.030 0.070 23.940 ;
    RECT 0 24.010 0.070 24.920 ;
    RECT 0 24.990 0.070 25.900 ;
    RECT 0 25.970 0.070 26.880 ;
    RECT 0 26.950 0.070 27.860 ;
    RECT 0 27.930 0.070 28.840 ;
    RECT 0 28.910 0.070 29.820 ;
    RECT 0 29.890 0.070 36.400 ;
    LAYER metal4 ;
    RECT 0 0 10.640 1.400 ;
    RECT 0 35.000 10.640 36.400 ;
    RECT 0.000 1.400 1.260 35.000 ;
    RECT 1.540 1.400 2.380 35.000 ;
    RECT 2.660 1.400 3.500 35.000 ;
    RECT 3.780 1.400 4.620 35.000 ;
    RECT 4.900 1.400 5.740 35.000 ;
    RECT 6.020 1.400 6.860 35.000 ;
    RECT 7.140 1.400 7.980 35.000 ;
    RECT 8.260 1.400 10.640 35.000 ;
    LAYER OVERLAP ;
    RECT 0 0 10.640 36.400 ;
  END
END fakeram45_64x7

END LIBRARY
