module MuxTest_width_1_inputs_4_outputs_16_pipeline_0( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [1:0] io_selects_0_0, // @[:@6.4]
  input  [1:0] io_selects_0_1, // @[:@6.4]
  input  [1:0] io_selects_1_0, // @[:@6.4]
  input  [1:0] io_selects_1_1, // @[:@6.4]
  input  [1:0] io_selects_2_0, // @[:@6.4]
  input  [1:0] io_selects_2_1, // @[:@6.4]
  input  [1:0] io_selects_3_0, // @[:@6.4]
  input  [1:0] io_selects_3_1, // @[:@6.4]
  input  [1:0] io_selects_4_0, // @[:@6.4]
  input  [1:0] io_selects_4_1, // @[:@6.4]
  input  [1:0] io_selects_5_0, // @[:@6.4]
  input  [1:0] io_selects_5_1, // @[:@6.4]
  input  [1:0] io_selects_6_0, // @[:@6.4]
  input  [1:0] io_selects_6_1, // @[:@6.4]
  input  [1:0] io_selects_7_0, // @[:@6.4]
  input  [1:0] io_selects_7_1, // @[:@6.4]
  input  [1:0] io_selects_8_0, // @[:@6.4]
  input  [1:0] io_selects_8_1, // @[:@6.4]
  input  [1:0] io_selects_9_0, // @[:@6.4]
  input  [1:0] io_selects_9_1, // @[:@6.4]
  input  [1:0] io_selects_10_0, // @[:@6.4]
  input  [1:0] io_selects_10_1, // @[:@6.4]
  input  [1:0] io_selects_11_0, // @[:@6.4]
  input  [1:0] io_selects_11_1, // @[:@6.4]
  input  [1:0] io_selects_12_0, // @[:@6.4]
  input  [1:0] io_selects_12_1, // @[:@6.4]
  input  [1:0] io_selects_13_0, // @[:@6.4]
  input  [1:0] io_selects_13_1, // @[:@6.4]
  input  [1:0] io_selects_14_0, // @[:@6.4]
  input  [1:0] io_selects_14_1, // @[:@6.4]
  input  [1:0] io_selects_15_0, // @[:@6.4]
  input  [1:0] io_selects_15_1, // @[:@6.4]
  input  [2:0] io_operation_0, // @[:@6.4]
  input  [2:0] io_operation_1, // @[:@6.4]
  input  [2:0] io_operation_2, // @[:@6.4]
  input  [2:0] io_operation_3, // @[:@6.4]
  input  [2:0] io_operation_4, // @[:@6.4]
  input  [2:0] io_operation_5, // @[:@6.4]
  input  [2:0] io_operation_6, // @[:@6.4]
  input  [2:0] io_operation_7, // @[:@6.4]
  input  [2:0] io_operation_8, // @[:@6.4]
  input  [2:0] io_operation_9, // @[:@6.4]
  input  [2:0] io_operation_10, // @[:@6.4]
  input  [2:0] io_operation_11, // @[:@6.4]
  input  [2:0] io_operation_12, // @[:@6.4]
  input  [2:0] io_operation_13, // @[:@6.4]
  input  [2:0] io_operation_14, // @[:@6.4]
  input  [2:0] io_operation_15, // @[:@6.4]
  input        io_inputs_0, // @[:@6.4]
  input        io_inputs_1, // @[:@6.4]
  input        io_inputs_2, // @[:@6.4]
  input        io_inputs_3, // @[:@6.4]
  output       io_outputs_0, // @[:@6.4]
  output       io_outputs_1, // @[:@6.4]
  output       io_outputs_2, // @[:@6.4]
  output       io_outputs_3, // @[:@6.4]
  output       io_outputs_4, // @[:@6.4]
  output       io_outputs_5, // @[:@6.4]
  output       io_outputs_6, // @[:@6.4]
  output       io_outputs_7, // @[:@6.4]
  output       io_outputs_8, // @[:@6.4]
  output       io_outputs_9, // @[:@6.4]
  output       io_outputs_10, // @[:@6.4]
  output       io_outputs_11, // @[:@6.4]
  output       io_outputs_12, // @[:@6.4]
  output       io_outputs_13, // @[:@6.4]
  output       io_outputs_14, // @[:@6.4]
  output       io_outputs_15 // @[:@6.4]
);
  wire  _GEN_1; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_2; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_3; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_5; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_6; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _GEN_7; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire [1:0] _T_698; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  wire  _T_699; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@9.4]
  wire [1:0] _T_701; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@10.4]
  wire  _T_703; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@11.4]
  wire  _T_704; // @[Mux.scala 46:19:@12.4]
  wire  _T_705; // @[Mux.scala 46:16:@13.4]
  wire  _T_706; // @[Mux.scala 46:19:@14.4]
  wire [1:0] _T_707; // @[Mux.scala 46:16:@15.4]
  wire  _T_708; // @[Mux.scala 46:19:@16.4]
  wire [1:0] _T_709; // @[Mux.scala 46:16:@17.4]
  wire  _T_710; // @[Mux.scala 46:19:@18.4]
  wire [1:0] _T_711; // @[Mux.scala 46:16:@19.4]
  wire  _GEN_9; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_10; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_11; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_13; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_14; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _GEN_15; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire [1:0] _T_715; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  wire  _T_716; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@21.4]
  wire [1:0] _T_718; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@22.4]
  wire  _T_720; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@23.4]
  wire  _T_721; // @[Mux.scala 46:19:@24.4]
  wire  _T_722; // @[Mux.scala 46:16:@25.4]
  wire  _T_723; // @[Mux.scala 46:19:@26.4]
  wire [1:0] _T_724; // @[Mux.scala 46:16:@27.4]
  wire  _T_725; // @[Mux.scala 46:19:@28.4]
  wire [1:0] _T_726; // @[Mux.scala 46:16:@29.4]
  wire  _T_727; // @[Mux.scala 46:19:@30.4]
  wire [1:0] _T_728; // @[Mux.scala 46:16:@31.4]
  wire  _GEN_17; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_18; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_19; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_21; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_22; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _GEN_23; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire [1:0] _T_732; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  wire  _T_733; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@33.4]
  wire [1:0] _T_735; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@34.4]
  wire  _T_737; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@35.4]
  wire  _T_738; // @[Mux.scala 46:19:@36.4]
  wire  _T_739; // @[Mux.scala 46:16:@37.4]
  wire  _T_740; // @[Mux.scala 46:19:@38.4]
  wire [1:0] _T_741; // @[Mux.scala 46:16:@39.4]
  wire  _T_742; // @[Mux.scala 46:19:@40.4]
  wire [1:0] _T_743; // @[Mux.scala 46:16:@41.4]
  wire  _T_744; // @[Mux.scala 46:19:@42.4]
  wire [1:0] _T_745; // @[Mux.scala 46:16:@43.4]
  wire  _GEN_25; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_26; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_27; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_29; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_30; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _GEN_31; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire [1:0] _T_749; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  wire  _T_750; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@45.4]
  wire [1:0] _T_752; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@46.4]
  wire  _T_754; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@47.4]
  wire  _T_755; // @[Mux.scala 46:19:@48.4]
  wire  _T_756; // @[Mux.scala 46:16:@49.4]
  wire  _T_757; // @[Mux.scala 46:19:@50.4]
  wire [1:0] _T_758; // @[Mux.scala 46:16:@51.4]
  wire  _T_759; // @[Mux.scala 46:19:@52.4]
  wire [1:0] _T_760; // @[Mux.scala 46:16:@53.4]
  wire  _T_761; // @[Mux.scala 46:19:@54.4]
  wire [1:0] _T_762; // @[Mux.scala 46:16:@55.4]
  wire  _GEN_33; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_34; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_35; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_37; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_38; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _GEN_39; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire [1:0] _T_766; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  wire  _T_767; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@57.4]
  wire [1:0] _T_769; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@58.4]
  wire  _T_771; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@59.4]
  wire  _T_772; // @[Mux.scala 46:19:@60.4]
  wire  _T_773; // @[Mux.scala 46:16:@61.4]
  wire  _T_774; // @[Mux.scala 46:19:@62.4]
  wire [1:0] _T_775; // @[Mux.scala 46:16:@63.4]
  wire  _T_776; // @[Mux.scala 46:19:@64.4]
  wire [1:0] _T_777; // @[Mux.scala 46:16:@65.4]
  wire  _T_778; // @[Mux.scala 46:19:@66.4]
  wire [1:0] _T_779; // @[Mux.scala 46:16:@67.4]
  wire  _GEN_41; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_42; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_43; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_45; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_46; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _GEN_47; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire [1:0] _T_783; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  wire  _T_784; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@69.4]
  wire [1:0] _T_786; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@70.4]
  wire  _T_788; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@71.4]
  wire  _T_789; // @[Mux.scala 46:19:@72.4]
  wire  _T_790; // @[Mux.scala 46:16:@73.4]
  wire  _T_791; // @[Mux.scala 46:19:@74.4]
  wire [1:0] _T_792; // @[Mux.scala 46:16:@75.4]
  wire  _T_793; // @[Mux.scala 46:19:@76.4]
  wire [1:0] _T_794; // @[Mux.scala 46:16:@77.4]
  wire  _T_795; // @[Mux.scala 46:19:@78.4]
  wire [1:0] _T_796; // @[Mux.scala 46:16:@79.4]
  wire  _GEN_49; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_50; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_51; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_53; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_54; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _GEN_55; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire [1:0] _T_800; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  wire  _T_801; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@81.4]
  wire [1:0] _T_803; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@82.4]
  wire  _T_805; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@83.4]
  wire  _T_806; // @[Mux.scala 46:19:@84.4]
  wire  _T_807; // @[Mux.scala 46:16:@85.4]
  wire  _T_808; // @[Mux.scala 46:19:@86.4]
  wire [1:0] _T_809; // @[Mux.scala 46:16:@87.4]
  wire  _T_810; // @[Mux.scala 46:19:@88.4]
  wire [1:0] _T_811; // @[Mux.scala 46:16:@89.4]
  wire  _T_812; // @[Mux.scala 46:19:@90.4]
  wire [1:0] _T_813; // @[Mux.scala 46:16:@91.4]
  wire  _GEN_57; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_58; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_59; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_61; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_62; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _GEN_63; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire [1:0] _T_817; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  wire  _T_818; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@93.4]
  wire [1:0] _T_820; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@94.4]
  wire  _T_822; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@95.4]
  wire  _T_823; // @[Mux.scala 46:19:@96.4]
  wire  _T_824; // @[Mux.scala 46:16:@97.4]
  wire  _T_825; // @[Mux.scala 46:19:@98.4]
  wire [1:0] _T_826; // @[Mux.scala 46:16:@99.4]
  wire  _T_827; // @[Mux.scala 46:19:@100.4]
  wire [1:0] _T_828; // @[Mux.scala 46:16:@101.4]
  wire  _T_829; // @[Mux.scala 46:19:@102.4]
  wire [1:0] _T_830; // @[Mux.scala 46:16:@103.4]
  wire  _GEN_65; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_66; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_67; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_69; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_70; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _GEN_71; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire [1:0] _T_834; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  wire  _T_835; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@105.4]
  wire [1:0] _T_837; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@106.4]
  wire  _T_839; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@107.4]
  wire  _T_840; // @[Mux.scala 46:19:@108.4]
  wire  _T_841; // @[Mux.scala 46:16:@109.4]
  wire  _T_842; // @[Mux.scala 46:19:@110.4]
  wire [1:0] _T_843; // @[Mux.scala 46:16:@111.4]
  wire  _T_844; // @[Mux.scala 46:19:@112.4]
  wire [1:0] _T_845; // @[Mux.scala 46:16:@113.4]
  wire  _T_846; // @[Mux.scala 46:19:@114.4]
  wire [1:0] _T_847; // @[Mux.scala 46:16:@115.4]
  wire  _GEN_73; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_74; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_75; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_77; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_78; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _GEN_79; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire [1:0] _T_851; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  wire  _T_852; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@117.4]
  wire [1:0] _T_854; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@118.4]
  wire  _T_856; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@119.4]
  wire  _T_857; // @[Mux.scala 46:19:@120.4]
  wire  _T_858; // @[Mux.scala 46:16:@121.4]
  wire  _T_859; // @[Mux.scala 46:19:@122.4]
  wire [1:0] _T_860; // @[Mux.scala 46:16:@123.4]
  wire  _T_861; // @[Mux.scala 46:19:@124.4]
  wire [1:0] _T_862; // @[Mux.scala 46:16:@125.4]
  wire  _T_863; // @[Mux.scala 46:19:@126.4]
  wire [1:0] _T_864; // @[Mux.scala 46:16:@127.4]
  wire  _GEN_81; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_82; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_83; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_85; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_86; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _GEN_87; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire [1:0] _T_868; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  wire  _T_869; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@129.4]
  wire [1:0] _T_871; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@130.4]
  wire  _T_873; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@131.4]
  wire  _T_874; // @[Mux.scala 46:19:@132.4]
  wire  _T_875; // @[Mux.scala 46:16:@133.4]
  wire  _T_876; // @[Mux.scala 46:19:@134.4]
  wire [1:0] _T_877; // @[Mux.scala 46:16:@135.4]
  wire  _T_878; // @[Mux.scala 46:19:@136.4]
  wire [1:0] _T_879; // @[Mux.scala 46:16:@137.4]
  wire  _T_880; // @[Mux.scala 46:19:@138.4]
  wire [1:0] _T_881; // @[Mux.scala 46:16:@139.4]
  wire  _GEN_89; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_90; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_91; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_93; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_94; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _GEN_95; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire [1:0] _T_885; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  wire  _T_886; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@141.4]
  wire [1:0] _T_888; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@142.4]
  wire  _T_890; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@143.4]
  wire  _T_891; // @[Mux.scala 46:19:@144.4]
  wire  _T_892; // @[Mux.scala 46:16:@145.4]
  wire  _T_893; // @[Mux.scala 46:19:@146.4]
  wire [1:0] _T_894; // @[Mux.scala 46:16:@147.4]
  wire  _T_895; // @[Mux.scala 46:19:@148.4]
  wire [1:0] _T_896; // @[Mux.scala 46:16:@149.4]
  wire  _T_897; // @[Mux.scala 46:19:@150.4]
  wire [1:0] _T_898; // @[Mux.scala 46:16:@151.4]
  wire  _GEN_97; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_98; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_99; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_101; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_102; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _GEN_103; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire [1:0] _T_902; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  wire  _T_903; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@153.4]
  wire [1:0] _T_905; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@154.4]
  wire  _T_907; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@155.4]
  wire  _T_908; // @[Mux.scala 46:19:@156.4]
  wire  _T_909; // @[Mux.scala 46:16:@157.4]
  wire  _T_910; // @[Mux.scala 46:19:@158.4]
  wire [1:0] _T_911; // @[Mux.scala 46:16:@159.4]
  wire  _T_912; // @[Mux.scala 46:19:@160.4]
  wire [1:0] _T_913; // @[Mux.scala 46:16:@161.4]
  wire  _T_914; // @[Mux.scala 46:19:@162.4]
  wire [1:0] _T_915; // @[Mux.scala 46:16:@163.4]
  wire  _GEN_105; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_106; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_107; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_109; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_110; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _GEN_111; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire [1:0] _T_919; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  wire  _T_920; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@165.4]
  wire [1:0] _T_922; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@166.4]
  wire  _T_924; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@167.4]
  wire  _T_925; // @[Mux.scala 46:19:@168.4]
  wire  _T_926; // @[Mux.scala 46:16:@169.4]
  wire  _T_927; // @[Mux.scala 46:19:@170.4]
  wire [1:0] _T_928; // @[Mux.scala 46:16:@171.4]
  wire  _T_929; // @[Mux.scala 46:19:@172.4]
  wire [1:0] _T_930; // @[Mux.scala 46:16:@173.4]
  wire  _T_931; // @[Mux.scala 46:19:@174.4]
  wire [1:0] _T_932; // @[Mux.scala 46:16:@175.4]
  wire  _GEN_113; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_114; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_115; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_117; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_118; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _GEN_119; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire [1:0] _T_936; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  wire  _T_937; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@177.4]
  wire [1:0] _T_939; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@178.4]
  wire  _T_941; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@179.4]
  wire  _T_942; // @[Mux.scala 46:19:@180.4]
  wire  _T_943; // @[Mux.scala 46:16:@181.4]
  wire  _T_944; // @[Mux.scala 46:19:@182.4]
  wire [1:0] _T_945; // @[Mux.scala 46:16:@183.4]
  wire  _T_946; // @[Mux.scala 46:19:@184.4]
  wire [1:0] _T_947; // @[Mux.scala 46:16:@185.4]
  wire  _T_948; // @[Mux.scala 46:19:@186.4]
  wire [1:0] _T_949; // @[Mux.scala 46:16:@187.4]
  wire  _GEN_121; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_122; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_123; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_125; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_126; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _GEN_127; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire [1:0] _T_953; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  wire  _T_954; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@189.4]
  wire [1:0] _T_956; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@190.4]
  wire  _T_958; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@191.4]
  wire  _T_959; // @[Mux.scala 46:19:@192.4]
  wire  _T_960; // @[Mux.scala 46:16:@193.4]
  wire  _T_961; // @[Mux.scala 46:19:@194.4]
  wire [1:0] _T_962; // @[Mux.scala 46:16:@195.4]
  wire  _T_963; // @[Mux.scala 46:19:@196.4]
  wire [1:0] _T_964; // @[Mux.scala 46:16:@197.4]
  wire  _T_965; // @[Mux.scala 46:19:@198.4]
  wire [1:0] _T_966; // @[Mux.scala 46:16:@199.4]
  assign _GEN_1 = 2'h1 == io_selects_0_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_2 = 2'h2 == io_selects_0_0 ? io_inputs_2 : _GEN_1; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_3 = 2'h3 == io_selects_0_0 ? io_inputs_3 : _GEN_2; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_5 = 2'h1 == io_selects_0_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_6 = 2'h2 == io_selects_0_1 ? io_inputs_2 : _GEN_5; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _GEN_7 = 2'h3 == io_selects_0_1 ? io_inputs_3 : _GEN_6; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _T_698 = _GEN_3 + _GEN_7; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@8.4]
  assign _T_699 = _GEN_3 + _GEN_7; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@9.4]
  assign _T_701 = _GEN_3 * _GEN_7; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@10.4]
  assign _T_703 = _GEN_3 / _GEN_7; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@11.4]
  assign _T_704 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_705 = _T_704 ? _T_703 : 1'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_706 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_707 = _T_706 ? _T_701 : {{1'd0}, _T_705}; // @[Mux.scala 46:16:@15.4]
  assign _T_708 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_709 = _T_708 ? {{1'd0}, _T_699} : _T_707; // @[Mux.scala 46:16:@17.4]
  assign _T_710 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _T_711 = _T_710 ? {{1'd0}, _GEN_3} : _T_709; // @[Mux.scala 46:16:@19.4]
  assign _GEN_9 = 2'h1 == io_selects_1_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_10 = 2'h2 == io_selects_1_0 ? io_inputs_2 : _GEN_9; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_11 = 2'h3 == io_selects_1_0 ? io_inputs_3 : _GEN_10; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_13 = 2'h1 == io_selects_1_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_14 = 2'h2 == io_selects_1_1 ? io_inputs_2 : _GEN_13; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _GEN_15 = 2'h3 == io_selects_1_1 ? io_inputs_3 : _GEN_14; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _T_715 = _GEN_11 + _GEN_15; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@20.4]
  assign _T_716 = _GEN_11 + _GEN_15; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@21.4]
  assign _T_718 = _GEN_11 * _GEN_15; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@22.4]
  assign _T_720 = _GEN_11 / _GEN_15; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@23.4]
  assign _T_721 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_722 = _T_721 ? _T_720 : 1'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_723 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_724 = _T_723 ? _T_718 : {{1'd0}, _T_722}; // @[Mux.scala 46:16:@27.4]
  assign _T_725 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_726 = _T_725 ? {{1'd0}, _T_716} : _T_724; // @[Mux.scala 46:16:@29.4]
  assign _T_727 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _T_728 = _T_727 ? {{1'd0}, _GEN_11} : _T_726; // @[Mux.scala 46:16:@31.4]
  assign _GEN_17 = 2'h1 == io_selects_2_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_18 = 2'h2 == io_selects_2_0 ? io_inputs_2 : _GEN_17; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_19 = 2'h3 == io_selects_2_0 ? io_inputs_3 : _GEN_18; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_21 = 2'h1 == io_selects_2_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_22 = 2'h2 == io_selects_2_1 ? io_inputs_2 : _GEN_21; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _GEN_23 = 2'h3 == io_selects_2_1 ? io_inputs_3 : _GEN_22; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _T_732 = _GEN_19 + _GEN_23; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@32.4]
  assign _T_733 = _GEN_19 + _GEN_23; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@33.4]
  assign _T_735 = _GEN_19 * _GEN_23; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@34.4]
  assign _T_737 = _GEN_19 / _GEN_23; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@35.4]
  assign _T_738 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_739 = _T_738 ? _T_737 : 1'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_740 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_741 = _T_740 ? _T_735 : {{1'd0}, _T_739}; // @[Mux.scala 46:16:@39.4]
  assign _T_742 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_743 = _T_742 ? {{1'd0}, _T_733} : _T_741; // @[Mux.scala 46:16:@41.4]
  assign _T_744 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _T_745 = _T_744 ? {{1'd0}, _GEN_19} : _T_743; // @[Mux.scala 46:16:@43.4]
  assign _GEN_25 = 2'h1 == io_selects_3_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_26 = 2'h2 == io_selects_3_0 ? io_inputs_2 : _GEN_25; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_27 = 2'h3 == io_selects_3_0 ? io_inputs_3 : _GEN_26; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_29 = 2'h1 == io_selects_3_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_30 = 2'h2 == io_selects_3_1 ? io_inputs_2 : _GEN_29; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _GEN_31 = 2'h3 == io_selects_3_1 ? io_inputs_3 : _GEN_30; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _T_749 = _GEN_27 + _GEN_31; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@44.4]
  assign _T_750 = _GEN_27 + _GEN_31; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@45.4]
  assign _T_752 = _GEN_27 * _GEN_31; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@46.4]
  assign _T_754 = _GEN_27 / _GEN_31; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@47.4]
  assign _T_755 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_756 = _T_755 ? _T_754 : 1'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_757 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_758 = _T_757 ? _T_752 : {{1'd0}, _T_756}; // @[Mux.scala 46:16:@51.4]
  assign _T_759 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_760 = _T_759 ? {{1'd0}, _T_750} : _T_758; // @[Mux.scala 46:16:@53.4]
  assign _T_761 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _T_762 = _T_761 ? {{1'd0}, _GEN_27} : _T_760; // @[Mux.scala 46:16:@55.4]
  assign _GEN_33 = 2'h1 == io_selects_4_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_34 = 2'h2 == io_selects_4_0 ? io_inputs_2 : _GEN_33; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_35 = 2'h3 == io_selects_4_0 ? io_inputs_3 : _GEN_34; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_37 = 2'h1 == io_selects_4_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_38 = 2'h2 == io_selects_4_1 ? io_inputs_2 : _GEN_37; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _GEN_39 = 2'h3 == io_selects_4_1 ? io_inputs_3 : _GEN_38; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _T_766 = _GEN_35 + _GEN_39; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@56.4]
  assign _T_767 = _GEN_35 + _GEN_39; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@57.4]
  assign _T_769 = _GEN_35 * _GEN_39; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@58.4]
  assign _T_771 = _GEN_35 / _GEN_39; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@59.4]
  assign _T_772 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_773 = _T_772 ? _T_771 : 1'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_774 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_775 = _T_774 ? _T_769 : {{1'd0}, _T_773}; // @[Mux.scala 46:16:@63.4]
  assign _T_776 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_777 = _T_776 ? {{1'd0}, _T_767} : _T_775; // @[Mux.scala 46:16:@65.4]
  assign _T_778 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _T_779 = _T_778 ? {{1'd0}, _GEN_35} : _T_777; // @[Mux.scala 46:16:@67.4]
  assign _GEN_41 = 2'h1 == io_selects_5_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_42 = 2'h2 == io_selects_5_0 ? io_inputs_2 : _GEN_41; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_43 = 2'h3 == io_selects_5_0 ? io_inputs_3 : _GEN_42; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_45 = 2'h1 == io_selects_5_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_46 = 2'h2 == io_selects_5_1 ? io_inputs_2 : _GEN_45; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _GEN_47 = 2'h3 == io_selects_5_1 ? io_inputs_3 : _GEN_46; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _T_783 = _GEN_43 + _GEN_47; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@68.4]
  assign _T_784 = _GEN_43 + _GEN_47; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@69.4]
  assign _T_786 = _GEN_43 * _GEN_47; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@70.4]
  assign _T_788 = _GEN_43 / _GEN_47; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@71.4]
  assign _T_789 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_790 = _T_789 ? _T_788 : 1'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_791 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_792 = _T_791 ? _T_786 : {{1'd0}, _T_790}; // @[Mux.scala 46:16:@75.4]
  assign _T_793 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_794 = _T_793 ? {{1'd0}, _T_784} : _T_792; // @[Mux.scala 46:16:@77.4]
  assign _T_795 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _T_796 = _T_795 ? {{1'd0}, _GEN_43} : _T_794; // @[Mux.scala 46:16:@79.4]
  assign _GEN_49 = 2'h1 == io_selects_6_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_50 = 2'h2 == io_selects_6_0 ? io_inputs_2 : _GEN_49; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_51 = 2'h3 == io_selects_6_0 ? io_inputs_3 : _GEN_50; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_53 = 2'h1 == io_selects_6_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_54 = 2'h2 == io_selects_6_1 ? io_inputs_2 : _GEN_53; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _GEN_55 = 2'h3 == io_selects_6_1 ? io_inputs_3 : _GEN_54; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _T_800 = _GEN_51 + _GEN_55; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@80.4]
  assign _T_801 = _GEN_51 + _GEN_55; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@81.4]
  assign _T_803 = _GEN_51 * _GEN_55; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@82.4]
  assign _T_805 = _GEN_51 / _GEN_55; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@83.4]
  assign _T_806 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_807 = _T_806 ? _T_805 : 1'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_808 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_809 = _T_808 ? _T_803 : {{1'd0}, _T_807}; // @[Mux.scala 46:16:@87.4]
  assign _T_810 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_811 = _T_810 ? {{1'd0}, _T_801} : _T_809; // @[Mux.scala 46:16:@89.4]
  assign _T_812 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _T_813 = _T_812 ? {{1'd0}, _GEN_51} : _T_811; // @[Mux.scala 46:16:@91.4]
  assign _GEN_57 = 2'h1 == io_selects_7_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_58 = 2'h2 == io_selects_7_0 ? io_inputs_2 : _GEN_57; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_59 = 2'h3 == io_selects_7_0 ? io_inputs_3 : _GEN_58; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_61 = 2'h1 == io_selects_7_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_62 = 2'h2 == io_selects_7_1 ? io_inputs_2 : _GEN_61; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _GEN_63 = 2'h3 == io_selects_7_1 ? io_inputs_3 : _GEN_62; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _T_817 = _GEN_59 + _GEN_63; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@92.4]
  assign _T_818 = _GEN_59 + _GEN_63; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@93.4]
  assign _T_820 = _GEN_59 * _GEN_63; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@94.4]
  assign _T_822 = _GEN_59 / _GEN_63; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@95.4]
  assign _T_823 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_824 = _T_823 ? _T_822 : 1'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_825 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_826 = _T_825 ? _T_820 : {{1'd0}, _T_824}; // @[Mux.scala 46:16:@99.4]
  assign _T_827 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_828 = _T_827 ? {{1'd0}, _T_818} : _T_826; // @[Mux.scala 46:16:@101.4]
  assign _T_829 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign _T_830 = _T_829 ? {{1'd0}, _GEN_59} : _T_828; // @[Mux.scala 46:16:@103.4]
  assign _GEN_65 = 2'h1 == io_selects_8_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_66 = 2'h2 == io_selects_8_0 ? io_inputs_2 : _GEN_65; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_67 = 2'h3 == io_selects_8_0 ? io_inputs_3 : _GEN_66; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_69 = 2'h1 == io_selects_8_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_70 = 2'h2 == io_selects_8_1 ? io_inputs_2 : _GEN_69; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _GEN_71 = 2'h3 == io_selects_8_1 ? io_inputs_3 : _GEN_70; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _T_834 = _GEN_67 + _GEN_71; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@104.4]
  assign _T_835 = _GEN_67 + _GEN_71; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@105.4]
  assign _T_837 = _GEN_67 * _GEN_71; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@106.4]
  assign _T_839 = _GEN_67 / _GEN_71; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@107.4]
  assign _T_840 = 3'h3 == io_operation_8; // @[Mux.scala 46:19:@108.4]
  assign _T_841 = _T_840 ? _T_839 : 1'h0; // @[Mux.scala 46:16:@109.4]
  assign _T_842 = 3'h2 == io_operation_8; // @[Mux.scala 46:19:@110.4]
  assign _T_843 = _T_842 ? _T_837 : {{1'd0}, _T_841}; // @[Mux.scala 46:16:@111.4]
  assign _T_844 = 3'h1 == io_operation_8; // @[Mux.scala 46:19:@112.4]
  assign _T_845 = _T_844 ? {{1'd0}, _T_835} : _T_843; // @[Mux.scala 46:16:@113.4]
  assign _T_846 = 3'h0 == io_operation_8; // @[Mux.scala 46:19:@114.4]
  assign _T_847 = _T_846 ? {{1'd0}, _GEN_67} : _T_845; // @[Mux.scala 46:16:@115.4]
  assign _GEN_73 = 2'h1 == io_selects_9_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_74 = 2'h2 == io_selects_9_0 ? io_inputs_2 : _GEN_73; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_75 = 2'h3 == io_selects_9_0 ? io_inputs_3 : _GEN_74; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_77 = 2'h1 == io_selects_9_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_78 = 2'h2 == io_selects_9_1 ? io_inputs_2 : _GEN_77; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _GEN_79 = 2'h3 == io_selects_9_1 ? io_inputs_3 : _GEN_78; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _T_851 = _GEN_75 + _GEN_79; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@116.4]
  assign _T_852 = _GEN_75 + _GEN_79; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@117.4]
  assign _T_854 = _GEN_75 * _GEN_79; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@118.4]
  assign _T_856 = _GEN_75 / _GEN_79; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@119.4]
  assign _T_857 = 3'h3 == io_operation_9; // @[Mux.scala 46:19:@120.4]
  assign _T_858 = _T_857 ? _T_856 : 1'h0; // @[Mux.scala 46:16:@121.4]
  assign _T_859 = 3'h2 == io_operation_9; // @[Mux.scala 46:19:@122.4]
  assign _T_860 = _T_859 ? _T_854 : {{1'd0}, _T_858}; // @[Mux.scala 46:16:@123.4]
  assign _T_861 = 3'h1 == io_operation_9; // @[Mux.scala 46:19:@124.4]
  assign _T_862 = _T_861 ? {{1'd0}, _T_852} : _T_860; // @[Mux.scala 46:16:@125.4]
  assign _T_863 = 3'h0 == io_operation_9; // @[Mux.scala 46:19:@126.4]
  assign _T_864 = _T_863 ? {{1'd0}, _GEN_75} : _T_862; // @[Mux.scala 46:16:@127.4]
  assign _GEN_81 = 2'h1 == io_selects_10_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_82 = 2'h2 == io_selects_10_0 ? io_inputs_2 : _GEN_81; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_83 = 2'h3 == io_selects_10_0 ? io_inputs_3 : _GEN_82; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_85 = 2'h1 == io_selects_10_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_86 = 2'h2 == io_selects_10_1 ? io_inputs_2 : _GEN_85; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _GEN_87 = 2'h3 == io_selects_10_1 ? io_inputs_3 : _GEN_86; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _T_868 = _GEN_83 + _GEN_87; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@128.4]
  assign _T_869 = _GEN_83 + _GEN_87; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@129.4]
  assign _T_871 = _GEN_83 * _GEN_87; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@130.4]
  assign _T_873 = _GEN_83 / _GEN_87; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@131.4]
  assign _T_874 = 3'h3 == io_operation_10; // @[Mux.scala 46:19:@132.4]
  assign _T_875 = _T_874 ? _T_873 : 1'h0; // @[Mux.scala 46:16:@133.4]
  assign _T_876 = 3'h2 == io_operation_10; // @[Mux.scala 46:19:@134.4]
  assign _T_877 = _T_876 ? _T_871 : {{1'd0}, _T_875}; // @[Mux.scala 46:16:@135.4]
  assign _T_878 = 3'h1 == io_operation_10; // @[Mux.scala 46:19:@136.4]
  assign _T_879 = _T_878 ? {{1'd0}, _T_869} : _T_877; // @[Mux.scala 46:16:@137.4]
  assign _T_880 = 3'h0 == io_operation_10; // @[Mux.scala 46:19:@138.4]
  assign _T_881 = _T_880 ? {{1'd0}, _GEN_83} : _T_879; // @[Mux.scala 46:16:@139.4]
  assign _GEN_89 = 2'h1 == io_selects_11_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_90 = 2'h2 == io_selects_11_0 ? io_inputs_2 : _GEN_89; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_91 = 2'h3 == io_selects_11_0 ? io_inputs_3 : _GEN_90; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_93 = 2'h1 == io_selects_11_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_94 = 2'h2 == io_selects_11_1 ? io_inputs_2 : _GEN_93; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _GEN_95 = 2'h3 == io_selects_11_1 ? io_inputs_3 : _GEN_94; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _T_885 = _GEN_91 + _GEN_95; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@140.4]
  assign _T_886 = _GEN_91 + _GEN_95; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@141.4]
  assign _T_888 = _GEN_91 * _GEN_95; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@142.4]
  assign _T_890 = _GEN_91 / _GEN_95; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@143.4]
  assign _T_891 = 3'h3 == io_operation_11; // @[Mux.scala 46:19:@144.4]
  assign _T_892 = _T_891 ? _T_890 : 1'h0; // @[Mux.scala 46:16:@145.4]
  assign _T_893 = 3'h2 == io_operation_11; // @[Mux.scala 46:19:@146.4]
  assign _T_894 = _T_893 ? _T_888 : {{1'd0}, _T_892}; // @[Mux.scala 46:16:@147.4]
  assign _T_895 = 3'h1 == io_operation_11; // @[Mux.scala 46:19:@148.4]
  assign _T_896 = _T_895 ? {{1'd0}, _T_886} : _T_894; // @[Mux.scala 46:16:@149.4]
  assign _T_897 = 3'h0 == io_operation_11; // @[Mux.scala 46:19:@150.4]
  assign _T_898 = _T_897 ? {{1'd0}, _GEN_91} : _T_896; // @[Mux.scala 46:16:@151.4]
  assign _GEN_97 = 2'h1 == io_selects_12_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_98 = 2'h2 == io_selects_12_0 ? io_inputs_2 : _GEN_97; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_99 = 2'h3 == io_selects_12_0 ? io_inputs_3 : _GEN_98; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_101 = 2'h1 == io_selects_12_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_102 = 2'h2 == io_selects_12_1 ? io_inputs_2 : _GEN_101; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _GEN_103 = 2'h3 == io_selects_12_1 ? io_inputs_3 : _GEN_102; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _T_902 = _GEN_99 + _GEN_103; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@152.4]
  assign _T_903 = _GEN_99 + _GEN_103; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@153.4]
  assign _T_905 = _GEN_99 * _GEN_103; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@154.4]
  assign _T_907 = _GEN_99 / _GEN_103; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@155.4]
  assign _T_908 = 3'h3 == io_operation_12; // @[Mux.scala 46:19:@156.4]
  assign _T_909 = _T_908 ? _T_907 : 1'h0; // @[Mux.scala 46:16:@157.4]
  assign _T_910 = 3'h2 == io_operation_12; // @[Mux.scala 46:19:@158.4]
  assign _T_911 = _T_910 ? _T_905 : {{1'd0}, _T_909}; // @[Mux.scala 46:16:@159.4]
  assign _T_912 = 3'h1 == io_operation_12; // @[Mux.scala 46:19:@160.4]
  assign _T_913 = _T_912 ? {{1'd0}, _T_903} : _T_911; // @[Mux.scala 46:16:@161.4]
  assign _T_914 = 3'h0 == io_operation_12; // @[Mux.scala 46:19:@162.4]
  assign _T_915 = _T_914 ? {{1'd0}, _GEN_99} : _T_913; // @[Mux.scala 46:16:@163.4]
  assign _GEN_105 = 2'h1 == io_selects_13_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_106 = 2'h2 == io_selects_13_0 ? io_inputs_2 : _GEN_105; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_107 = 2'h3 == io_selects_13_0 ? io_inputs_3 : _GEN_106; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_109 = 2'h1 == io_selects_13_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_110 = 2'h2 == io_selects_13_1 ? io_inputs_2 : _GEN_109; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _GEN_111 = 2'h3 == io_selects_13_1 ? io_inputs_3 : _GEN_110; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _T_919 = _GEN_107 + _GEN_111; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@164.4]
  assign _T_920 = _GEN_107 + _GEN_111; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@165.4]
  assign _T_922 = _GEN_107 * _GEN_111; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@166.4]
  assign _T_924 = _GEN_107 / _GEN_111; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@167.4]
  assign _T_925 = 3'h3 == io_operation_13; // @[Mux.scala 46:19:@168.4]
  assign _T_926 = _T_925 ? _T_924 : 1'h0; // @[Mux.scala 46:16:@169.4]
  assign _T_927 = 3'h2 == io_operation_13; // @[Mux.scala 46:19:@170.4]
  assign _T_928 = _T_927 ? _T_922 : {{1'd0}, _T_926}; // @[Mux.scala 46:16:@171.4]
  assign _T_929 = 3'h1 == io_operation_13; // @[Mux.scala 46:19:@172.4]
  assign _T_930 = _T_929 ? {{1'd0}, _T_920} : _T_928; // @[Mux.scala 46:16:@173.4]
  assign _T_931 = 3'h0 == io_operation_13; // @[Mux.scala 46:19:@174.4]
  assign _T_932 = _T_931 ? {{1'd0}, _GEN_107} : _T_930; // @[Mux.scala 46:16:@175.4]
  assign _GEN_113 = 2'h1 == io_selects_14_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_114 = 2'h2 == io_selects_14_0 ? io_inputs_2 : _GEN_113; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_115 = 2'h3 == io_selects_14_0 ? io_inputs_3 : _GEN_114; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_117 = 2'h1 == io_selects_14_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_118 = 2'h2 == io_selects_14_1 ? io_inputs_2 : _GEN_117; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _GEN_119 = 2'h3 == io_selects_14_1 ? io_inputs_3 : _GEN_118; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _T_936 = _GEN_115 + _GEN_119; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@176.4]
  assign _T_937 = _GEN_115 + _GEN_119; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@177.4]
  assign _T_939 = _GEN_115 * _GEN_119; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@178.4]
  assign _T_941 = _GEN_115 / _GEN_119; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@179.4]
  assign _T_942 = 3'h3 == io_operation_14; // @[Mux.scala 46:19:@180.4]
  assign _T_943 = _T_942 ? _T_941 : 1'h0; // @[Mux.scala 46:16:@181.4]
  assign _T_944 = 3'h2 == io_operation_14; // @[Mux.scala 46:19:@182.4]
  assign _T_945 = _T_944 ? _T_939 : {{1'd0}, _T_943}; // @[Mux.scala 46:16:@183.4]
  assign _T_946 = 3'h1 == io_operation_14; // @[Mux.scala 46:19:@184.4]
  assign _T_947 = _T_946 ? {{1'd0}, _T_937} : _T_945; // @[Mux.scala 46:16:@185.4]
  assign _T_948 = 3'h0 == io_operation_14; // @[Mux.scala 46:19:@186.4]
  assign _T_949 = _T_948 ? {{1'd0}, _GEN_115} : _T_947; // @[Mux.scala 46:16:@187.4]
  assign _GEN_121 = 2'h1 == io_selects_15_0 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_122 = 2'h2 == io_selects_15_0 ? io_inputs_2 : _GEN_121; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_123 = 2'h3 == io_selects_15_0 ? io_inputs_3 : _GEN_122; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_125 = 2'h1 == io_selects_15_1 ? io_inputs_1 : io_inputs_0; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_126 = 2'h2 == io_selects_15_1 ? io_inputs_2 : _GEN_125; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _GEN_127 = 2'h3 == io_selects_15_1 ? io_inputs_3 : _GEN_126; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _T_953 = _GEN_123 + _GEN_127; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@188.4]
  assign _T_954 = _GEN_123 + _GEN_127; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 32:53:@189.4]
  assign _T_956 = _GEN_123 * _GEN_127; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 33:58:@190.4]
  assign _T_958 = _GEN_123 / _GEN_127; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 34:56:@191.4]
  assign _T_959 = 3'h3 == io_operation_15; // @[Mux.scala 46:19:@192.4]
  assign _T_960 = _T_959 ? _T_958 : 1'h0; // @[Mux.scala 46:16:@193.4]
  assign _T_961 = 3'h2 == io_operation_15; // @[Mux.scala 46:19:@194.4]
  assign _T_962 = _T_961 ? _T_956 : {{1'd0}, _T_960}; // @[Mux.scala 46:16:@195.4]
  assign _T_963 = 3'h1 == io_operation_15; // @[Mux.scala 46:19:@196.4]
  assign _T_964 = _T_963 ? {{1'd0}, _T_954} : _T_962; // @[Mux.scala 46:16:@197.4]
  assign _T_965 = 3'h0 == io_operation_15; // @[Mux.scala 46:19:@198.4]
  assign _T_966 = _T_965 ? {{1'd0}, _GEN_123} : _T_964; // @[Mux.scala 46:16:@199.4]
  assign io_outputs_0 = _T_711[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@200.4]
  assign io_outputs_1 = _T_728[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@201.4]
  assign io_outputs_2 = _T_745[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@202.4]
  assign io_outputs_3 = _T_762[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@203.4]
  assign io_outputs_4 = _T_779[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@204.4]
  assign io_outputs_5 = _T_796[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@205.4]
  assign io_outputs_6 = _T_813[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@206.4]
  assign io_outputs_7 = _T_830[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@207.4]
  assign io_outputs_8 = _T_847[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@208.4]
  assign io_outputs_9 = _T_864[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@209.4]
  assign io_outputs_10 = _T_881[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@210.4]
  assign io_outputs_11 = _T_898[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@211.4]
  assign io_outputs_12 = _T_915[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@212.4]
  assign io_outputs_13 = _T_932[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@213.4]
  assign io_outputs_14 = _T_949[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@214.4]
  assign io_outputs_15 = _T_966[0]; // @[MuxTest_width_1_inputs_4_outputs_16_pipeline_0s.scala 23:14:@215.4]
endmodule
