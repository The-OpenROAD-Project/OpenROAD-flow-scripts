VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_64x22
  FOREIGN fakeram_64x22 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 3.040 BY 16.800 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.048 0.024 0.072 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.336 0.024 0.360 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.624 0.024 0.648 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.912 0.024 0.936 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.200 0.024 1.224 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.488 0.024 1.512 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.776 0.024 1.800 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.064 0.024 2.088 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.352 0.024 2.376 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.640 0.024 2.664 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.928 0.024 2.952 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.216 0.024 3.240 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.504 0.024 3.528 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.792 0.024 3.816 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.080 0.024 4.104 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.368 0.024 4.392 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.656 0.024 4.680 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.944 0.024 4.968 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.232 0.024 5.256 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.520 0.024 5.544 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.808 0.024 5.832 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.096 0.024 6.120 ;
    END
  END rd_out[21]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.432 0.024 6.456 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.720 0.024 6.744 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.008 0.024 7.032 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.296 0.024 7.320 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.584 0.024 7.608 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.872 0.024 7.896 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.160 0.024 8.184 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.448 0.024 8.472 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 8.736 0.024 8.760 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.024 0.024 9.048 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.312 0.024 9.336 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.600 0.024 9.624 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 9.888 0.024 9.912 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.176 0.024 10.200 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.464 0.024 10.488 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 10.752 0.024 10.776 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.040 0.024 11.064 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.328 0.024 11.352 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.616 0.024 11.640 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 11.904 0.024 11.928 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.192 0.024 12.216 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.480 0.024 12.504 ;
    END
  END wd_in[21]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 12.816 0.024 12.840 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.104 0.024 13.128 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.392 0.024 13.416 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.680 0.024 13.704 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 13.968 0.024 13.992 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.256 0.024 14.280 ;
    END
  END addr_in[5]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.592 0.024 14.616 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 14.880 0.024 14.904 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 15.168 0.024 15.192 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.000 2.992 0.096 ;
      RECT 0.048 0.768 2.992 0.864 ;
      RECT 0.048 1.536 2.992 1.632 ;
      RECT 0.048 2.304 2.992 2.400 ;
      RECT 0.048 3.072 2.992 3.168 ;
      RECT 0.048 3.840 2.992 3.936 ;
      RECT 0.048 4.608 2.992 4.704 ;
      RECT 0.048 5.376 2.992 5.472 ;
      RECT 0.048 6.144 2.992 6.240 ;
      RECT 0.048 6.912 2.992 7.008 ;
      RECT 0.048 7.680 2.992 7.776 ;
      RECT 0.048 8.448 2.992 8.544 ;
      RECT 0.048 9.216 2.992 9.312 ;
      RECT 0.048 9.984 2.992 10.080 ;
      RECT 0.048 10.752 2.992 10.848 ;
      RECT 0.048 11.520 2.992 11.616 ;
      RECT 0.048 12.288 2.992 12.384 ;
      RECT 0.048 13.056 2.992 13.152 ;
      RECT 0.048 13.824 2.992 13.920 ;
      RECT 0.048 14.592 2.992 14.688 ;
      RECT 0.048 15.360 2.992 15.456 ;
      RECT 0.048 16.128 2.992 16.224 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.384 2.992 0.480 ;
      RECT 0.048 1.152 2.992 1.248 ;
      RECT 0.048 1.920 2.992 2.016 ;
      RECT 0.048 2.688 2.992 2.784 ;
      RECT 0.048 3.456 2.992 3.552 ;
      RECT 0.048 4.224 2.992 4.320 ;
      RECT 0.048 4.992 2.992 5.088 ;
      RECT 0.048 5.760 2.992 5.856 ;
      RECT 0.048 6.528 2.992 6.624 ;
      RECT 0.048 7.296 2.992 7.392 ;
      RECT 0.048 8.064 2.992 8.160 ;
      RECT 0.048 8.832 2.992 8.928 ;
      RECT 0.048 9.600 2.992 9.696 ;
      RECT 0.048 10.368 2.992 10.464 ;
      RECT 0.048 11.136 2.992 11.232 ;
      RECT 0.048 11.904 2.992 12.000 ;
      RECT 0.048 12.672 2.992 12.768 ;
      RECT 0.048 13.440 2.992 13.536 ;
      RECT 0.048 14.208 2.992 14.304 ;
      RECT 0.048 14.976 2.992 15.072 ;
      RECT 0.048 15.744 2.992 15.840 ;
      RECT 0.048 16.512 2.992 16.608 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 3.040 16.800 ;
    LAYER M2 ;
    RECT 0 0 3.040 16.800 ;
    LAYER M3 ;
    RECT 0 0 3.040 16.800 ;
    LAYER M4 ;
    RECT 0.024 0 0.048 16.800 ;
    RECT 2.992 0 3.040 16.800 ;
    RECT 0.048 0.000 2.992 0.000 ;
    RECT 0.048 0.096 2.992 0.384 ;
    RECT 0.048 0.480 2.992 0.768 ;
    RECT 0.048 0.864 2.992 1.152 ;
    RECT 0.048 1.248 2.992 1.536 ;
    RECT 0.048 1.632 2.992 1.920 ;
    RECT 0.048 2.016 2.992 2.304 ;
    RECT 0.048 2.400 2.992 2.688 ;
    RECT 0.048 2.784 2.992 3.072 ;
    RECT 0.048 3.168 2.992 3.456 ;
    RECT 0.048 3.552 2.992 3.840 ;
    RECT 0.048 3.936 2.992 4.224 ;
    RECT 0.048 4.320 2.992 4.608 ;
    RECT 0.048 4.704 2.992 4.992 ;
    RECT 0.048 5.088 2.992 5.376 ;
    RECT 0.048 5.472 2.992 5.760 ;
    RECT 0.048 5.856 2.992 6.144 ;
    RECT 0.048 6.240 2.992 6.528 ;
    RECT 0.048 6.624 2.992 6.912 ;
    RECT 0.048 7.008 2.992 7.296 ;
    RECT 0.048 7.392 2.992 7.680 ;
    RECT 0.048 7.776 2.992 8.064 ;
    RECT 0.048 8.160 2.992 8.448 ;
    RECT 0.048 8.544 2.992 8.832 ;
    RECT 0.048 8.928 2.992 9.216 ;
    RECT 0.048 9.312 2.992 9.600 ;
    RECT 0.048 9.696 2.992 9.984 ;
    RECT 0.048 10.080 2.992 10.368 ;
    RECT 0.048 10.464 2.992 10.752 ;
    RECT 0.048 10.848 2.992 11.136 ;
    RECT 0.048 11.232 2.992 11.520 ;
    RECT 0.048 11.616 2.992 11.904 ;
    RECT 0.048 12.000 2.992 12.288 ;
    RECT 0.048 12.384 2.992 12.672 ;
    RECT 0.048 12.768 2.992 13.056 ;
    RECT 0.048 13.152 2.992 13.440 ;
    RECT 0.048 13.536 2.992 13.824 ;
    RECT 0.048 13.920 2.992 14.208 ;
    RECT 0.048 14.304 2.992 14.592 ;
    RECT 0.048 14.688 2.992 14.976 ;
    RECT 0.048 15.072 2.992 15.360 ;
    RECT 0.048 15.456 2.992 15.744 ;
    RECT 0.048 15.840 2.992 16.128 ;
    RECT 0.048 16.224 2.992 16.512 ;
    RECT 0.048 16.608 2.992 16.800 ;
    RECT 0 0.000 0.024 0.048 ;
    RECT 0 0.072 0.024 0.336 ;
    RECT 0 0.360 0.024 0.624 ;
    RECT 0 0.648 0.024 0.912 ;
    RECT 0 0.936 0.024 1.200 ;
    RECT 0 1.224 0.024 1.488 ;
    RECT 0 1.512 0.024 1.776 ;
    RECT 0 1.800 0.024 2.064 ;
    RECT 0 2.088 0.024 2.352 ;
    RECT 0 2.376 0.024 2.640 ;
    RECT 0 2.664 0.024 2.928 ;
    RECT 0 2.952 0.024 3.216 ;
    RECT 0 3.240 0.024 3.504 ;
    RECT 0 3.528 0.024 3.792 ;
    RECT 0 3.816 0.024 4.080 ;
    RECT 0 4.104 0.024 4.368 ;
    RECT 0 4.392 0.024 4.656 ;
    RECT 0 4.680 0.024 4.944 ;
    RECT 0 4.968 0.024 5.232 ;
    RECT 0 5.256 0.024 5.520 ;
    RECT 0 5.544 0.024 5.808 ;
    RECT 0 5.832 0.024 6.096 ;
    RECT 0 6.120 0.024 6.432 ;
    RECT 0 6.456 0.024 6.720 ;
    RECT 0 6.744 0.024 7.008 ;
    RECT 0 7.032 0.024 7.296 ;
    RECT 0 7.320 0.024 7.584 ;
    RECT 0 7.608 0.024 7.872 ;
    RECT 0 7.896 0.024 8.160 ;
    RECT 0 8.184 0.024 8.448 ;
    RECT 0 8.472 0.024 8.736 ;
    RECT 0 8.760 0.024 9.024 ;
    RECT 0 9.048 0.024 9.312 ;
    RECT 0 9.336 0.024 9.600 ;
    RECT 0 9.624 0.024 9.888 ;
    RECT 0 9.912 0.024 10.176 ;
    RECT 0 10.200 0.024 10.464 ;
    RECT 0 10.488 0.024 10.752 ;
    RECT 0 10.776 0.024 11.040 ;
    RECT 0 11.064 0.024 11.328 ;
    RECT 0 11.352 0.024 11.616 ;
    RECT 0 11.640 0.024 11.904 ;
    RECT 0 11.928 0.024 12.192 ;
    RECT 0 12.216 0.024 12.480 ;
    RECT 0 12.504 0.024 12.816 ;
    RECT 0 12.840 0.024 13.104 ;
    RECT 0 13.128 0.024 13.392 ;
    RECT 0 13.416 0.024 13.680 ;
    RECT 0 13.704 0.024 13.968 ;
    RECT 0 13.992 0.024 14.256 ;
    RECT 0 14.280 0.024 14.544 ;
    RECT 0 14.568 0.024 14.832 ;
    RECT 0 14.856 0.024 15.120 ;
    RECT 0 15.144 0.024 15.408 ;
    RECT 0 15.432 0.024 15.696 ;
    RECT 0 15.720 0.024 15.984 ;
    RECT 0 16.008 0.024 16.272 ;
    RECT 0 16.296 0.024 16.560 ;
    RECT 0 16.584 0.024 16.848 ;
    RECT 0 16.872 0.024 17.136 ;
    RECT 0 17.160 0.024 17.424 ;
    RECT 0 17.448 0.024 17.712 ;
    RECT 0 17.736 0.024 18.000 ;
    RECT 0 18.024 0.024 18.288 ;
    RECT 0 18.312 0.024 18.576 ;
    RECT 0 18.600 0.024 18.864 ;
    RECT 0 18.888 0.024 19.200 ;
    RECT 0 19.224 0.024 19.488 ;
    RECT 0 19.512 0.024 19.776 ;
    RECT 0 19.800 0.024 20.064 ;
    RECT 0 20.088 0.024 20.352 ;
    RECT 0 20.376 0.024 20.640 ;
    RECT 0 20.664 0.024 20.976 ;
    RECT 0 21.000 0.024 21.264 ;
    RECT 0 21.288 0.024 21.552 ;
    RECT 0 21.576 0.024 16.800 ;
#    LAYER OVERLAP ;
#    RECT 0 0 3.040 16.800 ;
  END
END fakeram_64x22

END LIBRARY
