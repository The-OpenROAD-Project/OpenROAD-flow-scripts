../../../platforms/nangate45/lef/fakeram45_2048x39.lef