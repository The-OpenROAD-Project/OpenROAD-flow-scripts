VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_256x32
  FOREIGN fakeram45_256x32 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 78.660 BY 64.400 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.400 0.070 1.470 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.960 0.070 2.030 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.520 0.070 2.590 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.080 0.070 3.150 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.640 0.070 3.710 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.200 0.070 4.270 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.760 0.070 4.830 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.320 0.070 5.390 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.880 0.070 5.950 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.440 0.070 6.510 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.000 0.070 7.070 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.560 0.070 7.630 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.120 0.070 8.190 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.680 0.070 8.750 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.240 0.070 9.310 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.800 0.070 9.870 ;
    END
  END w_mask_in[15]
  PIN w_mask_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.360 0.070 10.430 ;
    END
  END w_mask_in[16]
  PIN w_mask_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.920 0.070 10.990 ;
    END
  END w_mask_in[17]
  PIN w_mask_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.480 0.070 11.550 ;
    END
  END w_mask_in[18]
  PIN w_mask_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.040 0.070 12.110 ;
    END
  END w_mask_in[19]
  PIN w_mask_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.600 0.070 12.670 ;
    END
  END w_mask_in[20]
  PIN w_mask_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.160 0.070 13.230 ;
    END
  END w_mask_in[21]
  PIN w_mask_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.720 0.070 13.790 ;
    END
  END w_mask_in[22]
  PIN w_mask_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.280 0.070 14.350 ;
    END
  END w_mask_in[23]
  PIN w_mask_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.840 0.070 14.910 ;
    END
  END w_mask_in[24]
  PIN w_mask_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.400 0.070 15.470 ;
    END
  END w_mask_in[25]
  PIN w_mask_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.960 0.070 16.030 ;
    END
  END w_mask_in[26]
  PIN w_mask_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.520 0.070 16.590 ;
    END
  END w_mask_in[27]
  PIN w_mask_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.080 0.070 17.150 ;
    END
  END w_mask_in[28]
  PIN w_mask_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.640 0.070 17.710 ;
    END
  END w_mask_in[29]
  PIN w_mask_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.200 0.070 18.270 ;
    END
  END w_mask_in[30]
  PIN w_mask_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.760 0.070 18.830 ;
    END
  END w_mask_in[31]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.180 0.070 19.250 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.740 0.070 19.810 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.300 0.070 20.370 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.860 0.070 20.930 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.420 0.070 21.490 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.980 0.070 22.050 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.540 0.070 22.610 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.100 0.070 23.170 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.660 0.070 23.730 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.220 0.070 24.290 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.780 0.070 24.850 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.340 0.070 25.410 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.900 0.070 25.970 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.460 0.070 26.530 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.020 0.070 27.090 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.580 0.070 27.650 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.140 0.070 28.210 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.700 0.070 28.770 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.260 0.070 29.330 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.820 0.070 29.890 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.380 0.070 30.450 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.940 0.070 31.010 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.500 0.070 31.570 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.060 0.070 32.130 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.620 0.070 32.690 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.180 0.070 33.250 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.740 0.070 33.810 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.300 0.070 34.370 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 34.860 0.070 34.930 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.420 0.070 35.490 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.980 0.070 36.050 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.540 0.070 36.610 ;
    END
  END rd_out[31]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.960 0.070 37.030 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 37.520 0.070 37.590 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.080 0.070 38.150 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 38.640 0.070 38.710 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.200 0.070 39.270 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 39.760 0.070 39.830 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.320 0.070 40.390 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 40.880 0.070 40.950 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 41.440 0.070 41.510 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.000 0.070 42.070 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 42.560 0.070 42.630 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.120 0.070 43.190 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 43.680 0.070 43.750 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.240 0.070 44.310 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 44.800 0.070 44.870 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.360 0.070 45.430 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 45.920 0.070 45.990 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 46.480 0.070 46.550 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.040 0.070 47.110 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 47.600 0.070 47.670 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.160 0.070 48.230 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 48.720 0.070 48.790 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.280 0.070 49.350 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 49.840 0.070 49.910 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.400 0.070 50.470 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 50.960 0.070 51.030 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 51.520 0.070 51.590 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.080 0.070 52.150 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 52.640 0.070 52.710 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.200 0.070 53.270 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 53.760 0.070 53.830 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.320 0.070 54.390 ;
    END
  END wd_in[31]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 54.740 0.070 54.810 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.300 0.070 55.370 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 55.860 0.070 55.930 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.420 0.070 56.490 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 56.980 0.070 57.050 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 57.540 0.070 57.610 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.100 0.070 58.170 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 58.660 0.070 58.730 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.080 0.070 59.150 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 59.640 0.070 59.710 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 60.200 0.070 60.270 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 63.000 ;
      RECT 3.500 1.400 3.780 63.000 ;
      RECT 5.740 1.400 6.020 63.000 ;
      RECT 7.980 1.400 8.260 63.000 ;
      RECT 10.220 1.400 10.500 63.000 ;
      RECT 12.460 1.400 12.740 63.000 ;
      RECT 14.700 1.400 14.980 63.000 ;
      RECT 16.940 1.400 17.220 63.000 ;
      RECT 19.180 1.400 19.460 63.000 ;
      RECT 21.420 1.400 21.700 63.000 ;
      RECT 23.660 1.400 23.940 63.000 ;
      RECT 25.900 1.400 26.180 63.000 ;
      RECT 28.140 1.400 28.420 63.000 ;
      RECT 30.380 1.400 30.660 63.000 ;
      RECT 32.620 1.400 32.900 63.000 ;
      RECT 34.860 1.400 35.140 63.000 ;
      RECT 37.100 1.400 37.380 63.000 ;
      RECT 39.340 1.400 39.620 63.000 ;
      RECT 41.580 1.400 41.860 63.000 ;
      RECT 43.820 1.400 44.100 63.000 ;
      RECT 46.060 1.400 46.340 63.000 ;
      RECT 48.300 1.400 48.580 63.000 ;
      RECT 50.540 1.400 50.820 63.000 ;
      RECT 52.780 1.400 53.060 63.000 ;
      RECT 55.020 1.400 55.300 63.000 ;
      RECT 57.260 1.400 57.540 63.000 ;
      RECT 59.500 1.400 59.780 63.000 ;
      RECT 61.740 1.400 62.020 63.000 ;
      RECT 63.980 1.400 64.260 63.000 ;
      RECT 66.220 1.400 66.500 63.000 ;
      RECT 68.460 1.400 68.740 63.000 ;
      RECT 70.700 1.400 70.980 63.000 ;
      RECT 72.940 1.400 73.220 63.000 ;
      RECT 75.180 1.400 75.460 63.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 63.000 ;
      RECT 4.620 1.400 4.900 63.000 ;
      RECT 6.860 1.400 7.140 63.000 ;
      RECT 9.100 1.400 9.380 63.000 ;
      RECT 11.340 1.400 11.620 63.000 ;
      RECT 13.580 1.400 13.860 63.000 ;
      RECT 15.820 1.400 16.100 63.000 ;
      RECT 18.060 1.400 18.340 63.000 ;
      RECT 20.300 1.400 20.580 63.000 ;
      RECT 22.540 1.400 22.820 63.000 ;
      RECT 24.780 1.400 25.060 63.000 ;
      RECT 27.020 1.400 27.300 63.000 ;
      RECT 29.260 1.400 29.540 63.000 ;
      RECT 31.500 1.400 31.780 63.000 ;
      RECT 33.740 1.400 34.020 63.000 ;
      RECT 35.980 1.400 36.260 63.000 ;
      RECT 38.220 1.400 38.500 63.000 ;
      RECT 40.460 1.400 40.740 63.000 ;
      RECT 42.700 1.400 42.980 63.000 ;
      RECT 44.940 1.400 45.220 63.000 ;
      RECT 47.180 1.400 47.460 63.000 ;
      RECT 49.420 1.400 49.700 63.000 ;
      RECT 51.660 1.400 51.940 63.000 ;
      RECT 53.900 1.400 54.180 63.000 ;
      RECT 56.140 1.400 56.420 63.000 ;
      RECT 58.380 1.400 58.660 63.000 ;
      RECT 60.620 1.400 60.900 63.000 ;
      RECT 62.860 1.400 63.140 63.000 ;
      RECT 65.100 1.400 65.380 63.000 ;
      RECT 67.340 1.400 67.620 63.000 ;
      RECT 69.580 1.400 69.860 63.000 ;
      RECT 71.820 1.400 72.100 63.000 ;
      RECT 74.060 1.400 74.340 63.000 ;
      RECT 76.300 1.400 76.580 63.000 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 78.660 64.400 ;
    LAYER metal2 ;
    RECT 0 0 78.660 64.400 ;
    LAYER metal3 ;
    RECT 0.070 0 78.660 64.400 ;
    RECT 0 0.000 0.070 1.400 ;
    RECT 0 1.470 0.070 1.960 ;
    RECT 0 2.030 0.070 2.520 ;
    RECT 0 2.590 0.070 3.080 ;
    RECT 0 3.150 0.070 3.640 ;
    RECT 0 3.710 0.070 4.200 ;
    RECT 0 4.270 0.070 4.760 ;
    RECT 0 4.830 0.070 5.320 ;
    RECT 0 5.390 0.070 5.880 ;
    RECT 0 5.950 0.070 6.440 ;
    RECT 0 6.510 0.070 7.000 ;
    RECT 0 7.070 0.070 7.560 ;
    RECT 0 7.630 0.070 8.120 ;
    RECT 0 8.190 0.070 8.680 ;
    RECT 0 8.750 0.070 9.240 ;
    RECT 0 9.310 0.070 9.800 ;
    RECT 0 9.870 0.070 10.360 ;
    RECT 0 10.430 0.070 10.920 ;
    RECT 0 10.990 0.070 11.480 ;
    RECT 0 11.550 0.070 12.040 ;
    RECT 0 12.110 0.070 12.600 ;
    RECT 0 12.670 0.070 13.160 ;
    RECT 0 13.230 0.070 13.720 ;
    RECT 0 13.790 0.070 14.280 ;
    RECT 0 14.350 0.070 14.840 ;
    RECT 0 14.910 0.070 15.400 ;
    RECT 0 15.470 0.070 15.960 ;
    RECT 0 16.030 0.070 16.520 ;
    RECT 0 16.590 0.070 17.080 ;
    RECT 0 17.150 0.070 17.640 ;
    RECT 0 17.710 0.070 18.200 ;
    RECT 0 18.270 0.070 18.760 ;
    RECT 0 18.830 0.070 19.180 ;
    RECT 0 19.250 0.070 19.740 ;
    RECT 0 19.810 0.070 20.300 ;
    RECT 0 20.370 0.070 20.860 ;
    RECT 0 20.930 0.070 21.420 ;
    RECT 0 21.490 0.070 21.980 ;
    RECT 0 22.050 0.070 22.540 ;
    RECT 0 22.610 0.070 23.100 ;
    RECT 0 23.170 0.070 23.660 ;
    RECT 0 23.730 0.070 24.220 ;
    RECT 0 24.290 0.070 24.780 ;
    RECT 0 24.850 0.070 25.340 ;
    RECT 0 25.410 0.070 25.900 ;
    RECT 0 25.970 0.070 26.460 ;
    RECT 0 26.530 0.070 27.020 ;
    RECT 0 27.090 0.070 27.580 ;
    RECT 0 27.650 0.070 28.140 ;
    RECT 0 28.210 0.070 28.700 ;
    RECT 0 28.770 0.070 29.260 ;
    RECT 0 29.330 0.070 29.820 ;
    RECT 0 29.890 0.070 30.380 ;
    RECT 0 30.450 0.070 30.940 ;
    RECT 0 31.010 0.070 31.500 ;
    RECT 0 31.570 0.070 32.060 ;
    RECT 0 32.130 0.070 32.620 ;
    RECT 0 32.690 0.070 33.180 ;
    RECT 0 33.250 0.070 33.740 ;
    RECT 0 33.810 0.070 34.300 ;
    RECT 0 34.370 0.070 34.860 ;
    RECT 0 34.930 0.070 35.420 ;
    RECT 0 35.490 0.070 35.980 ;
    RECT 0 36.050 0.070 36.540 ;
    RECT 0 36.610 0.070 36.960 ;
    RECT 0 37.030 0.070 37.520 ;
    RECT 0 37.590 0.070 38.080 ;
    RECT 0 38.150 0.070 38.640 ;
    RECT 0 38.710 0.070 39.200 ;
    RECT 0 39.270 0.070 39.760 ;
    RECT 0 39.830 0.070 40.320 ;
    RECT 0 40.390 0.070 40.880 ;
    RECT 0 40.950 0.070 41.440 ;
    RECT 0 41.510 0.070 42.000 ;
    RECT 0 42.070 0.070 42.560 ;
    RECT 0 42.630 0.070 43.120 ;
    RECT 0 43.190 0.070 43.680 ;
    RECT 0 43.750 0.070 44.240 ;
    RECT 0 44.310 0.070 44.800 ;
    RECT 0 44.870 0.070 45.360 ;
    RECT 0 45.430 0.070 45.920 ;
    RECT 0 45.990 0.070 46.480 ;
    RECT 0 46.550 0.070 47.040 ;
    RECT 0 47.110 0.070 47.600 ;
    RECT 0 47.670 0.070 48.160 ;
    RECT 0 48.230 0.070 48.720 ;
    RECT 0 48.790 0.070 49.280 ;
    RECT 0 49.350 0.070 49.840 ;
    RECT 0 49.910 0.070 50.400 ;
    RECT 0 50.470 0.070 50.960 ;
    RECT 0 51.030 0.070 51.520 ;
    RECT 0 51.590 0.070 52.080 ;
    RECT 0 52.150 0.070 52.640 ;
    RECT 0 52.710 0.070 53.200 ;
    RECT 0 53.270 0.070 53.760 ;
    RECT 0 53.830 0.070 54.320 ;
    RECT 0 54.390 0.070 54.740 ;
    RECT 0 54.810 0.070 55.300 ;
    RECT 0 55.370 0.070 55.860 ;
    RECT 0 55.930 0.070 56.420 ;
    RECT 0 56.490 0.070 56.980 ;
    RECT 0 57.050 0.070 57.540 ;
    RECT 0 57.610 0.070 58.100 ;
    RECT 0 58.170 0.070 58.660 ;
    RECT 0 58.730 0.070 59.080 ;
    RECT 0 59.150 0.070 59.640 ;
    RECT 0 59.710 0.070 60.200 ;
    RECT 0 60.270 0.070 64.400 ;
    LAYER metal4 ;
    RECT 0 0 78.660 1.400 ;
    RECT 0 63.000 78.660 64.400 ;
    RECT 0.000 1.400 1.260 63.000 ;
    RECT 1.540 1.400 2.380 63.000 ;
    RECT 2.660 1.400 3.500 63.000 ;
    RECT 3.780 1.400 4.620 63.000 ;
    RECT 4.900 1.400 5.740 63.000 ;
    RECT 6.020 1.400 6.860 63.000 ;
    RECT 7.140 1.400 7.980 63.000 ;
    RECT 8.260 1.400 9.100 63.000 ;
    RECT 9.380 1.400 10.220 63.000 ;
    RECT 10.500 1.400 11.340 63.000 ;
    RECT 11.620 1.400 12.460 63.000 ;
    RECT 12.740 1.400 13.580 63.000 ;
    RECT 13.860 1.400 14.700 63.000 ;
    RECT 14.980 1.400 15.820 63.000 ;
    RECT 16.100 1.400 16.940 63.000 ;
    RECT 17.220 1.400 18.060 63.000 ;
    RECT 18.340 1.400 19.180 63.000 ;
    RECT 19.460 1.400 20.300 63.000 ;
    RECT 20.580 1.400 21.420 63.000 ;
    RECT 21.700 1.400 22.540 63.000 ;
    RECT 22.820 1.400 23.660 63.000 ;
    RECT 23.940 1.400 24.780 63.000 ;
    RECT 25.060 1.400 25.900 63.000 ;
    RECT 26.180 1.400 27.020 63.000 ;
    RECT 27.300 1.400 28.140 63.000 ;
    RECT 28.420 1.400 29.260 63.000 ;
    RECT 29.540 1.400 30.380 63.000 ;
    RECT 30.660 1.400 31.500 63.000 ;
    RECT 31.780 1.400 32.620 63.000 ;
    RECT 32.900 1.400 33.740 63.000 ;
    RECT 34.020 1.400 34.860 63.000 ;
    RECT 35.140 1.400 35.980 63.000 ;
    RECT 36.260 1.400 37.100 63.000 ;
    RECT 37.380 1.400 38.220 63.000 ;
    RECT 38.500 1.400 39.340 63.000 ;
    RECT 39.620 1.400 40.460 63.000 ;
    RECT 40.740 1.400 41.580 63.000 ;
    RECT 41.860 1.400 42.700 63.000 ;
    RECT 42.980 1.400 43.820 63.000 ;
    RECT 44.100 1.400 44.940 63.000 ;
    RECT 45.220 1.400 46.060 63.000 ;
    RECT 46.340 1.400 47.180 63.000 ;
    RECT 47.460 1.400 48.300 63.000 ;
    RECT 48.580 1.400 49.420 63.000 ;
    RECT 49.700 1.400 50.540 63.000 ;
    RECT 50.820 1.400 51.660 63.000 ;
    RECT 51.940 1.400 52.780 63.000 ;
    RECT 53.060 1.400 53.900 63.000 ;
    RECT 54.180 1.400 55.020 63.000 ;
    RECT 55.300 1.400 56.140 63.000 ;
    RECT 56.420 1.400 57.260 63.000 ;
    RECT 57.540 1.400 58.380 63.000 ;
    RECT 58.660 1.400 59.500 63.000 ;
    RECT 59.780 1.400 60.620 63.000 ;
    RECT 60.900 1.400 61.740 63.000 ;
    RECT 62.020 1.400 62.860 63.000 ;
    RECT 63.140 1.400 63.980 63.000 ;
    RECT 64.260 1.400 65.100 63.000 ;
    RECT 65.380 1.400 66.220 63.000 ;
    RECT 66.500 1.400 67.340 63.000 ;
    RECT 67.620 1.400 68.460 63.000 ;
    RECT 68.740 1.400 69.580 63.000 ;
    RECT 69.860 1.400 70.700 63.000 ;
    RECT 70.980 1.400 71.820 63.000 ;
    RECT 72.100 1.400 72.940 63.000 ;
    RECT 73.220 1.400 74.060 63.000 ;
    RECT 74.340 1.400 75.180 63.000 ;
    RECT 75.460 1.400 76.300 63.000 ;
    RECT 76.580 1.400 78.660 63.000 ;
    LAYER OVERLAP ;
    RECT 0 0 78.660 64.400 ;
  END
END fakeram45_256x32

END LIBRARY
