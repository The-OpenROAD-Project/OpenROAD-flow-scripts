../../../platforms/nangate45/lef/fakeram45_64x21.lef