VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram130_256x16
  FOREIGN fakeram130_256x16 0 0 ;
  SYMMETRY X Y ;
  SIZE 285.660 BY 187.680 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 4.370 0.460 4.830 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 7.130 0.460 7.590 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 9.890 0.460 10.350 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 12.650 0.460 13.110 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 15.410 0.460 15.870 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 18.170 0.460 18.630 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 20.930 0.460 21.390 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 23.690 0.460 24.150 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 26.450 0.460 26.910 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 29.210 0.460 29.670 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 31.970 0.460 32.430 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 34.730 0.460 35.190 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 37.490 0.460 37.950 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 40.250 0.460 40.710 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 43.010 0.460 43.470 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 45.770 0.460 46.230 ;
    END
  END w_mask_in[15]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 49.450 0.460 49.910 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 52.210 0.460 52.670 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 54.970 0.460 55.430 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 57.730 0.460 58.190 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 60.490 0.460 60.950 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 63.250 0.460 63.710 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 66.010 0.460 66.470 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 68.770 0.460 69.230 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 71.530 0.460 71.990 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 74.290 0.460 74.750 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 77.050 0.460 77.510 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 79.810 0.460 80.270 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 82.570 0.460 83.030 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 85.330 0.460 85.790 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 88.090 0.460 88.550 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 90.850 0.460 91.310 ;
    END
  END rd_out[15]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 94.530 0.460 94.990 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 97.290 0.460 97.750 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 100.050 0.460 100.510 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 102.810 0.460 103.270 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 105.570 0.460 106.030 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 108.330 0.460 108.790 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 111.090 0.460 111.550 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 113.850 0.460 114.310 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 116.610 0.460 117.070 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 119.370 0.460 119.830 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 122.130 0.460 122.590 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 124.890 0.460 125.350 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 127.650 0.460 128.110 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 130.410 0.460 130.870 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 133.170 0.460 133.630 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 135.930 0.460 136.390 ;
    END
  END wd_in[15]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 139.610 0.460 140.070 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 142.370 0.460 142.830 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 145.130 0.460 145.590 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 147.890 0.460 148.350 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 150.650 0.460 151.110 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 153.410 0.460 153.870 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 156.170 0.460 156.630 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 158.930 0.460 159.390 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 162.610 0.460 163.070 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 165.370 0.460 165.830 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
      RECT 0.000 168.130 0.460 168.590 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
      RECT 3.680 4.600 5.520 183.080 ;
      RECT 11.040 4.600 12.880 183.080 ;
      RECT 18.400 4.600 20.240 183.080 ;
      RECT 25.760 4.600 27.600 183.080 ;
      RECT 33.120 4.600 34.960 183.080 ;
      RECT 40.480 4.600 42.320 183.080 ;
      RECT 47.840 4.600 49.680 183.080 ;
      RECT 55.200 4.600 57.040 183.080 ;
      RECT 62.560 4.600 64.400 183.080 ;
      RECT 69.920 4.600 71.760 183.080 ;
      RECT 77.280 4.600 79.120 183.080 ;
      RECT 84.640 4.600 86.480 183.080 ;
      RECT 92.000 4.600 93.840 183.080 ;
      RECT 99.360 4.600 101.200 183.080 ;
      RECT 106.720 4.600 108.560 183.080 ;
      RECT 114.080 4.600 115.920 183.080 ;
      RECT 121.440 4.600 123.280 183.080 ;
      RECT 128.800 4.600 130.640 183.080 ;
      RECT 136.160 4.600 138.000 183.080 ;
      RECT 143.520 4.600 145.360 183.080 ;
      RECT 150.880 4.600 152.720 183.080 ;
      RECT 158.240 4.600 160.080 183.080 ;
      RECT 165.600 4.600 167.440 183.080 ;
      RECT 172.960 4.600 174.800 183.080 ;
      RECT 180.320 4.600 182.160 183.080 ;
      RECT 187.680 4.600 189.520 183.080 ;
      RECT 195.040 4.600 196.880 183.080 ;
      RECT 202.400 4.600 204.240 183.080 ;
      RECT 209.760 4.600 211.600 183.080 ;
      RECT 217.120 4.600 218.960 183.080 ;
      RECT 224.480 4.600 226.320 183.080 ;
      RECT 231.840 4.600 233.680 183.080 ;
      RECT 239.200 4.600 241.040 183.080 ;
      RECT 246.560 4.600 248.400 183.080 ;
      RECT 253.920 4.600 255.760 183.080 ;
      RECT 261.280 4.600 263.120 183.080 ;
      RECT 268.640 4.600 270.480 183.080 ;
      RECT 276.000 4.600 277.840 183.080 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
      RECT 7.360 4.600 9.200 183.080 ;
      RECT 14.720 4.600 16.560 183.080 ;
      RECT 22.080 4.600 23.920 183.080 ;
      RECT 29.440 4.600 31.280 183.080 ;
      RECT 36.800 4.600 38.640 183.080 ;
      RECT 44.160 4.600 46.000 183.080 ;
      RECT 51.520 4.600 53.360 183.080 ;
      RECT 58.880 4.600 60.720 183.080 ;
      RECT 66.240 4.600 68.080 183.080 ;
      RECT 73.600 4.600 75.440 183.080 ;
      RECT 80.960 4.600 82.800 183.080 ;
      RECT 88.320 4.600 90.160 183.080 ;
      RECT 95.680 4.600 97.520 183.080 ;
      RECT 103.040 4.600 104.880 183.080 ;
      RECT 110.400 4.600 112.240 183.080 ;
      RECT 117.760 4.600 119.600 183.080 ;
      RECT 125.120 4.600 126.960 183.080 ;
      RECT 132.480 4.600 134.320 183.080 ;
      RECT 139.840 4.600 141.680 183.080 ;
      RECT 147.200 4.600 149.040 183.080 ;
      RECT 154.560 4.600 156.400 183.080 ;
      RECT 161.920 4.600 163.760 183.080 ;
      RECT 169.280 4.600 171.120 183.080 ;
      RECT 176.640 4.600 178.480 183.080 ;
      RECT 184.000 4.600 185.840 183.080 ;
      RECT 191.360 4.600 193.200 183.080 ;
      RECT 198.720 4.600 200.560 183.080 ;
      RECT 206.080 4.600 207.920 183.080 ;
      RECT 213.440 4.600 215.280 183.080 ;
      RECT 220.800 4.600 222.640 183.080 ;
      RECT 228.160 4.600 230.000 183.080 ;
      RECT 235.520 4.600 237.360 183.080 ;
      RECT 242.880 4.600 244.720 183.080 ;
      RECT 250.240 4.600 252.080 183.080 ;
      RECT 257.600 4.600 259.440 183.080 ;
      RECT 264.960 4.600 266.800 183.080 ;
      RECT 272.320 4.600 274.160 183.080 ;
      RECT 279.680 4.600 281.520 183.080 ;
    END
  END VDD
  OBS
    LAYER met1 ;
    RECT 0 0 285.660 187.680 ;
    LAYER met2 ;
    RECT 0 0 285.660 187.680 ;
    LAYER met3 ;
    RECT 0.460 0 285.660 187.680 ;
    RECT 0 0.000 0.460 4.370 ;
    RECT 0 4.830 0.460 7.130 ;
    RECT 0 7.590 0.460 9.890 ;
    RECT 0 10.350 0.460 12.650 ;
    RECT 0 13.110 0.460 15.410 ;
    RECT 0 15.870 0.460 18.170 ;
    RECT 0 18.630 0.460 20.930 ;
    RECT 0 21.390 0.460 23.690 ;
    RECT 0 24.150 0.460 26.450 ;
    RECT 0 26.910 0.460 29.210 ;
    RECT 0 29.670 0.460 31.970 ;
    RECT 0 32.430 0.460 34.730 ;
    RECT 0 35.190 0.460 37.490 ;
    RECT 0 37.950 0.460 40.250 ;
    RECT 0 40.710 0.460 43.010 ;
    RECT 0 43.470 0.460 45.770 ;
    RECT 0 46.230 0.460 49.450 ;
    RECT 0 49.910 0.460 52.210 ;
    RECT 0 52.670 0.460 54.970 ;
    RECT 0 55.430 0.460 57.730 ;
    RECT 0 58.190 0.460 60.490 ;
    RECT 0 60.950 0.460 63.250 ;
    RECT 0 63.710 0.460 66.010 ;
    RECT 0 66.470 0.460 68.770 ;
    RECT 0 69.230 0.460 71.530 ;
    RECT 0 71.990 0.460 74.290 ;
    RECT 0 74.750 0.460 77.050 ;
    RECT 0 77.510 0.460 79.810 ;
    RECT 0 80.270 0.460 82.570 ;
    RECT 0 83.030 0.460 85.330 ;
    RECT 0 85.790 0.460 88.090 ;
    RECT 0 88.550 0.460 90.850 ;
    RECT 0 91.310 0.460 94.530 ;
    RECT 0 94.990 0.460 97.290 ;
    RECT 0 97.750 0.460 100.050 ;
    RECT 0 100.510 0.460 102.810 ;
    RECT 0 103.270 0.460 105.570 ;
    RECT 0 106.030 0.460 108.330 ;
    RECT 0 108.790 0.460 111.090 ;
    RECT 0 111.550 0.460 113.850 ;
    RECT 0 114.310 0.460 116.610 ;
    RECT 0 117.070 0.460 119.370 ;
    RECT 0 119.830 0.460 122.130 ;
    RECT 0 122.590 0.460 124.890 ;
    RECT 0 125.350 0.460 127.650 ;
    RECT 0 128.110 0.460 130.410 ;
    RECT 0 130.870 0.460 133.170 ;
    RECT 0 133.630 0.460 135.930 ;
    RECT 0 136.390 0.460 139.610 ;
    RECT 0 140.070 0.460 142.370 ;
    RECT 0 142.830 0.460 145.130 ;
    RECT 0 145.590 0.460 147.890 ;
    RECT 0 148.350 0.460 150.650 ;
    RECT 0 151.110 0.460 153.410 ;
    RECT 0 153.870 0.460 156.170 ;
    RECT 0 156.630 0.460 158.930 ;
    RECT 0 159.390 0.460 162.610 ;
    RECT 0 163.070 0.460 165.370 ;
    RECT 0 165.830 0.460 168.130 ;
    RECT 0 168.590 0.460 187.680 ;
    LAYER met4 ;
    RECT 0 0 285.660 4.600 ;
    RECT 0 183.080 285.660 187.680 ;
    RECT 0.000 4.600 3.680 183.080 ;
    RECT 5.520 4.600 7.360 183.080 ;
    RECT 9.200 4.600 11.040 183.080 ;
    RECT 12.880 4.600 14.720 183.080 ;
    RECT 16.560 4.600 18.400 183.080 ;
    RECT 20.240 4.600 22.080 183.080 ;
    RECT 23.920 4.600 25.760 183.080 ;
    RECT 27.600 4.600 29.440 183.080 ;
    RECT 31.280 4.600 33.120 183.080 ;
    RECT 34.960 4.600 36.800 183.080 ;
    RECT 38.640 4.600 40.480 183.080 ;
    RECT 42.320 4.600 44.160 183.080 ;
    RECT 46.000 4.600 47.840 183.080 ;
    RECT 49.680 4.600 51.520 183.080 ;
    RECT 53.360 4.600 55.200 183.080 ;
    RECT 57.040 4.600 58.880 183.080 ;
    RECT 60.720 4.600 62.560 183.080 ;
    RECT 64.400 4.600 66.240 183.080 ;
    RECT 68.080 4.600 69.920 183.080 ;
    RECT 71.760 4.600 73.600 183.080 ;
    RECT 75.440 4.600 77.280 183.080 ;
    RECT 79.120 4.600 80.960 183.080 ;
    RECT 82.800 4.600 84.640 183.080 ;
    RECT 86.480 4.600 88.320 183.080 ;
    RECT 90.160 4.600 92.000 183.080 ;
    RECT 93.840 4.600 95.680 183.080 ;
    RECT 97.520 4.600 99.360 183.080 ;
    RECT 101.200 4.600 103.040 183.080 ;
    RECT 104.880 4.600 106.720 183.080 ;
    RECT 108.560 4.600 110.400 183.080 ;
    RECT 112.240 4.600 114.080 183.080 ;
    RECT 115.920 4.600 117.760 183.080 ;
    RECT 119.600 4.600 121.440 183.080 ;
    RECT 123.280 4.600 125.120 183.080 ;
    RECT 126.960 4.600 128.800 183.080 ;
    RECT 130.640 4.600 132.480 183.080 ;
    RECT 134.320 4.600 136.160 183.080 ;
    RECT 138.000 4.600 139.840 183.080 ;
    RECT 141.680 4.600 143.520 183.080 ;
    RECT 145.360 4.600 147.200 183.080 ;
    RECT 149.040 4.600 150.880 183.080 ;
    RECT 152.720 4.600 154.560 183.080 ;
    RECT 156.400 4.600 158.240 183.080 ;
    RECT 160.080 4.600 161.920 183.080 ;
    RECT 163.760 4.600 165.600 183.080 ;
    RECT 167.440 4.600 169.280 183.080 ;
    RECT 171.120 4.600 172.960 183.080 ;
    RECT 174.800 4.600 176.640 183.080 ;
    RECT 178.480 4.600 180.320 183.080 ;
    RECT 182.160 4.600 184.000 183.080 ;
    RECT 185.840 4.600 187.680 183.080 ;
    RECT 189.520 4.600 191.360 183.080 ;
    RECT 193.200 4.600 195.040 183.080 ;
    RECT 196.880 4.600 198.720 183.080 ;
    RECT 200.560 4.600 202.400 183.080 ;
    RECT 204.240 4.600 206.080 183.080 ;
    RECT 207.920 4.600 209.760 183.080 ;
    RECT 211.600 4.600 213.440 183.080 ;
    RECT 215.280 4.600 217.120 183.080 ;
    RECT 218.960 4.600 220.800 183.080 ;
    RECT 222.640 4.600 224.480 183.080 ;
    RECT 226.320 4.600 228.160 183.080 ;
    RECT 230.000 4.600 231.840 183.080 ;
    RECT 233.680 4.600 235.520 183.080 ;
    RECT 237.360 4.600 239.200 183.080 ;
    RECT 241.040 4.600 242.880 183.080 ;
    RECT 244.720 4.600 246.560 183.080 ;
    RECT 248.400 4.600 250.240 183.080 ;
    RECT 252.080 4.600 253.920 183.080 ;
    RECT 255.760 4.600 257.600 183.080 ;
    RECT 259.440 4.600 261.280 183.080 ;
    RECT 263.120 4.600 264.960 183.080 ;
    RECT 266.800 4.600 268.640 183.080 ;
    RECT 270.480 4.600 272.320 183.080 ;
    RECT 274.160 4.600 276.000 183.080 ;
    RECT 277.840 4.600 279.680 183.080 ;
    RECT 281.520 4.600 285.660 183.080 ;
    LAYER OVERLAP ;
    RECT 0 0 285.660 187.680 ;
  END
END fakeram130_256x16

END LIBRARY
