module Element (clock,
    io_lsbIns_1,
    io_lsbIns_2,
    io_lsbIns_3,
    io_lsbIns_4,
    io_lsbIns_5,
    io_lsbIns_6,
    io_lsbIns_7,
    io_lsbOuts_0,
    io_lsbOuts_1,
    io_lsbOuts_2,
    io_lsbOuts_3,
    io_lsbOuts_4,
    io_lsbOuts_5,
    io_lsbOuts_6,
    io_lsbOuts_7,
    io_ins_down,
    io_ins_left,
    io_ins_right,
    io_ins_up,
    io_outs_down,
    io_outs_left,
    io_outs_right,
    io_outs_up);
 input clock;
 input io_lsbIns_1;
 input io_lsbIns_2;
 input io_lsbIns_3;
 input io_lsbIns_4;
 input io_lsbIns_5;
 input io_lsbIns_6;
 input io_lsbIns_7;
 output io_lsbOuts_0;
 output io_lsbOuts_1;
 output io_lsbOuts_2;
 output io_lsbOuts_3;
 output io_lsbOuts_4;
 output io_lsbOuts_5;
 output io_lsbOuts_6;
 output io_lsbOuts_7;
 input [63:0] io_ins_down;
 input [63:0] io_ins_left;
 input [63:0] io_ins_right;
 input [63:0] io_ins_up;
 output [63:0] io_outs_down;
 output [63:0] io_outs_left;
 output [63:0] io_outs_right;
 output [63:0] io_outs_up;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire clknet_leaf_0_clock;
 wire clknet_leaf_1_clock;
 wire clknet_leaf_2_clock;
 wire clknet_leaf_3_clock;
 wire clknet_leaf_4_clock;
 wire clknet_leaf_5_clock;
 wire clknet_leaf_6_clock;
 wire clknet_leaf_7_clock;
 wire clknet_leaf_8_clock;
 wire clknet_leaf_9_clock;
 wire clknet_leaf_10_clock;
 wire clknet_leaf_11_clock;
 wire clknet_leaf_12_clock;
 wire clknet_leaf_13_clock;
 wire clknet_leaf_14_clock;
 wire clknet_leaf_15_clock;
 wire clknet_leaf_16_clock;
 wire clknet_leaf_17_clock;
 wire clknet_leaf_18_clock;
 wire clknet_leaf_19_clock;
 wire clknet_leaf_20_clock;
 wire clknet_0_clock;
 wire clknet_1_0__leaf_clock;
 wire clknet_1_1__leaf_clock;

 DFFHQNx2_ASAP7_75t_R \REG[0]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(net1),
    .QN(_0257_));
 DFFHQNx2_ASAP7_75t_R \REG[10]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net2),
    .QN(_0267_));
 DFFHQNx2_ASAP7_75t_R \REG[11]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(net3),
    .QN(_0268_));
 DFFHQNx2_ASAP7_75t_R \REG[12]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net4),
    .QN(_0269_));
 DFFHQNx2_ASAP7_75t_R \REG[13]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(net5),
    .QN(_0270_));
 DFFHQNx2_ASAP7_75t_R \REG[14]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(net6),
    .QN(_0271_));
 DFFHQNx2_ASAP7_75t_R \REG[15]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(net7),
    .QN(_0272_));
 DFFHQNx2_ASAP7_75t_R \REG[16]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(net8),
    .QN(_0273_));
 DFFHQNx2_ASAP7_75t_R \REG[17]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net9),
    .QN(_0274_));
 DFFHQNx2_ASAP7_75t_R \REG[18]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(net10),
    .QN(_0275_));
 DFFHQNx2_ASAP7_75t_R \REG[19]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net11),
    .QN(_0276_));
 DFFHQNx2_ASAP7_75t_R \REG[1]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(net12),
    .QN(_0258_));
 DFFHQNx2_ASAP7_75t_R \REG[20]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net13),
    .QN(_0277_));
 DFFHQNx2_ASAP7_75t_R \REG[21]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net14),
    .QN(_0278_));
 DFFHQNx2_ASAP7_75t_R \REG[22]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net15),
    .QN(_0279_));
 DFFHQNx2_ASAP7_75t_R \REG[23]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net16),
    .QN(_0280_));
 DFFHQNx2_ASAP7_75t_R \REG[24]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net17),
    .QN(_0281_));
 DFFHQNx2_ASAP7_75t_R \REG[25]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net18),
    .QN(_0282_));
 DFFHQNx2_ASAP7_75t_R \REG[26]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net19),
    .QN(_0283_));
 DFFHQNx2_ASAP7_75t_R \REG[27]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net20),
    .QN(_0284_));
 DFFHQNx2_ASAP7_75t_R \REG[28]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net21),
    .QN(_0285_));
 DFFHQNx2_ASAP7_75t_R \REG[29]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net22),
    .QN(_0286_));
 DFFHQNx2_ASAP7_75t_R \REG[2]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(net23),
    .QN(_0259_));
 DFFHQNx2_ASAP7_75t_R \REG[30]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net24),
    .QN(_0287_));
 DFFHQNx2_ASAP7_75t_R \REG[31]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(net25),
    .QN(_0288_));
 DFFHQNx2_ASAP7_75t_R \REG[32]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net26),
    .QN(_0289_));
 DFFHQNx2_ASAP7_75t_R \REG[33]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net27),
    .QN(_0290_));
 DFFHQNx2_ASAP7_75t_R \REG[34]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net28),
    .QN(_0291_));
 DFFHQNx2_ASAP7_75t_R \REG[35]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net29),
    .QN(_0292_));
 DFFHQNx2_ASAP7_75t_R \REG[36]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net30),
    .QN(_0293_));
 DFFHQNx2_ASAP7_75t_R \REG[37]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net31),
    .QN(_0294_));
 DFFHQNx2_ASAP7_75t_R \REG[38]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net32),
    .QN(_0295_));
 DFFHQNx2_ASAP7_75t_R \REG[39]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(net33),
    .QN(_0296_));
 DFFHQNx2_ASAP7_75t_R \REG[3]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net34),
    .QN(_0260_));
 DFFHQNx2_ASAP7_75t_R \REG[40]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(net35),
    .QN(_0297_));
 DFFHQNx2_ASAP7_75t_R \REG[41]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net36),
    .QN(_0298_));
 DFFHQNx2_ASAP7_75t_R \REG[42]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net37),
    .QN(_0299_));
 DFFHQNx2_ASAP7_75t_R \REG[43]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net38),
    .QN(_0300_));
 DFFHQNx2_ASAP7_75t_R \REG[44]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net39),
    .QN(_0301_));
 DFFHQNx2_ASAP7_75t_R \REG[45]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net40),
    .QN(_0302_));
 DFFHQNx2_ASAP7_75t_R \REG[46]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net41),
    .QN(_0303_));
 DFFHQNx2_ASAP7_75t_R \REG[47]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net42),
    .QN(_0304_));
 DFFHQNx2_ASAP7_75t_R \REG[48]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net43),
    .QN(_0305_));
 DFFHQNx2_ASAP7_75t_R \REG[49]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net44),
    .QN(_0306_));
 DFFHQNx2_ASAP7_75t_R \REG[4]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(net45),
    .QN(_0261_));
 DFFHQNx2_ASAP7_75t_R \REG[50]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net46),
    .QN(_0307_));
 DFFHQNx2_ASAP7_75t_R \REG[51]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net47),
    .QN(_0308_));
 DFFHQNx2_ASAP7_75t_R \REG[52]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net48),
    .QN(_0309_));
 DFFHQNx2_ASAP7_75t_R \REG[53]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net49),
    .QN(_0310_));
 DFFHQNx2_ASAP7_75t_R \REG[54]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(net50),
    .QN(_0311_));
 DFFHQNx2_ASAP7_75t_R \REG[55]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net51),
    .QN(_0312_));
 DFFHQNx2_ASAP7_75t_R \REG[56]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net52),
    .QN(_0313_));
 DFFHQNx2_ASAP7_75t_R \REG[57]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(net53),
    .QN(_0314_));
 DFFHQNx2_ASAP7_75t_R \REG[58]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(net54),
    .QN(_0315_));
 DFFHQNx2_ASAP7_75t_R \REG[59]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net55),
    .QN(_0316_));
 DFFHQNx2_ASAP7_75t_R \REG[5]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(net56),
    .QN(_0262_));
 DFFHQNx2_ASAP7_75t_R \REG[60]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net57),
    .QN(_0317_));
 DFFHQNx2_ASAP7_75t_R \REG[61]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net58),
    .QN(_0318_));
 DFFHQNx2_ASAP7_75t_R \REG[62]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net59),
    .QN(_0319_));
 DFFHQNx2_ASAP7_75t_R \REG[63]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(net60),
    .QN(_0320_));
 DFFHQNx2_ASAP7_75t_R \REG[6]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net61),
    .QN(_0263_));
 DFFHQNx2_ASAP7_75t_R \REG[7]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(net62),
    .QN(_0264_));
 DFFHQNx2_ASAP7_75t_R \REG[8]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net63),
    .QN(_0265_));
 DFFHQNx2_ASAP7_75t_R \REG[9]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(net64),
    .QN(_0266_));
 DFFHQNx2_ASAP7_75t_R \REG_1[0]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(net65),
    .QN(_0449_));
 DFFHQNx2_ASAP7_75t_R \REG_1[10]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net66),
    .QN(_0459_));
 DFFHQNx2_ASAP7_75t_R \REG_1[11]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net67),
    .QN(_0460_));
 DFFHQNx2_ASAP7_75t_R \REG_1[12]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(net68),
    .QN(_0461_));
 DFFHQNx2_ASAP7_75t_R \REG_1[13]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net69),
    .QN(_0462_));
 DFFHQNx2_ASAP7_75t_R \REG_1[14]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net70),
    .QN(_0463_));
 DFFHQNx2_ASAP7_75t_R \REG_1[15]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net71),
    .QN(_0464_));
 DFFHQNx2_ASAP7_75t_R \REG_1[16]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net72),
    .QN(_0465_));
 DFFHQNx2_ASAP7_75t_R \REG_1[17]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net73),
    .QN(_0466_));
 DFFHQNx2_ASAP7_75t_R \REG_1[18]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net74),
    .QN(_0467_));
 DFFHQNx2_ASAP7_75t_R \REG_1[19]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(net75),
    .QN(_0468_));
 DFFHQNx2_ASAP7_75t_R \REG_1[1]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net76),
    .QN(_0450_));
 DFFHQNx2_ASAP7_75t_R \REG_1[20]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net77),
    .QN(_0469_));
 DFFHQNx2_ASAP7_75t_R \REG_1[21]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net78),
    .QN(_0470_));
 DFFHQNx2_ASAP7_75t_R \REG_1[22]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net79),
    .QN(_0471_));
 DFFHQNx2_ASAP7_75t_R \REG_1[23]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net80),
    .QN(_0472_));
 DFFHQNx2_ASAP7_75t_R \REG_1[24]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net81),
    .QN(_0473_));
 DFFHQNx2_ASAP7_75t_R \REG_1[25]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net82),
    .QN(_0474_));
 DFFHQNx2_ASAP7_75t_R \REG_1[26]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net83),
    .QN(_0475_));
 DFFHQNx2_ASAP7_75t_R \REG_1[27]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net84),
    .QN(_0476_));
 DFFHQNx2_ASAP7_75t_R \REG_1[28]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net85),
    .QN(_0477_));
 DFFHQNx2_ASAP7_75t_R \REG_1[29]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net86),
    .QN(_0478_));
 DFFHQNx2_ASAP7_75t_R \REG_1[2]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net87),
    .QN(_0451_));
 DFFHQNx2_ASAP7_75t_R \REG_1[30]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net88),
    .QN(_0479_));
 DFFHQNx2_ASAP7_75t_R \REG_1[31]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net89),
    .QN(_0480_));
 DFFHQNx2_ASAP7_75t_R \REG_1[32]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net90),
    .QN(_0481_));
 DFFHQNx2_ASAP7_75t_R \REG_1[33]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net91),
    .QN(_0482_));
 DFFHQNx2_ASAP7_75t_R \REG_1[34]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net92),
    .QN(_0483_));
 DFFHQNx2_ASAP7_75t_R \REG_1[35]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net93),
    .QN(_0484_));
 DFFHQNx2_ASAP7_75t_R \REG_1[36]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net94),
    .QN(_0485_));
 DFFHQNx2_ASAP7_75t_R \REG_1[37]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net95),
    .QN(_0486_));
 DFFHQNx2_ASAP7_75t_R \REG_1[38]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net96),
    .QN(_0487_));
 DFFHQNx2_ASAP7_75t_R \REG_1[39]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net97),
    .QN(_0488_));
 DFFHQNx2_ASAP7_75t_R \REG_1[3]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net98),
    .QN(_0452_));
 DFFHQNx2_ASAP7_75t_R \REG_1[40]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net99),
    .QN(_0489_));
 DFFHQNx2_ASAP7_75t_R \REG_1[41]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net100),
    .QN(_0490_));
 DFFHQNx2_ASAP7_75t_R \REG_1[42]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net101),
    .QN(_0491_));
 DFFHQNx2_ASAP7_75t_R \REG_1[43]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net102),
    .QN(_0492_));
 DFFHQNx2_ASAP7_75t_R \REG_1[44]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net103),
    .QN(_0493_));
 DFFHQNx2_ASAP7_75t_R \REG_1[45]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(net104),
    .QN(_0494_));
 DFFHQNx2_ASAP7_75t_R \REG_1[46]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net105),
    .QN(_0495_));
 DFFHQNx2_ASAP7_75t_R \REG_1[47]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net106),
    .QN(_0496_));
 DFFHQNx2_ASAP7_75t_R \REG_1[48]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net107),
    .QN(_0497_));
 DFFHQNx2_ASAP7_75t_R \REG_1[49]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net108),
    .QN(_0498_));
 DFFHQNx2_ASAP7_75t_R \REG_1[4]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net109),
    .QN(_0453_));
 DFFHQNx2_ASAP7_75t_R \REG_1[50]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net110),
    .QN(_0499_));
 DFFHQNx2_ASAP7_75t_R \REG_1[51]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net111),
    .QN(_0500_));
 DFFHQNx2_ASAP7_75t_R \REG_1[52]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net112),
    .QN(_0501_));
 DFFHQNx2_ASAP7_75t_R \REG_1[53]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net113),
    .QN(_0502_));
 DFFHQNx2_ASAP7_75t_R \REG_1[54]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net114),
    .QN(_0503_));
 DFFHQNx2_ASAP7_75t_R \REG_1[55]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net115),
    .QN(_0504_));
 DFFHQNx2_ASAP7_75t_R \REG_1[56]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(net116),
    .QN(_0505_));
 DFFHQNx2_ASAP7_75t_R \REG_1[57]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net117),
    .QN(_0506_));
 DFFHQNx2_ASAP7_75t_R \REG_1[58]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net118),
    .QN(_0507_));
 DFFHQNx2_ASAP7_75t_R \REG_1[59]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net119),
    .QN(_0508_));
 DFFHQNx2_ASAP7_75t_R \REG_1[5]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(net120),
    .QN(_0454_));
 DFFHQNx2_ASAP7_75t_R \REG_1[60]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net121),
    .QN(_0509_));
 DFFHQNx2_ASAP7_75t_R \REG_1[61]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net122),
    .QN(_0510_));
 DFFHQNx2_ASAP7_75t_R \REG_1[62]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net123),
    .QN(_0511_));
 DFFHQNx2_ASAP7_75t_R \REG_1[63]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(net124),
    .QN(_0512_));
 DFFHQNx2_ASAP7_75t_R \REG_1[6]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(net125),
    .QN(_0455_));
 DFFHQNx2_ASAP7_75t_R \REG_1[7]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net126),
    .QN(_0456_));
 DFFHQNx2_ASAP7_75t_R \REG_1[8]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net127),
    .QN(_0457_));
 DFFHQNx2_ASAP7_75t_R \REG_1[9]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net128),
    .QN(_0458_));
 DFFHQNx2_ASAP7_75t_R \REG_2[0]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net129),
    .QN(_0385_));
 DFFHQNx2_ASAP7_75t_R \REG_2[10]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net130),
    .QN(_0395_));
 DFFHQNx2_ASAP7_75t_R \REG_2[11]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net131),
    .QN(_0396_));
 DFFHQNx2_ASAP7_75t_R \REG_2[12]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net132),
    .QN(_0397_));
 DFFHQNx2_ASAP7_75t_R \REG_2[13]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net133),
    .QN(_0398_));
 DFFHQNx2_ASAP7_75t_R \REG_2[14]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net134),
    .QN(_0399_));
 DFFHQNx2_ASAP7_75t_R \REG_2[15]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net135),
    .QN(_0400_));
 DFFHQNx2_ASAP7_75t_R \REG_2[16]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net136),
    .QN(_0401_));
 DFFHQNx2_ASAP7_75t_R \REG_2[17]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net137),
    .QN(_0402_));
 DFFHQNx2_ASAP7_75t_R \REG_2[18]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net138),
    .QN(_0403_));
 DFFHQNx2_ASAP7_75t_R \REG_2[19]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net139),
    .QN(_0404_));
 DFFHQNx2_ASAP7_75t_R \REG_2[1]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net140),
    .QN(_0386_));
 DFFHQNx2_ASAP7_75t_R \REG_2[20]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net141),
    .QN(_0405_));
 DFFHQNx2_ASAP7_75t_R \REG_2[21]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net142),
    .QN(_0406_));
 DFFHQNx2_ASAP7_75t_R \REG_2[22]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(net143),
    .QN(_0407_));
 DFFHQNx2_ASAP7_75t_R \REG_2[23]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net144),
    .QN(_0408_));
 DFFHQNx2_ASAP7_75t_R \REG_2[24]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net145),
    .QN(_0409_));
 DFFHQNx2_ASAP7_75t_R \REG_2[25]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net146),
    .QN(_0410_));
 DFFHQNx2_ASAP7_75t_R \REG_2[26]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net147),
    .QN(_0411_));
 DFFHQNx2_ASAP7_75t_R \REG_2[27]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net148),
    .QN(_0412_));
 DFFHQNx2_ASAP7_75t_R \REG_2[28]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net149),
    .QN(_0413_));
 DFFHQNx2_ASAP7_75t_R \REG_2[29]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net150),
    .QN(_0414_));
 DFFHQNx2_ASAP7_75t_R \REG_2[2]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net151),
    .QN(_0387_));
 DFFHQNx2_ASAP7_75t_R \REG_2[30]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net152),
    .QN(_0415_));
 DFFHQNx2_ASAP7_75t_R \REG_2[31]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net153),
    .QN(_0416_));
 DFFHQNx2_ASAP7_75t_R \REG_2[32]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net154),
    .QN(_0417_));
 DFFHQNx2_ASAP7_75t_R \REG_2[33]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net155),
    .QN(_0418_));
 DFFHQNx2_ASAP7_75t_R \REG_2[34]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net156),
    .QN(_0419_));
 DFFHQNx2_ASAP7_75t_R \REG_2[35]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net157),
    .QN(_0420_));
 DFFHQNx2_ASAP7_75t_R \REG_2[36]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net158),
    .QN(_0421_));
 DFFHQNx2_ASAP7_75t_R \REG_2[37]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net159),
    .QN(_0422_));
 DFFHQNx2_ASAP7_75t_R \REG_2[38]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net160),
    .QN(_0423_));
 DFFHQNx2_ASAP7_75t_R \REG_2[39]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net161),
    .QN(_0424_));
 DFFHQNx2_ASAP7_75t_R \REG_2[3]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net162),
    .QN(_0388_));
 DFFHQNx2_ASAP7_75t_R \REG_2[40]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net163),
    .QN(_0425_));
 DFFHQNx2_ASAP7_75t_R \REG_2[41]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net164),
    .QN(_0426_));
 DFFHQNx2_ASAP7_75t_R \REG_2[42]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net165),
    .QN(_0427_));
 DFFHQNx2_ASAP7_75t_R \REG_2[43]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net166),
    .QN(_0428_));
 DFFHQNx2_ASAP7_75t_R \REG_2[44]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net167),
    .QN(_0429_));
 DFFHQNx2_ASAP7_75t_R \REG_2[45]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net168),
    .QN(_0430_));
 DFFHQNx2_ASAP7_75t_R \REG_2[46]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net169),
    .QN(_0431_));
 DFFHQNx2_ASAP7_75t_R \REG_2[47]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net170),
    .QN(_0432_));
 DFFHQNx2_ASAP7_75t_R \REG_2[48]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net171),
    .QN(_0433_));
 DFFHQNx2_ASAP7_75t_R \REG_2[49]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(net172),
    .QN(_0434_));
 DFFHQNx2_ASAP7_75t_R \REG_2[4]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net173),
    .QN(_0389_));
 DFFHQNx2_ASAP7_75t_R \REG_2[50]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net174),
    .QN(_0435_));
 DFFHQNx2_ASAP7_75t_R \REG_2[51]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net175),
    .QN(_0436_));
 DFFHQNx2_ASAP7_75t_R \REG_2[52]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net176),
    .QN(_0437_));
 DFFHQNx2_ASAP7_75t_R \REG_2[53]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net177),
    .QN(_0438_));
 DFFHQNx2_ASAP7_75t_R \REG_2[54]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net178),
    .QN(_0439_));
 DFFHQNx2_ASAP7_75t_R \REG_2[55]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(net179),
    .QN(_0440_));
 DFFHQNx2_ASAP7_75t_R \REG_2[56]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net180),
    .QN(_0441_));
 DFFHQNx2_ASAP7_75t_R \REG_2[57]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(net181),
    .QN(_0442_));
 DFFHQNx2_ASAP7_75t_R \REG_2[58]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net182),
    .QN(_0443_));
 DFFHQNx2_ASAP7_75t_R \REG_2[59]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(net183),
    .QN(_0444_));
 DFFHQNx2_ASAP7_75t_R \REG_2[5]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net184),
    .QN(_0390_));
 DFFHQNx2_ASAP7_75t_R \REG_2[60]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(net185),
    .QN(_0445_));
 DFFHQNx2_ASAP7_75t_R \REG_2[61]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(net186),
    .QN(_0446_));
 DFFHQNx2_ASAP7_75t_R \REG_2[62]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(net187),
    .QN(_0447_));
 DFFHQNx2_ASAP7_75t_R \REG_2[63]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(net188),
    .QN(_0448_));
 DFFHQNx2_ASAP7_75t_R \REG_2[6]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net189),
    .QN(_0391_));
 DFFHQNx2_ASAP7_75t_R \REG_2[7]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(net190),
    .QN(_0392_));
 DFFHQNx2_ASAP7_75t_R \REG_2[8]$_DFF_P_  (.CLK(clknet_leaf_0_clock),
    .D(net191),
    .QN(_0393_));
 DFFHQNx2_ASAP7_75t_R \REG_2[9]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(net192),
    .QN(_0394_));
 DFFHQNx2_ASAP7_75t_R \REG_4[0]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net193),
    .QN(_0321_));
 DFFHQNx2_ASAP7_75t_R \REG_4[10]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net194),
    .QN(_0331_));
 DFFHQNx2_ASAP7_75t_R \REG_4[11]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net195),
    .QN(_0332_));
 DFFHQNx2_ASAP7_75t_R \REG_4[12]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net196),
    .QN(_0333_));
 DFFHQNx2_ASAP7_75t_R \REG_4[13]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net197),
    .QN(_0334_));
 DFFHQNx2_ASAP7_75t_R \REG_4[14]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net198),
    .QN(_0335_));
 DFFHQNx2_ASAP7_75t_R \REG_4[15]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net199),
    .QN(_0336_));
 DFFHQNx2_ASAP7_75t_R \REG_4[16]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net200),
    .QN(_0337_));
 DFFHQNx2_ASAP7_75t_R \REG_4[17]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net201),
    .QN(_0338_));
 DFFHQNx2_ASAP7_75t_R \REG_4[18]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net202),
    .QN(_0339_));
 DFFHQNx2_ASAP7_75t_R \REG_4[19]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net203),
    .QN(_0340_));
 DFFHQNx2_ASAP7_75t_R \REG_4[1]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net204),
    .QN(_0322_));
 DFFHQNx2_ASAP7_75t_R \REG_4[20]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net205),
    .QN(_0341_));
 DFFHQNx2_ASAP7_75t_R \REG_4[21]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net206),
    .QN(_0342_));
 DFFHQNx2_ASAP7_75t_R \REG_4[22]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net207),
    .QN(_0343_));
 DFFHQNx2_ASAP7_75t_R \REG_4[23]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net208),
    .QN(_0344_));
 DFFHQNx2_ASAP7_75t_R \REG_4[24]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net209),
    .QN(_0345_));
 DFFHQNx2_ASAP7_75t_R \REG_4[25]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net210),
    .QN(_0346_));
 DFFHQNx2_ASAP7_75t_R \REG_4[26]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net211),
    .QN(_0347_));
 DFFHQNx2_ASAP7_75t_R \REG_4[27]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net212),
    .QN(_0348_));
 DFFHQNx2_ASAP7_75t_R \REG_4[28]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net213),
    .QN(_0349_));
 DFFHQNx2_ASAP7_75t_R \REG_4[29]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net214),
    .QN(_0350_));
 DFFHQNx2_ASAP7_75t_R \REG_4[2]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(net215),
    .QN(_0323_));
 DFFHQNx2_ASAP7_75t_R \REG_4[30]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net216),
    .QN(_0351_));
 DFFHQNx2_ASAP7_75t_R \REG_4[31]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net217),
    .QN(_0352_));
 DFFHQNx2_ASAP7_75t_R \REG_4[32]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net218),
    .QN(_0353_));
 DFFHQNx2_ASAP7_75t_R \REG_4[33]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net219),
    .QN(_0354_));
 DFFHQNx2_ASAP7_75t_R \REG_4[34]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net220),
    .QN(_0355_));
 DFFHQNx2_ASAP7_75t_R \REG_4[35]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net221),
    .QN(_0356_));
 DFFHQNx2_ASAP7_75t_R \REG_4[36]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net222),
    .QN(_0357_));
 DFFHQNx2_ASAP7_75t_R \REG_4[37]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(net223),
    .QN(_0358_));
 DFFHQNx2_ASAP7_75t_R \REG_4[38]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net224),
    .QN(_0359_));
 DFFHQNx2_ASAP7_75t_R \REG_4[39]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net225),
    .QN(_0360_));
 DFFHQNx2_ASAP7_75t_R \REG_4[3]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net226),
    .QN(_0324_));
 DFFHQNx2_ASAP7_75t_R \REG_4[40]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net227),
    .QN(_0361_));
 DFFHQNx2_ASAP7_75t_R \REG_4[41]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net228),
    .QN(_0362_));
 DFFHQNx2_ASAP7_75t_R \REG_4[42]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net229),
    .QN(_0363_));
 DFFHQNx2_ASAP7_75t_R \REG_4[43]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net230),
    .QN(_0364_));
 DFFHQNx2_ASAP7_75t_R \REG_4[44]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net231),
    .QN(_0365_));
 DFFHQNx2_ASAP7_75t_R \REG_4[45]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(net232),
    .QN(_0366_));
 DFFHQNx2_ASAP7_75t_R \REG_4[46]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net233),
    .QN(_0367_));
 DFFHQNx2_ASAP7_75t_R \REG_4[47]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(net234),
    .QN(_0368_));
 DFFHQNx2_ASAP7_75t_R \REG_4[48]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net235),
    .QN(_0369_));
 DFFHQNx2_ASAP7_75t_R \REG_4[49]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net236),
    .QN(_0370_));
 DFFHQNx2_ASAP7_75t_R \REG_4[4]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net237),
    .QN(_0325_));
 DFFHQNx2_ASAP7_75t_R \REG_4[50]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net238),
    .QN(_0371_));
 DFFHQNx2_ASAP7_75t_R \REG_4[51]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net239),
    .QN(_0372_));
 DFFHQNx2_ASAP7_75t_R \REG_4[52]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net240),
    .QN(_0373_));
 DFFHQNx2_ASAP7_75t_R \REG_4[53]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(net241),
    .QN(_0374_));
 DFFHQNx2_ASAP7_75t_R \REG_4[54]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net242),
    .QN(_0375_));
 DFFHQNx2_ASAP7_75t_R \REG_4[55]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(net243),
    .QN(_0376_));
 DFFHQNx2_ASAP7_75t_R \REG_4[56]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(net244),
    .QN(_0377_));
 DFFHQNx2_ASAP7_75t_R \REG_4[57]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(net245),
    .QN(_0378_));
 DFFHQNx2_ASAP7_75t_R \REG_4[58]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(net246),
    .QN(_0379_));
 DFFHQNx2_ASAP7_75t_R \REG_4[59]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(net247),
    .QN(_0380_));
 DFFHQNx2_ASAP7_75t_R \REG_4[5]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net248),
    .QN(_0326_));
 DFFHQNx2_ASAP7_75t_R \REG_4[60]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(net249),
    .QN(_0381_));
 DFFHQNx2_ASAP7_75t_R \REG_4[61]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(net250),
    .QN(_0382_));
 DFFHQNx2_ASAP7_75t_R \REG_4[62]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(net251),
    .QN(_0383_));
 DFFHQNx2_ASAP7_75t_R \REG_4[63]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(net252),
    .QN(_0384_));
 DFFHQNx2_ASAP7_75t_R \REG_4[6]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(net253),
    .QN(_0327_));
 DFFHQNx2_ASAP7_75t_R \REG_4[7]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net254),
    .QN(_0328_));
 DFFHQNx2_ASAP7_75t_R \REG_4[8]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net255),
    .QN(_0329_));
 DFFHQNx2_ASAP7_75t_R \REG_4[9]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(net256),
    .QN(_0330_));
 NAND2x1_ASAP7_75t_R _0769_ (.A(_0319_),
    .B(_0447_),
    .Y(_0250_));
 NAND2x1_ASAP7_75t_R _0770_ (.A(_0320_),
    .B(_0448_),
    .Y(_0251_));
 NAND2x1_ASAP7_75t_R _0771_ (.A(_0321_),
    .B(_0385_),
    .Y(_0128_));
 NAND2x1_ASAP7_75t_R _0772_ (.A(_0322_),
    .B(_0386_),
    .Y(_0139_));
 NAND2x1_ASAP7_75t_R _0773_ (.A(_0323_),
    .B(_0387_),
    .Y(_0150_));
 NAND2x1_ASAP7_75t_R _0774_ (.A(_0324_),
    .B(_0388_),
    .Y(_0161_));
 NAND2x1_ASAP7_75t_R _0775_ (.A(_0325_),
    .B(_0389_),
    .Y(_0172_));
 NAND2x1_ASAP7_75t_R _0776_ (.A(_0326_),
    .B(_0390_),
    .Y(_0183_));
 NAND2x1_ASAP7_75t_R _0777_ (.A(_0327_),
    .B(_0391_),
    .Y(_0188_));
 NAND2x1_ASAP7_75t_R _0778_ (.A(_0328_),
    .B(_0392_),
    .Y(_0189_));
 NAND2x1_ASAP7_75t_R _0779_ (.A(_0329_),
    .B(_0393_),
    .Y(_0190_));
 NAND2x1_ASAP7_75t_R _0780_ (.A(_0330_),
    .B(_0394_),
    .Y(_0191_));
 NAND2x1_ASAP7_75t_R _0781_ (.A(_0331_),
    .B(_0395_),
    .Y(_0129_));
 NAND2x1_ASAP7_75t_R _0782_ (.A(_0332_),
    .B(_0396_),
    .Y(_0130_));
 NAND2x1_ASAP7_75t_R _0783_ (.A(_0333_),
    .B(_0397_),
    .Y(_0131_));
 NAND2x1_ASAP7_75t_R _0784_ (.A(_0334_),
    .B(_0398_),
    .Y(_0132_));
 NAND2x1_ASAP7_75t_R _0785_ (.A(_0335_),
    .B(_0399_),
    .Y(_0133_));
 NAND2x1_ASAP7_75t_R _0786_ (.A(_0336_),
    .B(_0400_),
    .Y(_0134_));
 NAND2x1_ASAP7_75t_R _0787_ (.A(_0337_),
    .B(_0401_),
    .Y(_0135_));
 NAND2x1_ASAP7_75t_R _0788_ (.A(_0338_),
    .B(_0402_),
    .Y(_0136_));
 NAND2x1_ASAP7_75t_R _0789_ (.A(_0339_),
    .B(_0403_),
    .Y(_0137_));
 NAND2x1_ASAP7_75t_R _0790_ (.A(_0340_),
    .B(_0404_),
    .Y(_0138_));
 NAND2x1_ASAP7_75t_R _0791_ (.A(_0341_),
    .B(_0405_),
    .Y(_0140_));
 NAND2x1_ASAP7_75t_R _0792_ (.A(_0342_),
    .B(_0406_),
    .Y(_0141_));
 NAND2x1_ASAP7_75t_R _0793_ (.A(_0343_),
    .B(_0407_),
    .Y(_0142_));
 NAND2x1_ASAP7_75t_R _0794_ (.A(_0344_),
    .B(_0408_),
    .Y(_0143_));
 NAND2x1_ASAP7_75t_R _0795_ (.A(_0345_),
    .B(_0409_),
    .Y(_0144_));
 NAND2x1_ASAP7_75t_R _0796_ (.A(_0346_),
    .B(_0410_),
    .Y(_0145_));
 NAND2x1_ASAP7_75t_R _0797_ (.A(_0347_),
    .B(_0411_),
    .Y(_0146_));
 NAND2x1_ASAP7_75t_R _0798_ (.A(_0348_),
    .B(_0412_),
    .Y(_0147_));
 NAND2x1_ASAP7_75t_R _0799_ (.A(_0349_),
    .B(_0413_),
    .Y(_0148_));
 NAND2x1_ASAP7_75t_R _0800_ (.A(_0350_),
    .B(_0414_),
    .Y(_0149_));
 NAND2x1_ASAP7_75t_R _0801_ (.A(_0351_),
    .B(_0415_),
    .Y(_0151_));
 NAND2x1_ASAP7_75t_R _0802_ (.A(_0352_),
    .B(_0416_),
    .Y(_0152_));
 NAND2x1_ASAP7_75t_R _0803_ (.A(_0353_),
    .B(_0417_),
    .Y(_0153_));
 NAND2x1_ASAP7_75t_R _0804_ (.A(_0354_),
    .B(_0418_),
    .Y(_0154_));
 NAND2x1_ASAP7_75t_R _0805_ (.A(_0355_),
    .B(_0419_),
    .Y(_0155_));
 NAND2x1_ASAP7_75t_R _0806_ (.A(_0356_),
    .B(_0420_),
    .Y(_0156_));
 NAND2x1_ASAP7_75t_R _0807_ (.A(_0357_),
    .B(_0421_),
    .Y(_0157_));
 NAND2x1_ASAP7_75t_R _0808_ (.A(_0358_),
    .B(_0422_),
    .Y(_0158_));
 NAND2x1_ASAP7_75t_R _0809_ (.A(_0359_),
    .B(_0423_),
    .Y(_0159_));
 NAND2x1_ASAP7_75t_R _0810_ (.A(_0360_),
    .B(_0424_),
    .Y(_0160_));
 NAND2x1_ASAP7_75t_R _0811_ (.A(_0361_),
    .B(_0425_),
    .Y(_0162_));
 NAND2x1_ASAP7_75t_R _0812_ (.A(_0362_),
    .B(_0426_),
    .Y(_0163_));
 NAND2x1_ASAP7_75t_R _0813_ (.A(_0363_),
    .B(_0427_),
    .Y(_0164_));
 NAND2x1_ASAP7_75t_R _0814_ (.A(_0364_),
    .B(_0428_),
    .Y(_0165_));
 NAND2x1_ASAP7_75t_R _0815_ (.A(_0365_),
    .B(_0429_),
    .Y(_0166_));
 NAND2x1_ASAP7_75t_R _0816_ (.A(_0366_),
    .B(_0430_),
    .Y(_0167_));
 NAND2x1_ASAP7_75t_R _0817_ (.A(_0367_),
    .B(_0431_),
    .Y(_0168_));
 NAND2x1_ASAP7_75t_R _0818_ (.A(_0368_),
    .B(_0432_),
    .Y(_0169_));
 NAND2x1_ASAP7_75t_R _0819_ (.A(_0369_),
    .B(_0433_),
    .Y(_0170_));
 NAND2x1_ASAP7_75t_R _0820_ (.A(_0370_),
    .B(_0434_),
    .Y(_0171_));
 NAND2x1_ASAP7_75t_R _0821_ (.A(_0371_),
    .B(_0435_),
    .Y(_0173_));
 NAND2x1_ASAP7_75t_R _0822_ (.A(_0372_),
    .B(_0436_),
    .Y(_0174_));
 NAND2x1_ASAP7_75t_R _0823_ (.A(_0373_),
    .B(_0437_),
    .Y(_0175_));
 NAND2x1_ASAP7_75t_R _0824_ (.A(_0374_),
    .B(_0438_),
    .Y(_0176_));
 NAND2x1_ASAP7_75t_R _0825_ (.A(_0375_),
    .B(_0439_),
    .Y(_0177_));
 NAND2x1_ASAP7_75t_R _0826_ (.A(_0376_),
    .B(_0440_),
    .Y(_0178_));
 NAND2x1_ASAP7_75t_R _0827_ (.A(_0377_),
    .B(_0441_),
    .Y(_0179_));
 NAND2x1_ASAP7_75t_R _0828_ (.A(_0378_),
    .B(_0442_),
    .Y(_0180_));
 NAND2x1_ASAP7_75t_R _0829_ (.A(_0379_),
    .B(_0443_),
    .Y(_0181_));
 NAND2x1_ASAP7_75t_R _0830_ (.A(_0380_),
    .B(_0444_),
    .Y(_0182_));
 NAND2x1_ASAP7_75t_R _0831_ (.A(_0381_),
    .B(_0445_),
    .Y(_0184_));
 NAND2x1_ASAP7_75t_R _0832_ (.A(_0382_),
    .B(_0446_),
    .Y(_0185_));
 NAND2x1_ASAP7_75t_R _0833_ (.A(_0383_),
    .B(_0447_),
    .Y(_0186_));
 NAND2x1_ASAP7_75t_R _0834_ (.A(_0384_),
    .B(_0448_),
    .Y(_0187_));
 NAND2x1_ASAP7_75t_R _0835_ (.A(_0321_),
    .B(_0449_),
    .Y(_0000_));
 NAND2x1_ASAP7_75t_R _0836_ (.A(_0322_),
    .B(_0450_),
    .Y(_0011_));
 NAND2x1_ASAP7_75t_R _0837_ (.A(_0323_),
    .B(_0451_),
    .Y(_0022_));
 NAND2x1_ASAP7_75t_R _0838_ (.A(_0324_),
    .B(_0452_),
    .Y(_0033_));
 NAND2x1_ASAP7_75t_R _0839_ (.A(_0325_),
    .B(_0453_),
    .Y(_0044_));
 NAND2x1_ASAP7_75t_R _0840_ (.A(_0326_),
    .B(_0454_),
    .Y(_0055_));
 NAND2x1_ASAP7_75t_R _0841_ (.A(_0327_),
    .B(_0455_),
    .Y(_0060_));
 NAND2x1_ASAP7_75t_R _0842_ (.A(_0328_),
    .B(_0456_),
    .Y(_0061_));
 NAND2x1_ASAP7_75t_R _0843_ (.A(_0329_),
    .B(_0457_),
    .Y(_0062_));
 NAND2x1_ASAP7_75t_R _0844_ (.A(_0330_),
    .B(_0458_),
    .Y(_0063_));
 NAND2x1_ASAP7_75t_R _0845_ (.A(_0331_),
    .B(_0459_),
    .Y(_0001_));
 NAND2x1_ASAP7_75t_R _0846_ (.A(_0332_),
    .B(_0460_),
    .Y(_0002_));
 NAND2x1_ASAP7_75t_R _0847_ (.A(_0333_),
    .B(_0461_),
    .Y(_0003_));
 NAND2x1_ASAP7_75t_R _0848_ (.A(_0334_),
    .B(_0462_),
    .Y(_0004_));
 NAND2x1_ASAP7_75t_R _0849_ (.A(_0335_),
    .B(_0463_),
    .Y(_0005_));
 NAND2x1_ASAP7_75t_R _0850_ (.A(_0336_),
    .B(_0464_),
    .Y(_0006_));
 NAND2x1_ASAP7_75t_R _0851_ (.A(_0337_),
    .B(_0465_),
    .Y(_0007_));
 NAND2x1_ASAP7_75t_R _0852_ (.A(_0338_),
    .B(_0466_),
    .Y(_0008_));
 NAND2x1_ASAP7_75t_R _0853_ (.A(_0339_),
    .B(_0467_),
    .Y(_0009_));
 NAND2x1_ASAP7_75t_R _0854_ (.A(_0340_),
    .B(_0468_),
    .Y(_0010_));
 NAND2x1_ASAP7_75t_R _0855_ (.A(_0341_),
    .B(_0469_),
    .Y(_0012_));
 NAND2x1_ASAP7_75t_R _0856_ (.A(_0342_),
    .B(_0470_),
    .Y(_0013_));
 NAND2x1_ASAP7_75t_R _0857_ (.A(_0343_),
    .B(_0471_),
    .Y(_0014_));
 NAND2x1_ASAP7_75t_R _0858_ (.A(_0344_),
    .B(_0472_),
    .Y(_0015_));
 NAND2x1_ASAP7_75t_R _0859_ (.A(_0345_),
    .B(_0473_),
    .Y(_0016_));
 NAND2x1_ASAP7_75t_R _0860_ (.A(_0346_),
    .B(_0474_),
    .Y(_0017_));
 NAND2x1_ASAP7_75t_R _0861_ (.A(_0347_),
    .B(_0475_),
    .Y(_0018_));
 NAND2x1_ASAP7_75t_R _0862_ (.A(_0348_),
    .B(_0476_),
    .Y(_0019_));
 NAND2x1_ASAP7_75t_R _0863_ (.A(_0349_),
    .B(_0477_),
    .Y(_0020_));
 NAND2x1_ASAP7_75t_R _0864_ (.A(_0350_),
    .B(_0478_),
    .Y(_0021_));
 NAND2x1_ASAP7_75t_R _0865_ (.A(_0351_),
    .B(_0479_),
    .Y(_0023_));
 NAND2x1_ASAP7_75t_R _0866_ (.A(_0352_),
    .B(_0480_),
    .Y(_0024_));
 NAND2x1_ASAP7_75t_R _0867_ (.A(_0353_),
    .B(_0481_),
    .Y(_0025_));
 NAND2x1_ASAP7_75t_R _0868_ (.A(_0354_),
    .B(_0482_),
    .Y(_0026_));
 NAND2x1_ASAP7_75t_R _0869_ (.A(_0355_),
    .B(_0483_),
    .Y(_0027_));
 NAND2x1_ASAP7_75t_R _0870_ (.A(_0356_),
    .B(_0484_),
    .Y(_0028_));
 NAND2x1_ASAP7_75t_R _0871_ (.A(_0357_),
    .B(_0485_),
    .Y(_0029_));
 NAND2x1_ASAP7_75t_R _0872_ (.A(_0358_),
    .B(_0486_),
    .Y(_0030_));
 NAND2x1_ASAP7_75t_R _0873_ (.A(_0359_),
    .B(_0487_),
    .Y(_0031_));
 NAND2x1_ASAP7_75t_R _0874_ (.A(_0360_),
    .B(_0488_),
    .Y(_0032_));
 NAND2x1_ASAP7_75t_R _0875_ (.A(_0361_),
    .B(_0489_),
    .Y(_0034_));
 NAND2x1_ASAP7_75t_R _0876_ (.A(_0362_),
    .B(_0490_),
    .Y(_0035_));
 NAND2x1_ASAP7_75t_R _0877_ (.A(_0363_),
    .B(_0491_),
    .Y(_0036_));
 NAND2x1_ASAP7_75t_R _0878_ (.A(_0364_),
    .B(_0492_),
    .Y(_0037_));
 NAND2x1_ASAP7_75t_R _0879_ (.A(_0365_),
    .B(_0493_),
    .Y(_0038_));
 NAND2x1_ASAP7_75t_R _0880_ (.A(_0366_),
    .B(_0494_),
    .Y(_0039_));
 NAND2x1_ASAP7_75t_R _0881_ (.A(_0367_),
    .B(_0495_),
    .Y(_0040_));
 NAND2x1_ASAP7_75t_R _0882_ (.A(_0368_),
    .B(_0496_),
    .Y(_0041_));
 NAND2x1_ASAP7_75t_R _0883_ (.A(_0369_),
    .B(_0497_),
    .Y(_0042_));
 NAND2x1_ASAP7_75t_R _0884_ (.A(_0370_),
    .B(_0498_),
    .Y(_0043_));
 NAND2x1_ASAP7_75t_R _0885_ (.A(_0371_),
    .B(_0499_),
    .Y(_0045_));
 NAND2x1_ASAP7_75t_R _0886_ (.A(_0372_),
    .B(_0500_),
    .Y(_0046_));
 NAND2x1_ASAP7_75t_R _0887_ (.A(_0373_),
    .B(_0501_),
    .Y(_0047_));
 NAND2x1_ASAP7_75t_R _0888_ (.A(_0374_),
    .B(_0502_),
    .Y(_0048_));
 NAND2x1_ASAP7_75t_R _0889_ (.A(_0375_),
    .B(_0503_),
    .Y(_0049_));
 NAND2x1_ASAP7_75t_R _0890_ (.A(_0376_),
    .B(_0504_),
    .Y(_0050_));
 NAND2x1_ASAP7_75t_R _0891_ (.A(_0377_),
    .B(_0505_),
    .Y(_0051_));
 NAND2x1_ASAP7_75t_R _0892_ (.A(_0378_),
    .B(_0506_),
    .Y(_0052_));
 NAND2x1_ASAP7_75t_R _0893_ (.A(_0379_),
    .B(_0507_),
    .Y(_0053_));
 NAND2x1_ASAP7_75t_R _0894_ (.A(_0380_),
    .B(_0508_),
    .Y(_0054_));
 NAND2x1_ASAP7_75t_R _0895_ (.A(_0381_),
    .B(_0509_),
    .Y(_0056_));
 NAND2x1_ASAP7_75t_R _0896_ (.A(_0382_),
    .B(_0510_),
    .Y(_0057_));
 NAND2x1_ASAP7_75t_R _0897_ (.A(_0383_),
    .B(_0511_),
    .Y(_0058_));
 NAND2x1_ASAP7_75t_R _0898_ (.A(_0384_),
    .B(_0512_),
    .Y(_0059_));
 NAND2x1_ASAP7_75t_R _0899_ (.A(_0257_),
    .B(_0449_),
    .Y(_0064_));
 NAND2x1_ASAP7_75t_R _0900_ (.A(_0258_),
    .B(_0450_),
    .Y(_0075_));
 NAND2x1_ASAP7_75t_R _0901_ (.A(_0259_),
    .B(_0451_),
    .Y(_0086_));
 NAND2x1_ASAP7_75t_R _0902_ (.A(_0260_),
    .B(_0452_),
    .Y(_0097_));
 NAND2x1_ASAP7_75t_R _0903_ (.A(_0261_),
    .B(_0453_),
    .Y(_0108_));
 NAND2x1_ASAP7_75t_R _0904_ (.A(_0262_),
    .B(_0454_),
    .Y(_0119_));
 NAND2x1_ASAP7_75t_R _0905_ (.A(_0263_),
    .B(_0455_),
    .Y(_0124_));
 NAND2x1_ASAP7_75t_R _0906_ (.A(_0264_),
    .B(_0456_),
    .Y(_0125_));
 NAND2x1_ASAP7_75t_R _0907_ (.A(_0265_),
    .B(_0457_),
    .Y(_0126_));
 NAND2x1_ASAP7_75t_R _0908_ (.A(_0266_),
    .B(_0458_),
    .Y(_0127_));
 NAND2x1_ASAP7_75t_R _0909_ (.A(_0267_),
    .B(_0459_),
    .Y(_0065_));
 NAND2x1_ASAP7_75t_R _0910_ (.A(_0268_),
    .B(_0460_),
    .Y(_0066_));
 NAND2x1_ASAP7_75t_R _0911_ (.A(_0269_),
    .B(_0461_),
    .Y(_0067_));
 NAND2x1_ASAP7_75t_R _0912_ (.A(_0270_),
    .B(_0462_),
    .Y(_0068_));
 NAND2x1_ASAP7_75t_R _0913_ (.A(_0271_),
    .B(_0463_),
    .Y(_0069_));
 NAND2x1_ASAP7_75t_R _0914_ (.A(_0272_),
    .B(_0464_),
    .Y(_0070_));
 NAND2x1_ASAP7_75t_R _0915_ (.A(_0273_),
    .B(_0465_),
    .Y(_0071_));
 NAND2x1_ASAP7_75t_R _0916_ (.A(_0274_),
    .B(_0466_),
    .Y(_0072_));
 NAND2x1_ASAP7_75t_R _0917_ (.A(_0275_),
    .B(_0467_),
    .Y(_0073_));
 NAND2x1_ASAP7_75t_R _0918_ (.A(_0276_),
    .B(_0468_),
    .Y(_0074_));
 NAND2x1_ASAP7_75t_R _0919_ (.A(_0277_),
    .B(_0469_),
    .Y(_0076_));
 NAND2x1_ASAP7_75t_R _0920_ (.A(_0278_),
    .B(_0470_),
    .Y(_0077_));
 NAND2x1_ASAP7_75t_R _0921_ (.A(_0279_),
    .B(_0471_),
    .Y(_0078_));
 NAND2x1_ASAP7_75t_R _0922_ (.A(_0280_),
    .B(_0472_),
    .Y(_0079_));
 NAND2x1_ASAP7_75t_R _0923_ (.A(_0281_),
    .B(_0473_),
    .Y(_0080_));
 NAND2x1_ASAP7_75t_R _0924_ (.A(_0282_),
    .B(_0474_),
    .Y(_0081_));
 NAND2x1_ASAP7_75t_R _0925_ (.A(_0283_),
    .B(_0475_),
    .Y(_0082_));
 NAND2x1_ASAP7_75t_R _0926_ (.A(_0284_),
    .B(_0476_),
    .Y(_0083_));
 NAND2x1_ASAP7_75t_R _0927_ (.A(_0285_),
    .B(_0477_),
    .Y(_0084_));
 NAND2x1_ASAP7_75t_R _0928_ (.A(_0286_),
    .B(_0478_),
    .Y(_0085_));
 NAND2x1_ASAP7_75t_R _0929_ (.A(_0287_),
    .B(_0479_),
    .Y(_0087_));
 NAND2x1_ASAP7_75t_R _0930_ (.A(_0288_),
    .B(_0480_),
    .Y(_0088_));
 NAND2x1_ASAP7_75t_R _0931_ (.A(_0289_),
    .B(_0481_),
    .Y(_0089_));
 NAND2x1_ASAP7_75t_R _0932_ (.A(_0290_),
    .B(_0482_),
    .Y(_0090_));
 NAND2x1_ASAP7_75t_R _0933_ (.A(_0291_),
    .B(_0483_),
    .Y(_0091_));
 NAND2x1_ASAP7_75t_R _0934_ (.A(_0292_),
    .B(_0484_),
    .Y(_0092_));
 NAND2x1_ASAP7_75t_R _0935_ (.A(_0293_),
    .B(_0485_),
    .Y(_0093_));
 NAND2x1_ASAP7_75t_R _0936_ (.A(_0294_),
    .B(_0486_),
    .Y(_0094_));
 NAND2x1_ASAP7_75t_R _0937_ (.A(_0295_),
    .B(_0487_),
    .Y(_0095_));
 NAND2x1_ASAP7_75t_R _0938_ (.A(_0296_),
    .B(_0488_),
    .Y(_0096_));
 NAND2x1_ASAP7_75t_R _0939_ (.A(_0297_),
    .B(_0489_),
    .Y(_0098_));
 NAND2x1_ASAP7_75t_R _0940_ (.A(_0298_),
    .B(_0490_),
    .Y(_0099_));
 NAND2x1_ASAP7_75t_R _0941_ (.A(_0299_),
    .B(_0491_),
    .Y(_0100_));
 NAND2x1_ASAP7_75t_R _0942_ (.A(_0300_),
    .B(_0492_),
    .Y(_0101_));
 NAND2x1_ASAP7_75t_R _0943_ (.A(_0301_),
    .B(_0493_),
    .Y(_0102_));
 NAND2x1_ASAP7_75t_R _0944_ (.A(_0302_),
    .B(_0494_),
    .Y(_0103_));
 NAND2x1_ASAP7_75t_R _0945_ (.A(_0303_),
    .B(_0495_),
    .Y(_0104_));
 NAND2x1_ASAP7_75t_R _0946_ (.A(_0304_),
    .B(_0496_),
    .Y(_0105_));
 NAND2x1_ASAP7_75t_R _0947_ (.A(_0305_),
    .B(_0497_),
    .Y(_0106_));
 NAND2x1_ASAP7_75t_R _0948_ (.A(_0306_),
    .B(_0498_),
    .Y(_0107_));
 NAND2x1_ASAP7_75t_R _0949_ (.A(_0307_),
    .B(_0499_),
    .Y(_0109_));
 NAND2x1_ASAP7_75t_R _0950_ (.A(_0308_),
    .B(_0500_),
    .Y(_0110_));
 NAND2x1_ASAP7_75t_R _0951_ (.A(_0309_),
    .B(_0501_),
    .Y(_0111_));
 NAND2x1_ASAP7_75t_R _0952_ (.A(_0310_),
    .B(_0502_),
    .Y(_0112_));
 NAND2x1_ASAP7_75t_R _0953_ (.A(_0311_),
    .B(_0503_),
    .Y(_0113_));
 NAND2x1_ASAP7_75t_R _0954_ (.A(_0312_),
    .B(_0504_),
    .Y(_0114_));
 NAND2x1_ASAP7_75t_R _0955_ (.A(_0313_),
    .B(_0505_),
    .Y(_0115_));
 NAND2x1_ASAP7_75t_R _0956_ (.A(_0314_),
    .B(_0506_),
    .Y(_0116_));
 NAND2x1_ASAP7_75t_R _0957_ (.A(_0315_),
    .B(_0507_),
    .Y(_0117_));
 NAND2x1_ASAP7_75t_R _0958_ (.A(_0316_),
    .B(_0508_),
    .Y(_0118_));
 NAND2x1_ASAP7_75t_R _0959_ (.A(_0317_),
    .B(_0509_),
    .Y(_0120_));
 NAND2x1_ASAP7_75t_R _0960_ (.A(_0318_),
    .B(_0510_),
    .Y(_0121_));
 NAND2x1_ASAP7_75t_R _0961_ (.A(_0319_),
    .B(_0511_),
    .Y(_0122_));
 NAND2x1_ASAP7_75t_R _0962_ (.A(_0320_),
    .B(_0512_),
    .Y(_0123_));
 NAND2x1_ASAP7_75t_R _0963_ (.A(_0257_),
    .B(_0385_),
    .Y(_0192_));
 NAND2x1_ASAP7_75t_R _0964_ (.A(_0258_),
    .B(_0386_),
    .Y(_0203_));
 NAND2x1_ASAP7_75t_R _0965_ (.A(_0259_),
    .B(_0387_),
    .Y(_0214_));
 NAND2x1_ASAP7_75t_R _0966_ (.A(_0260_),
    .B(_0388_),
    .Y(_0225_));
 NAND2x1_ASAP7_75t_R _0967_ (.A(_0261_),
    .B(_0389_),
    .Y(_0236_));
 NAND2x1_ASAP7_75t_R _0968_ (.A(_0262_),
    .B(_0390_),
    .Y(_0247_));
 NAND2x1_ASAP7_75t_R _0969_ (.A(_0263_),
    .B(_0391_),
    .Y(_0252_));
 NAND2x1_ASAP7_75t_R _0970_ (.A(_0264_),
    .B(_0392_),
    .Y(_0253_));
 NAND2x1_ASAP7_75t_R _0971_ (.A(_0265_),
    .B(_0393_),
    .Y(_0254_));
 NAND2x1_ASAP7_75t_R _0972_ (.A(_0266_),
    .B(_0394_),
    .Y(_0255_));
 NAND2x1_ASAP7_75t_R _0973_ (.A(_0267_),
    .B(_0395_),
    .Y(_0193_));
 NAND2x1_ASAP7_75t_R _0974_ (.A(_0268_),
    .B(_0396_),
    .Y(_0194_));
 NAND2x1_ASAP7_75t_R _0975_ (.A(_0269_),
    .B(_0397_),
    .Y(_0195_));
 NAND2x1_ASAP7_75t_R _0976_ (.A(_0270_),
    .B(_0398_),
    .Y(_0196_));
 NAND2x1_ASAP7_75t_R _0977_ (.A(_0271_),
    .B(_0399_),
    .Y(_0197_));
 NAND2x1_ASAP7_75t_R _0978_ (.A(_0272_),
    .B(_0400_),
    .Y(_0198_));
 NAND2x1_ASAP7_75t_R _0979_ (.A(_0273_),
    .B(_0401_),
    .Y(_0199_));
 NAND2x1_ASAP7_75t_R _0980_ (.A(_0274_),
    .B(_0402_),
    .Y(_0200_));
 NAND2x1_ASAP7_75t_R _0981_ (.A(_0275_),
    .B(_0403_),
    .Y(_0201_));
 NAND2x1_ASAP7_75t_R _0982_ (.A(_0276_),
    .B(_0404_),
    .Y(_0202_));
 NAND2x1_ASAP7_75t_R _0983_ (.A(_0277_),
    .B(_0405_),
    .Y(_0204_));
 NAND2x1_ASAP7_75t_R _0984_ (.A(_0278_),
    .B(_0406_),
    .Y(_0205_));
 NAND2x1_ASAP7_75t_R _0985_ (.A(_0279_),
    .B(_0407_),
    .Y(_0206_));
 NAND2x1_ASAP7_75t_R _0986_ (.A(_0280_),
    .B(_0408_),
    .Y(_0207_));
 NAND2x1_ASAP7_75t_R _0987_ (.A(_0281_),
    .B(_0409_),
    .Y(_0208_));
 NAND2x1_ASAP7_75t_R _0988_ (.A(_0282_),
    .B(_0410_),
    .Y(_0209_));
 NAND2x1_ASAP7_75t_R _0989_ (.A(_0283_),
    .B(_0411_),
    .Y(_0210_));
 NAND2x1_ASAP7_75t_R _0990_ (.A(_0284_),
    .B(_0412_),
    .Y(_0211_));
 NAND2x1_ASAP7_75t_R _0991_ (.A(_0285_),
    .B(_0413_),
    .Y(_0212_));
 NAND2x1_ASAP7_75t_R _0992_ (.A(_0286_),
    .B(_0414_),
    .Y(_0213_));
 NAND2x1_ASAP7_75t_R _0993_ (.A(_0287_),
    .B(_0415_),
    .Y(_0215_));
 NAND2x1_ASAP7_75t_R _0994_ (.A(_0288_),
    .B(_0416_),
    .Y(_0216_));
 NAND2x1_ASAP7_75t_R _0995_ (.A(_0289_),
    .B(_0417_),
    .Y(_0217_));
 NAND2x1_ASAP7_75t_R _0996_ (.A(_0290_),
    .B(_0418_),
    .Y(_0218_));
 NAND2x1_ASAP7_75t_R _0997_ (.A(_0291_),
    .B(_0419_),
    .Y(_0219_));
 NAND2x1_ASAP7_75t_R _0998_ (.A(_0292_),
    .B(_0420_),
    .Y(_0220_));
 NAND2x1_ASAP7_75t_R _0999_ (.A(_0293_),
    .B(_0421_),
    .Y(_0221_));
 NAND2x1_ASAP7_75t_R _1000_ (.A(_0294_),
    .B(_0422_),
    .Y(_0222_));
 NAND2x1_ASAP7_75t_R _1001_ (.A(_0295_),
    .B(_0423_),
    .Y(_0223_));
 NAND2x1_ASAP7_75t_R _1002_ (.A(_0296_),
    .B(_0424_),
    .Y(_0224_));
 NAND2x1_ASAP7_75t_R _1003_ (.A(_0297_),
    .B(_0425_),
    .Y(_0226_));
 NAND2x1_ASAP7_75t_R _1004_ (.A(_0298_),
    .B(_0426_),
    .Y(_0227_));
 NAND2x1_ASAP7_75t_R _1005_ (.A(_0299_),
    .B(_0427_),
    .Y(_0228_));
 NAND2x1_ASAP7_75t_R _1006_ (.A(_0300_),
    .B(_0428_),
    .Y(_0229_));
 NAND2x1_ASAP7_75t_R _1007_ (.A(_0301_),
    .B(_0429_),
    .Y(_0230_));
 NAND2x1_ASAP7_75t_R _1008_ (.A(_0302_),
    .B(_0430_),
    .Y(_0231_));
 NAND2x1_ASAP7_75t_R _1009_ (.A(_0303_),
    .B(_0431_),
    .Y(_0232_));
 NAND2x1_ASAP7_75t_R _1010_ (.A(_0304_),
    .B(_0432_),
    .Y(_0233_));
 NAND2x1_ASAP7_75t_R _1011_ (.A(_0305_),
    .B(_0433_),
    .Y(_0234_));
 NAND2x1_ASAP7_75t_R _1012_ (.A(_0306_),
    .B(_0434_),
    .Y(_0235_));
 NAND2x1_ASAP7_75t_R _1013_ (.A(_0307_),
    .B(_0435_),
    .Y(_0237_));
 NAND2x1_ASAP7_75t_R _1014_ (.A(_0308_),
    .B(_0436_),
    .Y(_0238_));
 NAND2x1_ASAP7_75t_R _1015_ (.A(_0309_),
    .B(_0437_),
    .Y(_0239_));
 NAND2x1_ASAP7_75t_R _1016_ (.A(_0310_),
    .B(_0438_),
    .Y(_0240_));
 NAND2x1_ASAP7_75t_R _1017_ (.A(_0311_),
    .B(_0439_),
    .Y(_0241_));
 NAND2x1_ASAP7_75t_R _1018_ (.A(_0312_),
    .B(_0440_),
    .Y(_0242_));
 NAND2x1_ASAP7_75t_R _1019_ (.A(_0313_),
    .B(_0441_),
    .Y(_0243_));
 NAND2x1_ASAP7_75t_R _1020_ (.A(_0314_),
    .B(_0442_),
    .Y(_0244_));
 NAND2x1_ASAP7_75t_R _1021_ (.A(_0315_),
    .B(_0443_),
    .Y(_0245_));
 NAND2x1_ASAP7_75t_R _1022_ (.A(_0316_),
    .B(_0444_),
    .Y(_0246_));
 NAND2x1_ASAP7_75t_R _1023_ (.A(_0317_),
    .B(_0445_),
    .Y(_0248_));
 NAND2x1_ASAP7_75t_R _1024_ (.A(_0318_),
    .B(_0446_),
    .Y(_0249_));
 INVx1_ASAP7_75t_R _1025_ (.A(_0256_),
    .Y(net261));
 INVx2_ASAP7_75t_R _1026_ (.A(_0513_),
    .Y(net265));
 INVx1_ASAP7_75t_R _1027_ (.A(_0514_),
    .Y(net341));
 INVx1_ASAP7_75t_R _1028_ (.A(_0515_),
    .Y(net352));
 INVx1_ASAP7_75t_R _1029_ (.A(_0516_),
    .Y(net363));
 INVx1_ASAP7_75t_R _1030_ (.A(_0517_),
    .Y(net374));
 INVx1_ASAP7_75t_R _1031_ (.A(_0518_),
    .Y(net385));
 INVx1_ASAP7_75t_R _1032_ (.A(_0519_),
    .Y(net390));
 INVx1_ASAP7_75t_R _1033_ (.A(_0520_),
    .Y(net391));
 INVx1_ASAP7_75t_R _1034_ (.A(_0521_),
    .Y(net392));
 INVx1_ASAP7_75t_R _1035_ (.A(_0522_),
    .Y(net393));
 INVx1_ASAP7_75t_R _1036_ (.A(_0523_),
    .Y(net331));
 INVx1_ASAP7_75t_R _1037_ (.A(_0524_),
    .Y(net332));
 INVx1_ASAP7_75t_R _1038_ (.A(_0525_),
    .Y(net333));
 INVx1_ASAP7_75t_R _1039_ (.A(_0526_),
    .Y(net334));
 INVx1_ASAP7_75t_R _1040_ (.A(_0527_),
    .Y(net335));
 INVx1_ASAP7_75t_R _1041_ (.A(_0528_),
    .Y(net336));
 INVx1_ASAP7_75t_R _1042_ (.A(_0529_),
    .Y(net337));
 INVx1_ASAP7_75t_R _1043_ (.A(_0530_),
    .Y(net338));
 INVx1_ASAP7_75t_R _1044_ (.A(_0531_),
    .Y(net339));
 INVx1_ASAP7_75t_R _1045_ (.A(_0532_),
    .Y(net340));
 INVx1_ASAP7_75t_R _1046_ (.A(_0533_),
    .Y(net342));
 INVx1_ASAP7_75t_R _1047_ (.A(_0534_),
    .Y(net343));
 INVx1_ASAP7_75t_R _1048_ (.A(_0535_),
    .Y(net344));
 INVx1_ASAP7_75t_R _1049_ (.A(_0536_),
    .Y(net345));
 INVx1_ASAP7_75t_R _1050_ (.A(_0537_),
    .Y(net346));
 INVx1_ASAP7_75t_R _1051_ (.A(_0538_),
    .Y(net347));
 INVx1_ASAP7_75t_R _1052_ (.A(_0539_),
    .Y(net348));
 INVx1_ASAP7_75t_R _1053_ (.A(_0540_),
    .Y(net349));
 INVx1_ASAP7_75t_R _1054_ (.A(_0541_),
    .Y(net350));
 INVx1_ASAP7_75t_R _1055_ (.A(_0542_),
    .Y(net351));
 INVx1_ASAP7_75t_R _1056_ (.A(_0543_),
    .Y(net353));
 INVx1_ASAP7_75t_R _1057_ (.A(_0544_),
    .Y(net354));
 INVx1_ASAP7_75t_R _1058_ (.A(_0545_),
    .Y(net355));
 INVx1_ASAP7_75t_R _1059_ (.A(_0546_),
    .Y(net356));
 INVx1_ASAP7_75t_R _1060_ (.A(_0547_),
    .Y(net357));
 INVx1_ASAP7_75t_R _1061_ (.A(_0548_),
    .Y(net358));
 INVx1_ASAP7_75t_R _1062_ (.A(_0549_),
    .Y(net359));
 INVx1_ASAP7_75t_R _1063_ (.A(_0550_),
    .Y(net360));
 INVx1_ASAP7_75t_R _1064_ (.A(_0551_),
    .Y(net361));
 INVx1_ASAP7_75t_R _1065_ (.A(_0552_),
    .Y(net362));
 INVx1_ASAP7_75t_R _1066_ (.A(_0553_),
    .Y(net364));
 INVx1_ASAP7_75t_R _1067_ (.A(_0554_),
    .Y(net365));
 INVx2_ASAP7_75t_R _1068_ (.A(_0555_),
    .Y(net366));
 INVx1_ASAP7_75t_R _1069_ (.A(_0556_),
    .Y(net367));
 INVx2_ASAP7_75t_R _1070_ (.A(_0557_),
    .Y(net368));
 INVx1_ASAP7_75t_R _1071_ (.A(_0558_),
    .Y(net369));
 INVx1_ASAP7_75t_R _1072_ (.A(_0559_),
    .Y(net370));
 INVx1_ASAP7_75t_R _1073_ (.A(_0560_),
    .Y(net371));
 INVx2_ASAP7_75t_R _1074_ (.A(_0561_),
    .Y(net372));
 INVx2_ASAP7_75t_R _1075_ (.A(_0562_),
    .Y(net373));
 INVx1_ASAP7_75t_R _1076_ (.A(_0563_),
    .Y(net375));
 INVx1_ASAP7_75t_R _1077_ (.A(_0564_),
    .Y(net376));
 INVx1_ASAP7_75t_R _1078_ (.A(_0565_),
    .Y(net377));
 INVx1_ASAP7_75t_R _1079_ (.A(_0566_),
    .Y(net378));
 INVx2_ASAP7_75t_R _1080_ (.A(_0567_),
    .Y(net379));
 INVx2_ASAP7_75t_R _1081_ (.A(_0568_),
    .Y(net380));
 INVx1_ASAP7_75t_R _1082_ (.A(_0569_),
    .Y(net381));
 INVx1_ASAP7_75t_R _1083_ (.A(_0570_),
    .Y(net382));
 INVx1_ASAP7_75t_R _1084_ (.A(_0571_),
    .Y(net383));
 INVx2_ASAP7_75t_R _1085_ (.A(_0572_),
    .Y(net384));
 INVx2_ASAP7_75t_R _1086_ (.A(_0573_),
    .Y(net386));
 INVx2_ASAP7_75t_R _1087_ (.A(_0574_),
    .Y(net387));
 INVx2_ASAP7_75t_R _1088_ (.A(_0575_),
    .Y(net388));
 INVx2_ASAP7_75t_R _1089_ (.A(_0576_),
    .Y(net389));
 INVx1_ASAP7_75t_R _1090_ (.A(_0577_),
    .Y(net458));
 INVx1_ASAP7_75t_R _1091_ (.A(_0578_),
    .Y(net469));
 INVx1_ASAP7_75t_R _1092_ (.A(_0579_),
    .Y(net480));
 INVx1_ASAP7_75t_R _1093_ (.A(_0580_),
    .Y(net491));
 INVx1_ASAP7_75t_R _1094_ (.A(_0581_),
    .Y(net502));
 INVx1_ASAP7_75t_R _1095_ (.A(_0582_),
    .Y(net513));
 INVx1_ASAP7_75t_R _1096_ (.A(_0583_),
    .Y(net518));
 INVx1_ASAP7_75t_R _1097_ (.A(_0584_),
    .Y(net519));
 INVx1_ASAP7_75t_R _1098_ (.A(_0585_),
    .Y(net520));
 INVx1_ASAP7_75t_R _1099_ (.A(_0586_),
    .Y(net521));
 INVx1_ASAP7_75t_R _1100_ (.A(_0587_),
    .Y(net459));
 INVx1_ASAP7_75t_R _1101_ (.A(_0588_),
    .Y(net460));
 INVx1_ASAP7_75t_R _1102_ (.A(_0589_),
    .Y(net461));
 INVx1_ASAP7_75t_R _1103_ (.A(_0590_),
    .Y(net462));
 INVx1_ASAP7_75t_R _1104_ (.A(_0591_),
    .Y(net463));
 INVx1_ASAP7_75t_R _1105_ (.A(_0592_),
    .Y(net464));
 INVx1_ASAP7_75t_R _1106_ (.A(_0593_),
    .Y(net465));
 INVx1_ASAP7_75t_R _1107_ (.A(_0594_),
    .Y(net466));
 INVx1_ASAP7_75t_R _1108_ (.A(_0595_),
    .Y(net467));
 INVx1_ASAP7_75t_R _1109_ (.A(_0596_),
    .Y(net468));
 INVx1_ASAP7_75t_R _1110_ (.A(_0597_),
    .Y(net470));
 INVx1_ASAP7_75t_R _1111_ (.A(_0598_),
    .Y(net471));
 INVx1_ASAP7_75t_R _1112_ (.A(_0599_),
    .Y(net472));
 INVx1_ASAP7_75t_R _1113_ (.A(_0600_),
    .Y(net473));
 INVx1_ASAP7_75t_R _1114_ (.A(_0601_),
    .Y(net474));
 INVx1_ASAP7_75t_R _1115_ (.A(_0602_),
    .Y(net475));
 INVx1_ASAP7_75t_R _1116_ (.A(_0603_),
    .Y(net476));
 INVx1_ASAP7_75t_R _1117_ (.A(_0604_),
    .Y(net477));
 INVx1_ASAP7_75t_R _1118_ (.A(_0605_),
    .Y(net478));
 INVx1_ASAP7_75t_R _1119_ (.A(_0606_),
    .Y(net479));
 INVx1_ASAP7_75t_R _1120_ (.A(_0607_),
    .Y(net481));
 INVx1_ASAP7_75t_R _1121_ (.A(_0608_),
    .Y(net482));
 INVx1_ASAP7_75t_R _1122_ (.A(_0609_),
    .Y(net483));
 INVx1_ASAP7_75t_R _1123_ (.A(_0610_),
    .Y(net484));
 INVx1_ASAP7_75t_R _1124_ (.A(_0611_),
    .Y(net485));
 INVx1_ASAP7_75t_R _1125_ (.A(_0612_),
    .Y(net486));
 INVx1_ASAP7_75t_R _1126_ (.A(_0613_),
    .Y(net487));
 INVx1_ASAP7_75t_R _1127_ (.A(_0614_),
    .Y(net488));
 INVx1_ASAP7_75t_R _1128_ (.A(_0615_),
    .Y(net489));
 INVx1_ASAP7_75t_R _1129_ (.A(_0616_),
    .Y(net490));
 INVx1_ASAP7_75t_R _1130_ (.A(_0617_),
    .Y(net492));
 INVx1_ASAP7_75t_R _1131_ (.A(_0618_),
    .Y(net493));
 INVx1_ASAP7_75t_R _1132_ (.A(_0619_),
    .Y(net494));
 INVx1_ASAP7_75t_R _1133_ (.A(_0620_),
    .Y(net495));
 INVx1_ASAP7_75t_R _1134_ (.A(_0621_),
    .Y(net496));
 INVx1_ASAP7_75t_R _1135_ (.A(_0622_),
    .Y(net497));
 INVx1_ASAP7_75t_R _1136_ (.A(_0623_),
    .Y(net498));
 INVx1_ASAP7_75t_R _1137_ (.A(_0624_),
    .Y(net499));
 INVx1_ASAP7_75t_R _1138_ (.A(_0625_),
    .Y(net500));
 INVx1_ASAP7_75t_R _1139_ (.A(_0626_),
    .Y(net501));
 INVx1_ASAP7_75t_R _1140_ (.A(_0627_),
    .Y(net503));
 INVx1_ASAP7_75t_R _1141_ (.A(_0628_),
    .Y(net504));
 INVx1_ASAP7_75t_R _1142_ (.A(_0629_),
    .Y(net505));
 INVx1_ASAP7_75t_R _1143_ (.A(_0630_),
    .Y(net506));
 INVx1_ASAP7_75t_R _1144_ (.A(_0631_),
    .Y(net507));
 INVx1_ASAP7_75t_R _1145_ (.A(_0632_),
    .Y(net508));
 INVx1_ASAP7_75t_R _1146_ (.A(_0633_),
    .Y(net509));
 INVx1_ASAP7_75t_R _1147_ (.A(_0634_),
    .Y(net510));
 INVx1_ASAP7_75t_R _1148_ (.A(_0635_),
    .Y(net511));
 INVx1_ASAP7_75t_R _1149_ (.A(_0636_),
    .Y(net512));
 INVx1_ASAP7_75t_R _1150_ (.A(_0637_),
    .Y(net514));
 INVx1_ASAP7_75t_R _1151_ (.A(_0638_),
    .Y(net515));
 INVx1_ASAP7_75t_R _1152_ (.A(_0639_),
    .Y(net516));
 INVx1_ASAP7_75t_R _1153_ (.A(_0640_),
    .Y(net517));
 INVx1_ASAP7_75t_R _1154_ (.A(_0641_),
    .Y(net394));
 INVx2_ASAP7_75t_R _1155_ (.A(_0642_),
    .Y(net405));
 INVx2_ASAP7_75t_R _1156_ (.A(_0643_),
    .Y(net416));
 INVx2_ASAP7_75t_R _1157_ (.A(_0644_),
    .Y(net427));
 INVx2_ASAP7_75t_R _1158_ (.A(_0645_),
    .Y(net438));
 INVx2_ASAP7_75t_R _1159_ (.A(_0646_),
    .Y(net449));
 INVx1_ASAP7_75t_R _1160_ (.A(_0647_),
    .Y(net454));
 INVx1_ASAP7_75t_R _1161_ (.A(_0648_),
    .Y(net455));
 INVx1_ASAP7_75t_R _1162_ (.A(_0649_),
    .Y(net456));
 INVx1_ASAP7_75t_R _1163_ (.A(_0650_),
    .Y(net457));
 INVx1_ASAP7_75t_R _1164_ (.A(_0651_),
    .Y(net395));
 INVx1_ASAP7_75t_R _1165_ (.A(_0652_),
    .Y(net396));
 INVx1_ASAP7_75t_R _1166_ (.A(_0653_),
    .Y(net397));
 INVx1_ASAP7_75t_R _1167_ (.A(_0654_),
    .Y(net398));
 INVx2_ASAP7_75t_R _1168_ (.A(_0655_),
    .Y(net399));
 INVx2_ASAP7_75t_R _1169_ (.A(_0656_),
    .Y(net400));
 INVx1_ASAP7_75t_R _1170_ (.A(_0657_),
    .Y(net401));
 INVx1_ASAP7_75t_R _1171_ (.A(_0658_),
    .Y(net402));
 INVx1_ASAP7_75t_R _1172_ (.A(_0659_),
    .Y(net403));
 INVx1_ASAP7_75t_R _1173_ (.A(_0660_),
    .Y(net404));
 INVx1_ASAP7_75t_R _1174_ (.A(_0661_),
    .Y(net406));
 INVx1_ASAP7_75t_R _1175_ (.A(_0662_),
    .Y(net407));
 INVx1_ASAP7_75t_R _1176_ (.A(_0663_),
    .Y(net408));
 INVx1_ASAP7_75t_R _1177_ (.A(_0664_),
    .Y(net409));
 INVx1_ASAP7_75t_R _1178_ (.A(_0665_),
    .Y(net410));
 INVx1_ASAP7_75t_R _1179_ (.A(_0666_),
    .Y(net411));
 INVx2_ASAP7_75t_R _1180_ (.A(_0667_),
    .Y(net412));
 INVx1_ASAP7_75t_R _1181_ (.A(_0668_),
    .Y(net413));
 INVx1_ASAP7_75t_R _1182_ (.A(_0669_),
    .Y(net414));
 INVx1_ASAP7_75t_R _1183_ (.A(_0670_),
    .Y(net415));
 INVx1_ASAP7_75t_R _1184_ (.A(_0671_),
    .Y(net417));
 INVx1_ASAP7_75t_R _1185_ (.A(_0672_),
    .Y(net418));
 INVx1_ASAP7_75t_R _1186_ (.A(_0673_),
    .Y(net419));
 INVx1_ASAP7_75t_R _1187_ (.A(_0674_),
    .Y(net420));
 INVx1_ASAP7_75t_R _1188_ (.A(_0675_),
    .Y(net421));
 INVx1_ASAP7_75t_R _1189_ (.A(_0676_),
    .Y(net422));
 INVx1_ASAP7_75t_R _1190_ (.A(_0677_),
    .Y(net423));
 INVx1_ASAP7_75t_R _1191_ (.A(_0678_),
    .Y(net424));
 INVx1_ASAP7_75t_R _1192_ (.A(_0679_),
    .Y(net425));
 INVx1_ASAP7_75t_R _1193_ (.A(_0680_),
    .Y(net426));
 INVx1_ASAP7_75t_R _1194_ (.A(_0681_),
    .Y(net428));
 INVx1_ASAP7_75t_R _1195_ (.A(_0682_),
    .Y(net429));
 INVx1_ASAP7_75t_R _1196_ (.A(_0683_),
    .Y(net430));
 INVx1_ASAP7_75t_R _1197_ (.A(_0684_),
    .Y(net431));
 INVx1_ASAP7_75t_R _1198_ (.A(_0685_),
    .Y(net432));
 INVx1_ASAP7_75t_R _1199_ (.A(_0686_),
    .Y(net433));
 INVx1_ASAP7_75t_R _1200_ (.A(_0687_),
    .Y(net434));
 INVx1_ASAP7_75t_R _1201_ (.A(_0688_),
    .Y(net435));
 INVx1_ASAP7_75t_R _1202_ (.A(_0689_),
    .Y(net436));
 INVx1_ASAP7_75t_R _1203_ (.A(_0690_),
    .Y(net437));
 INVx1_ASAP7_75t_R _1204_ (.A(_0691_),
    .Y(net439));
 INVx1_ASAP7_75t_R _1205_ (.A(_0692_),
    .Y(net440));
 INVx1_ASAP7_75t_R _1206_ (.A(_0693_),
    .Y(net441));
 INVx1_ASAP7_75t_R _1207_ (.A(_0694_),
    .Y(net442));
 INVx1_ASAP7_75t_R _1208_ (.A(_0695_),
    .Y(net443));
 INVx1_ASAP7_75t_R _1209_ (.A(_0696_),
    .Y(net444));
 INVx1_ASAP7_75t_R _1210_ (.A(_0697_),
    .Y(net445));
 INVx1_ASAP7_75t_R _1211_ (.A(_0698_),
    .Y(net446));
 INVx1_ASAP7_75t_R _1212_ (.A(_0699_),
    .Y(net447));
 INVx1_ASAP7_75t_R _1213_ (.A(_0700_),
    .Y(net448));
 INVx1_ASAP7_75t_R _1214_ (.A(_0701_),
    .Y(net450));
 INVx1_ASAP7_75t_R _1215_ (.A(_0702_),
    .Y(net451));
 INVx1_ASAP7_75t_R _1216_ (.A(_0703_),
    .Y(net452));
 INVx1_ASAP7_75t_R _1217_ (.A(_0704_),
    .Y(net453));
 INVx1_ASAP7_75t_R _1218_ (.A(_0705_),
    .Y(net266));
 INVx1_ASAP7_75t_R _1219_ (.A(_0706_),
    .Y(net277));
 INVx1_ASAP7_75t_R _1220_ (.A(_0707_),
    .Y(net288));
 INVx1_ASAP7_75t_R _1221_ (.A(_0708_),
    .Y(net299));
 INVx1_ASAP7_75t_R _1222_ (.A(_0709_),
    .Y(net310));
 INVx1_ASAP7_75t_R _1223_ (.A(_0710_),
    .Y(net321));
 INVx1_ASAP7_75t_R _1224_ (.A(_0711_),
    .Y(net326));
 INVx1_ASAP7_75t_R _1225_ (.A(_0712_),
    .Y(net327));
 INVx1_ASAP7_75t_R _1226_ (.A(_0713_),
    .Y(net328));
 INVx1_ASAP7_75t_R _1227_ (.A(_0714_),
    .Y(net329));
 INVx1_ASAP7_75t_R _1228_ (.A(_0715_),
    .Y(net267));
 INVx1_ASAP7_75t_R _1229_ (.A(_0716_),
    .Y(net268));
 INVx1_ASAP7_75t_R _1230_ (.A(_0717_),
    .Y(net269));
 INVx1_ASAP7_75t_R _1231_ (.A(_0718_),
    .Y(net270));
 INVx1_ASAP7_75t_R _1232_ (.A(_0719_),
    .Y(net271));
 INVx1_ASAP7_75t_R _1233_ (.A(_0720_),
    .Y(net272));
 INVx1_ASAP7_75t_R _1234_ (.A(_0721_),
    .Y(net273));
 INVx1_ASAP7_75t_R _1235_ (.A(_0722_),
    .Y(net274));
 INVx1_ASAP7_75t_R _1236_ (.A(_0723_),
    .Y(net275));
 INVx1_ASAP7_75t_R _1237_ (.A(_0724_),
    .Y(net276));
 INVx1_ASAP7_75t_R _1238_ (.A(_0725_),
    .Y(net278));
 INVx1_ASAP7_75t_R _1239_ (.A(_0726_),
    .Y(net279));
 INVx1_ASAP7_75t_R _1240_ (.A(_0727_),
    .Y(net280));
 INVx1_ASAP7_75t_R _1241_ (.A(_0728_),
    .Y(net281));
 INVx1_ASAP7_75t_R _1242_ (.A(_0729_),
    .Y(net282));
 INVx1_ASAP7_75t_R _1243_ (.A(_0730_),
    .Y(net283));
 INVx1_ASAP7_75t_R _1244_ (.A(_0731_),
    .Y(net284));
 INVx1_ASAP7_75t_R _1245_ (.A(_0732_),
    .Y(net285));
 INVx1_ASAP7_75t_R _1246_ (.A(_0733_),
    .Y(net286));
 INVx1_ASAP7_75t_R _1247_ (.A(_0734_),
    .Y(net287));
 INVx1_ASAP7_75t_R _1248_ (.A(_0735_),
    .Y(net289));
 INVx1_ASAP7_75t_R _1249_ (.A(_0736_),
    .Y(net290));
 INVx1_ASAP7_75t_R _1250_ (.A(_0737_),
    .Y(net291));
 INVx1_ASAP7_75t_R _1251_ (.A(_0738_),
    .Y(net292));
 INVx1_ASAP7_75t_R _1252_ (.A(_0739_),
    .Y(net293));
 INVx1_ASAP7_75t_R _1253_ (.A(_0740_),
    .Y(net294));
 INVx1_ASAP7_75t_R _1254_ (.A(_0741_),
    .Y(net295));
 INVx1_ASAP7_75t_R _1255_ (.A(_0742_),
    .Y(net296));
 INVx1_ASAP7_75t_R _1256_ (.A(_0743_),
    .Y(net297));
 INVx1_ASAP7_75t_R _1257_ (.A(_0744_),
    .Y(net298));
 INVx1_ASAP7_75t_R _1258_ (.A(_0745_),
    .Y(net300));
 INVx1_ASAP7_75t_R _1259_ (.A(_0746_),
    .Y(net301));
 INVx1_ASAP7_75t_R _1260_ (.A(_0747_),
    .Y(net302));
 INVx1_ASAP7_75t_R _1261_ (.A(_0748_),
    .Y(net303));
 INVx1_ASAP7_75t_R _1262_ (.A(_0749_),
    .Y(net304));
 INVx1_ASAP7_75t_R _1263_ (.A(_0750_),
    .Y(net305));
 INVx1_ASAP7_75t_R _1264_ (.A(_0751_),
    .Y(net306));
 INVx1_ASAP7_75t_R _1265_ (.A(_0752_),
    .Y(net307));
 INVx1_ASAP7_75t_R _1266_ (.A(_0753_),
    .Y(net308));
 INVx1_ASAP7_75t_R _1267_ (.A(_0754_),
    .Y(net309));
 INVx1_ASAP7_75t_R _1268_ (.A(_0755_),
    .Y(net311));
 INVx1_ASAP7_75t_R _1269_ (.A(_0756_),
    .Y(net312));
 INVx1_ASAP7_75t_R _1270_ (.A(_0757_),
    .Y(net313));
 INVx1_ASAP7_75t_R _1271_ (.A(_0758_),
    .Y(net314));
 INVx1_ASAP7_75t_R _1272_ (.A(_0759_),
    .Y(net315));
 INVx1_ASAP7_75t_R _1273_ (.A(_0760_),
    .Y(net316));
 INVx1_ASAP7_75t_R _1274_ (.A(_0761_),
    .Y(net317));
 INVx1_ASAP7_75t_R _1275_ (.A(_0762_),
    .Y(net318));
 INVx1_ASAP7_75t_R _1276_ (.A(_0763_),
    .Y(net319));
 INVx1_ASAP7_75t_R _1277_ (.A(_0764_),
    .Y(net320));
 INVx1_ASAP7_75t_R _1278_ (.A(_0765_),
    .Y(net322));
 INVx1_ASAP7_75t_R _1279_ (.A(_0766_),
    .Y(net323));
 INVx1_ASAP7_75t_R _1280_ (.A(_0767_),
    .Y(net324));
 INVx1_ASAP7_75t_R _1281_ (.A(_0768_),
    .Y(net325));
 BUFx2_ASAP7_75t_R _1282_ (.A(io_lsbIns_1),
    .Y(net258));
 BUFx3_ASAP7_75t_R _1283_ (.A(io_lsbIns_2),
    .Y(net259));
 BUFx2_ASAP7_75t_R _1284_ (.A(io_lsbIns_3),
    .Y(net260));
 BUFx2_ASAP7_75t_R _1285_ (.A(io_lsbIns_5),
    .Y(net262));
 BUFx3_ASAP7_75t_R _1286_ (.A(io_lsbIns_6),
    .Y(net263));
 BUFx2_ASAP7_75t_R _1287_ (.A(io_lsbIns_7),
    .Y(net264));
 BUFx2_ASAP7_75t_R _1288_ (.A(net265),
    .Y(net330));
 DFFHQNx3_ASAP7_75t_R \io_lsbOuts_3$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(net257),
    .QN(_0256_));
 DFFHQNx2_ASAP7_75t_R \io_lsbOuts_7$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0064_),
    .QN(_0513_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[0]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(_0000_),
    .QN(_0705_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[10]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0001_),
    .QN(_0715_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[11]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0002_),
    .QN(_0716_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[12]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0003_),
    .QN(_0717_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[13]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0004_),
    .QN(_0718_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[14]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0005_),
    .QN(_0719_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[15]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0006_),
    .QN(_0720_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[16]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0007_),
    .QN(_0721_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[17]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0008_),
    .QN(_0722_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[18]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0009_),
    .QN(_0723_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[19]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0010_),
    .QN(_0724_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[1]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(_0011_),
    .QN(_0706_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[20]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0012_),
    .QN(_0725_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[21]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0013_),
    .QN(_0726_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[22]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0014_),
    .QN(_0727_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[23]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0015_),
    .QN(_0728_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[24]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0016_),
    .QN(_0729_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[25]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0017_),
    .QN(_0730_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[26]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0018_),
    .QN(_0731_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[27]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0019_),
    .QN(_0732_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[28]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0020_),
    .QN(_0733_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[29]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0021_),
    .QN(_0734_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[2]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(_0022_),
    .QN(_0707_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[30]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0023_),
    .QN(_0735_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[31]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0024_),
    .QN(_0736_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[32]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0025_),
    .QN(_0737_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[33]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0026_),
    .QN(_0738_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[34]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0027_),
    .QN(_0739_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[35]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0028_),
    .QN(_0740_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[36]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0029_),
    .QN(_0741_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[37]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0030_),
    .QN(_0742_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[38]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0031_),
    .QN(_0743_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[39]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0032_),
    .QN(_0744_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[3]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0033_),
    .QN(_0708_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[40]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0034_),
    .QN(_0745_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[41]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0035_),
    .QN(_0746_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[42]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0036_),
    .QN(_0747_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[43]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(_0037_),
    .QN(_0748_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[44]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0038_),
    .QN(_0749_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[45]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0039_),
    .QN(_0750_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[46]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0040_),
    .QN(_0751_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[47]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0041_),
    .QN(_0752_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[48]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(_0042_),
    .QN(_0753_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[49]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0043_),
    .QN(_0754_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[4]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0044_),
    .QN(_0709_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[50]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(_0045_),
    .QN(_0755_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[51]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(_0046_),
    .QN(_0756_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[52]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(_0047_),
    .QN(_0757_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[53]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0048_),
    .QN(_0758_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[54]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(_0049_),
    .QN(_0759_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[55]$_DFF_P_  (.CLK(clknet_leaf_15_clock),
    .D(_0050_),
    .QN(_0760_));
 DFFHQNx3_ASAP7_75t_R \io_outs_down[56]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0051_),
    .QN(_0761_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[57]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0052_),
    .QN(_0762_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[58]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0053_),
    .QN(_0763_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[59]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0054_),
    .QN(_0764_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[5]$_DFF_P_  (.CLK(clknet_leaf_20_clock),
    .D(_0055_),
    .QN(_0710_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[60]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0056_),
    .QN(_0765_));
 DFFHQNx1_ASAP7_75t_R \io_outs_down[61]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0057_),
    .QN(_0766_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[62]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0058_),
    .QN(_0767_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[63]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0059_),
    .QN(_0768_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[6]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0060_),
    .QN(_0711_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[7]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0061_),
    .QN(_0712_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[8]$_DFF_P_  (.CLK(clknet_leaf_16_clock),
    .D(_0062_),
    .QN(_0713_));
 DFFHQNx2_ASAP7_75t_R \io_outs_down[9]$_DFF_P_  (.CLK(clknet_leaf_19_clock),
    .D(_0063_),
    .QN(_0714_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[10]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(_0065_),
    .QN(_0523_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[11]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0066_),
    .QN(_0524_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[12]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0067_),
    .QN(_0525_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[13]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0068_),
    .QN(_0526_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[14]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0069_),
    .QN(_0527_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[15]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0070_),
    .QN(_0528_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[16]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0071_),
    .QN(_0529_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[17]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0072_),
    .QN(_0530_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[18]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0073_),
    .QN(_0531_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[19]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0074_),
    .QN(_0532_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[1]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0075_),
    .QN(_0514_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[20]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0076_),
    .QN(_0533_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[21]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0077_),
    .QN(_0534_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[22]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0078_),
    .QN(_0535_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[23]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0079_),
    .QN(_0536_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[24]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0080_),
    .QN(_0537_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[25]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(_0081_),
    .QN(_0538_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[26]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0082_),
    .QN(_0539_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[27]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(_0083_),
    .QN(_0540_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[28]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0084_),
    .QN(_0541_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[29]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(_0085_),
    .QN(_0542_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[2]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(_0086_),
    .QN(_0515_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[30]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0087_),
    .QN(_0543_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[31]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0088_),
    .QN(_0544_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[32]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0089_),
    .QN(_0545_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[33]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(_0090_),
    .QN(_0546_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[34]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0091_),
    .QN(_0547_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[35]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0092_),
    .QN(_0548_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[36]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0093_),
    .QN(_0549_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[37]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0094_),
    .QN(_0550_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[38]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0095_),
    .QN(_0551_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[39]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0096_),
    .QN(_0552_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[3]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0097_),
    .QN(_0516_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[40]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(_0098_),
    .QN(_0553_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[41]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0099_),
    .QN(_0554_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[42]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0100_),
    .QN(_0555_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[43]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0101_),
    .QN(_0556_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[44]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0102_),
    .QN(_0557_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[45]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0103_),
    .QN(_0558_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[46]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0104_),
    .QN(_0559_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[47]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0105_),
    .QN(_0560_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[48]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0106_),
    .QN(_0561_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[49]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(_0107_),
    .QN(_0562_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[4]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0108_),
    .QN(_0517_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[50]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0109_),
    .QN(_0563_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[51]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0110_),
    .QN(_0564_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[52]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0111_),
    .QN(_0565_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[53]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0112_),
    .QN(_0566_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[54]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0113_),
    .QN(_0567_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[55]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0114_),
    .QN(_0568_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[56]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0115_),
    .QN(_0569_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[57]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0116_),
    .QN(_0570_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[58]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0117_),
    .QN(_0571_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[59]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0118_),
    .QN(_0572_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[5]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0119_),
    .QN(_0518_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[60]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(_0120_),
    .QN(_0573_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[61]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0121_),
    .QN(_0574_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[62]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(_0122_),
    .QN(_0575_));
 DFFHQNx2_ASAP7_75t_R \io_outs_left[63]$_DFF_P_  (.CLK(clknet_leaf_11_clock),
    .D(_0123_),
    .QN(_0576_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[6]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0124_),
    .QN(_0519_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[7]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(_0125_),
    .QN(_0520_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[8]$_DFF_P_  (.CLK(clknet_leaf_4_clock),
    .D(_0126_),
    .QN(_0521_));
 DFFHQNx3_ASAP7_75t_R \io_outs_left[9]$_DFF_P_  (.CLK(clknet_leaf_3_clock),
    .D(_0127_),
    .QN(_0522_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[0]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0128_),
    .QN(_0641_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[10]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0129_),
    .QN(_0651_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[11]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0130_),
    .QN(_0652_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[12]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0131_),
    .QN(_0653_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[13]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0132_),
    .QN(_0654_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[14]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0133_),
    .QN(_0655_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[15]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(_0134_),
    .QN(_0656_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[16]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0135_),
    .QN(_0657_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[17]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0136_),
    .QN(_0658_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[18]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0137_),
    .QN(_0659_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[19]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0138_),
    .QN(_0660_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[1]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0139_),
    .QN(_0642_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[20]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0140_),
    .QN(_0661_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[21]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0141_),
    .QN(_0662_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[22]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0142_),
    .QN(_0663_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[23]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0143_),
    .QN(_0664_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[24]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0144_),
    .QN(_0665_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[25]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0145_),
    .QN(_0666_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[26]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0146_),
    .QN(_0667_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[27]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0147_),
    .QN(_0668_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[28]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0148_),
    .QN(_0669_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[29]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0149_),
    .QN(_0670_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[2]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0150_),
    .QN(_0643_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[30]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0151_),
    .QN(_0671_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[31]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0152_),
    .QN(_0672_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[32]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0153_),
    .QN(_0673_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[33]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0154_),
    .QN(_0674_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[34]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0155_),
    .QN(_0675_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[35]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0156_),
    .QN(_0676_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[36]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0157_),
    .QN(_0677_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[37]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0158_),
    .QN(_0678_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[38]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0159_),
    .QN(_0679_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[39]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0160_),
    .QN(_0680_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[3]$_DFF_P_  (.CLK(clknet_leaf_1_clock),
    .D(_0161_),
    .QN(_0644_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[40]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0162_),
    .QN(_0681_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[41]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0163_),
    .QN(_0682_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[42]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0164_),
    .QN(_0683_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[43]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0165_),
    .QN(_0684_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[44]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0166_),
    .QN(_0685_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[45]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0167_),
    .QN(_0686_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[46]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0168_),
    .QN(_0687_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[47]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0169_),
    .QN(_0688_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[48]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0170_),
    .QN(_0689_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[49]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0171_),
    .QN(_0690_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[4]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0172_),
    .QN(_0645_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[50]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0173_),
    .QN(_0691_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[51]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0174_),
    .QN(_0692_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[52]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0175_),
    .QN(_0693_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[53]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0176_),
    .QN(_0694_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[54]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0177_),
    .QN(_0695_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[55]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0178_),
    .QN(_0696_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[56]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0179_),
    .QN(_0697_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[57]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0180_),
    .QN(_0698_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[58]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0181_),
    .QN(_0699_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[59]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0182_),
    .QN(_0700_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[5]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0183_),
    .QN(_0646_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[60]$_DFF_P_  (.CLK(clknet_leaf_14_clock),
    .D(_0184_),
    .QN(_0701_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[61]$_DFF_P_  (.CLK(clknet_leaf_12_clock),
    .D(_0185_),
    .QN(_0702_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[62]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0186_),
    .QN(_0703_));
 DFFHQNx2_ASAP7_75t_R \io_outs_right[63]$_DFF_P_  (.CLK(clknet_leaf_10_clock),
    .D(_0187_),
    .QN(_0704_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[6]$_DFF_P_  (.CLK(clknet_leaf_18_clock),
    .D(_0188_),
    .QN(_0647_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[7]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0189_),
    .QN(_0648_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[8]$_DFF_P_  (.CLK(clknet_leaf_17_clock),
    .D(_0190_),
    .QN(_0649_));
 DFFHQNx3_ASAP7_75t_R \io_outs_right[9]$_DFF_P_  (.CLK(clknet_leaf_13_clock),
    .D(_0191_),
    .QN(_0650_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[0]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(_0192_),
    .QN(_0577_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[10]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(_0193_),
    .QN(_0587_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[11]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0194_),
    .QN(_0588_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[12]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0195_),
    .QN(_0589_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[13]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(_0196_),
    .QN(_0590_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[14]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(_0197_),
    .QN(_0591_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[15]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(_0198_),
    .QN(_0592_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[16]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0199_),
    .QN(_0593_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[17]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(_0200_),
    .QN(_0594_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[18]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0201_),
    .QN(_0595_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[19]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(_0202_),
    .QN(_0596_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[1]$_DFF_P_  (.CLK(clknet_leaf_2_clock),
    .D(_0203_),
    .QN(_0578_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[20]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0204_),
    .QN(_0597_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[21]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0205_),
    .QN(_0598_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[22]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0206_),
    .QN(_0599_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[23]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(_0207_),
    .QN(_0600_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[24]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0208_),
    .QN(_0601_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[25]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0209_),
    .QN(_0602_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[26]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0210_),
    .QN(_0603_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[27]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0211_),
    .QN(_0604_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[28]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0212_),
    .QN(_0605_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[29]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0213_),
    .QN(_0606_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[2]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(_0214_),
    .QN(_0579_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[30]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0215_),
    .QN(_0607_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[31]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0216_),
    .QN(_0608_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[32]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0217_),
    .QN(_0609_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[33]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0218_),
    .QN(_0610_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[34]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(_0219_),
    .QN(_0611_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[35]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0220_),
    .QN(_0612_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[36]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0221_),
    .QN(_0613_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[37]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0222_),
    .QN(_0614_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[38]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0223_),
    .QN(_0615_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[39]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0224_),
    .QN(_0616_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[3]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(_0225_),
    .QN(_0580_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[40]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0226_),
    .QN(_0617_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[41]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0227_),
    .QN(_0618_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[42]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0228_),
    .QN(_0619_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[43]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0229_),
    .QN(_0620_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[44]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0230_),
    .QN(_0621_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[45]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0231_),
    .QN(_0622_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[46]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0232_),
    .QN(_0623_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[47]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0233_),
    .QN(_0624_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[48]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0234_),
    .QN(_0625_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[49]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0235_),
    .QN(_0626_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[4]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(_0236_),
    .QN(_0581_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[50]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0237_),
    .QN(_0627_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[51]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0238_),
    .QN(_0628_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[52]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0239_),
    .QN(_0629_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[53]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0240_),
    .QN(_0630_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[54]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0241_),
    .QN(_0631_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[55]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0242_),
    .QN(_0632_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[56]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0243_),
    .QN(_0633_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[57]$_DFF_P_  (.CLK(clknet_leaf_8_clock),
    .D(_0244_),
    .QN(_0634_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[58]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0245_),
    .QN(_0635_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[59]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0246_),
    .QN(_0636_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[5]$_DFF_P_  (.CLK(clknet_leaf_6_clock),
    .D(_0247_),
    .QN(_0582_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[60]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0248_),
    .QN(_0637_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[61]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0249_),
    .QN(_0638_));
 DFFHQNx2_ASAP7_75t_R \io_outs_up[62]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0250_),
    .QN(_0639_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[63]$_DFF_P_  (.CLK(clknet_leaf_9_clock),
    .D(_0251_),
    .QN(_0640_));
 DFFHQNx1_ASAP7_75t_R \io_outs_up[6]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0252_),
    .QN(_0583_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[7]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0253_),
    .QN(_0584_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[8]$_DFF_P_  (.CLK(clknet_leaf_5_clock),
    .D(_0254_),
    .QN(_0585_));
 DFFHQNx3_ASAP7_75t_R \io_outs_up[9]$_DFF_P_  (.CLK(clknet_leaf_7_clock),
    .D(_0255_),
    .QN(_0586_));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_152 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_153 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_154 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_155 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_156 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_157 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_158 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_159 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_160 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_161 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_162 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_163 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_164 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_165 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_166 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_167 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_168 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_169 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_170 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_171 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_172 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_173 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_174 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_175 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_176 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_177 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_178 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_179 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_180 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_29_Left_181 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_30_Left_182 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_31_Left_183 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_32_Left_184 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_33_Left_185 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_34_Left_186 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_35_Left_187 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_36_Left_188 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_37_Left_189 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_38_Left_190 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_39_Left_191 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_40_Left_192 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_41_Left_193 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_42_Left_194 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_43_Left_195 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_44_Left_196 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_45_Left_197 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_46_Left_198 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_47_Left_199 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_48_Left_200 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_49_Left_201 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_50_Left_202 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_51_Left_203 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_52_Left_204 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_53_Left_205 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_54_Left_206 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_55_Left_207 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_56_Left_208 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_57_Left_209 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_58_Left_210 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_59_Left_211 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_60_Left_212 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_61_Left_213 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_62_Left_214 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_63_Left_215 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_64_Left_216 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_65_Left_217 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_66_Left_218 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_67_Left_219 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_68_Left_220 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_69_Left_221 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_70_Left_222 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_71_Left_223 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_72_Left_224 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_73_Left_225 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_74_Left_226 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_75_Left_227 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_76_Left_228 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_77_Left_229 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_78_Left_230 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_79_Left_231 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_80_Left_232 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_81_Left_233 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_82_Left_234 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_83_Left_235 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_84_Left_236 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_85_Left_237 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_86_Left_238 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_87_Left_239 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_88_Left_240 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_89_Left_241 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_90_Left_242 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_91_Left_243 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_92_Left_244 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_93_Left_245 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_94_Left_246 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_95_Left_247 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_96_Left_248 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_97_Left_249 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_98_Left_250 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_99_Left_251 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_100_Left_252 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_101_Left_253 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_102_Left_254 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_103_Left_255 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_104_Left_256 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_105_Left_257 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_106_Left_258 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_107_Left_259 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_108_Left_260 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_109_Left_261 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_110_Left_262 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_111_Left_263 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_112_Left_264 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_113_Left_265 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_114_Left_266 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_115_Left_267 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_116_Left_268 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_117_Left_269 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_118_Left_270 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_119_Left_271 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_120_Left_272 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_121_Left_273 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_122_Left_274 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_123_Left_275 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_124_Left_276 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_125_Left_277 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_126_Left_278 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_127_Left_279 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_128_Left_280 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_129_Left_281 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_130_Left_282 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_131_Left_283 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_132_Left_284 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_133_Left_285 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_134_Left_286 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_135_Left_287 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_136_Left_288 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_137_Left_289 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_138_Left_290 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_139_Left_291 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_140_Left_292 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_141_Left_293 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_142_Left_294 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_143_Left_295 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_144_Left_296 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_145_Left_297 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_146_Left_298 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_147_Left_299 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_148_Left_300 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_149_Left_301 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_150_Left_302 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_151_Left_303 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_0_304 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_2_305 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_4_306 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_6_307 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_8_308 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_10_309 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_12_310 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_14_311 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_16_312 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_18_313 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_20_314 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_22_315 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_24_316 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_26_317 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_28_318 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_30_319 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_32_320 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_34_321 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_36_322 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_38_323 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_40_324 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_42_325 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_44_326 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_46_327 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_48_328 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_50_329 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_52_330 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_54_331 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_56_332 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_58_333 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_60_334 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_62_335 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_64_336 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_66_337 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_68_338 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_70_339 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_72_340 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_74_341 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_76_342 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_78_343 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_80_344 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_82_345 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_84_346 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_86_347 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_88_348 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_90_349 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_92_350 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_94_351 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_96_352 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_98_353 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_100_354 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_102_355 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_104_356 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_106_357 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_108_358 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_110_359 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_112_360 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_114_361 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_116_362 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_118_363 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_120_364 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_122_365 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_124_366 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_126_367 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_128_368 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_130_369 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_132_370 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_134_371 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_136_372 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_138_373 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_140_374 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_142_375 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_144_376 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_146_377 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_148_378 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_150_379 ();
 TAPCELL_ASAP7_75t_R TAP_TAPCELL_ROW_151_380 ();
 BUFx2_ASAP7_75t_R input1 (.A(io_ins_down[0]),
    .Y(net1));
 BUFx2_ASAP7_75t_R input2 (.A(io_ins_down[10]),
    .Y(net2));
 BUFx2_ASAP7_75t_R input3 (.A(io_ins_down[11]),
    .Y(net3));
 BUFx2_ASAP7_75t_R input4 (.A(io_ins_down[12]),
    .Y(net4));
 BUFx2_ASAP7_75t_R input5 (.A(io_ins_down[13]),
    .Y(net5));
 BUFx2_ASAP7_75t_R input6 (.A(io_ins_down[14]),
    .Y(net6));
 BUFx2_ASAP7_75t_R input7 (.A(io_ins_down[15]),
    .Y(net7));
 BUFx2_ASAP7_75t_R input8 (.A(io_ins_down[16]),
    .Y(net8));
 BUFx2_ASAP7_75t_R input9 (.A(io_ins_down[17]),
    .Y(net9));
 BUFx2_ASAP7_75t_R input10 (.A(io_ins_down[18]),
    .Y(net10));
 BUFx2_ASAP7_75t_R input11 (.A(io_ins_down[19]),
    .Y(net11));
 BUFx2_ASAP7_75t_R input12 (.A(io_ins_down[1]),
    .Y(net12));
 BUFx2_ASAP7_75t_R input13 (.A(io_ins_down[20]),
    .Y(net13));
 BUFx2_ASAP7_75t_R input14 (.A(io_ins_down[21]),
    .Y(net14));
 BUFx2_ASAP7_75t_R input15 (.A(io_ins_down[22]),
    .Y(net15));
 BUFx2_ASAP7_75t_R input16 (.A(io_ins_down[23]),
    .Y(net16));
 BUFx2_ASAP7_75t_R input17 (.A(io_ins_down[24]),
    .Y(net17));
 BUFx2_ASAP7_75t_R input18 (.A(io_ins_down[25]),
    .Y(net18));
 BUFx2_ASAP7_75t_R input19 (.A(io_ins_down[26]),
    .Y(net19));
 BUFx2_ASAP7_75t_R input20 (.A(io_ins_down[27]),
    .Y(net20));
 BUFx2_ASAP7_75t_R input21 (.A(io_ins_down[28]),
    .Y(net21));
 BUFx2_ASAP7_75t_R input22 (.A(io_ins_down[29]),
    .Y(net22));
 BUFx2_ASAP7_75t_R input23 (.A(io_ins_down[2]),
    .Y(net23));
 BUFx2_ASAP7_75t_R input24 (.A(io_ins_down[30]),
    .Y(net24));
 BUFx2_ASAP7_75t_R input25 (.A(io_ins_down[31]),
    .Y(net25));
 BUFx2_ASAP7_75t_R input26 (.A(io_ins_down[32]),
    .Y(net26));
 BUFx2_ASAP7_75t_R input27 (.A(io_ins_down[33]),
    .Y(net27));
 BUFx2_ASAP7_75t_R input28 (.A(io_ins_down[34]),
    .Y(net28));
 BUFx2_ASAP7_75t_R input29 (.A(io_ins_down[35]),
    .Y(net29));
 BUFx2_ASAP7_75t_R input30 (.A(io_ins_down[36]),
    .Y(net30));
 BUFx2_ASAP7_75t_R input31 (.A(io_ins_down[37]),
    .Y(net31));
 BUFx2_ASAP7_75t_R input32 (.A(io_ins_down[38]),
    .Y(net32));
 BUFx2_ASAP7_75t_R input33 (.A(io_ins_down[39]),
    .Y(net33));
 BUFx2_ASAP7_75t_R input34 (.A(io_ins_down[3]),
    .Y(net34));
 BUFx2_ASAP7_75t_R input35 (.A(io_ins_down[40]),
    .Y(net35));
 BUFx2_ASAP7_75t_R input36 (.A(io_ins_down[41]),
    .Y(net36));
 BUFx2_ASAP7_75t_R input37 (.A(io_ins_down[42]),
    .Y(net37));
 BUFx2_ASAP7_75t_R input38 (.A(io_ins_down[43]),
    .Y(net38));
 BUFx2_ASAP7_75t_R input39 (.A(io_ins_down[44]),
    .Y(net39));
 BUFx2_ASAP7_75t_R input40 (.A(io_ins_down[45]),
    .Y(net40));
 BUFx2_ASAP7_75t_R input41 (.A(io_ins_down[46]),
    .Y(net41));
 BUFx2_ASAP7_75t_R input42 (.A(io_ins_down[47]),
    .Y(net42));
 BUFx2_ASAP7_75t_R input43 (.A(io_ins_down[48]),
    .Y(net43));
 BUFx2_ASAP7_75t_R input44 (.A(io_ins_down[49]),
    .Y(net44));
 BUFx2_ASAP7_75t_R input45 (.A(io_ins_down[4]),
    .Y(net45));
 BUFx2_ASAP7_75t_R input46 (.A(io_ins_down[50]),
    .Y(net46));
 BUFx2_ASAP7_75t_R input47 (.A(io_ins_down[51]),
    .Y(net47));
 BUFx2_ASAP7_75t_R input48 (.A(io_ins_down[52]),
    .Y(net48));
 BUFx2_ASAP7_75t_R input49 (.A(io_ins_down[53]),
    .Y(net49));
 BUFx2_ASAP7_75t_R input50 (.A(io_ins_down[54]),
    .Y(net50));
 BUFx2_ASAP7_75t_R input51 (.A(io_ins_down[55]),
    .Y(net51));
 BUFx2_ASAP7_75t_R input52 (.A(io_ins_down[56]),
    .Y(net52));
 BUFx2_ASAP7_75t_R input53 (.A(io_ins_down[57]),
    .Y(net53));
 BUFx2_ASAP7_75t_R input54 (.A(io_ins_down[58]),
    .Y(net54));
 BUFx2_ASAP7_75t_R input55 (.A(io_ins_down[59]),
    .Y(net55));
 BUFx2_ASAP7_75t_R input56 (.A(io_ins_down[5]),
    .Y(net56));
 BUFx2_ASAP7_75t_R input57 (.A(io_ins_down[60]),
    .Y(net57));
 BUFx2_ASAP7_75t_R input58 (.A(io_ins_down[61]),
    .Y(net58));
 BUFx2_ASAP7_75t_R input59 (.A(io_ins_down[62]),
    .Y(net59));
 BUFx2_ASAP7_75t_R input60 (.A(io_ins_down[63]),
    .Y(net60));
 BUFx2_ASAP7_75t_R input61 (.A(io_ins_down[6]),
    .Y(net61));
 BUFx2_ASAP7_75t_R input62 (.A(io_ins_down[7]),
    .Y(net62));
 BUFx2_ASAP7_75t_R input63 (.A(io_ins_down[8]),
    .Y(net63));
 BUFx2_ASAP7_75t_R input64 (.A(io_ins_down[9]),
    .Y(net64));
 BUFx2_ASAP7_75t_R input65 (.A(io_ins_left[0]),
    .Y(net65));
 BUFx2_ASAP7_75t_R input66 (.A(io_ins_left[10]),
    .Y(net66));
 BUFx2_ASAP7_75t_R input67 (.A(io_ins_left[11]),
    .Y(net67));
 BUFx2_ASAP7_75t_R input68 (.A(io_ins_left[12]),
    .Y(net68));
 BUFx2_ASAP7_75t_R input69 (.A(io_ins_left[13]),
    .Y(net69));
 BUFx2_ASAP7_75t_R input70 (.A(io_ins_left[14]),
    .Y(net70));
 BUFx2_ASAP7_75t_R input71 (.A(io_ins_left[15]),
    .Y(net71));
 BUFx2_ASAP7_75t_R input72 (.A(io_ins_left[16]),
    .Y(net72));
 BUFx2_ASAP7_75t_R input73 (.A(io_ins_left[17]),
    .Y(net73));
 BUFx2_ASAP7_75t_R input74 (.A(io_ins_left[18]),
    .Y(net74));
 BUFx2_ASAP7_75t_R input75 (.A(io_ins_left[19]),
    .Y(net75));
 BUFx2_ASAP7_75t_R input76 (.A(io_ins_left[1]),
    .Y(net76));
 BUFx2_ASAP7_75t_R input77 (.A(io_ins_left[20]),
    .Y(net77));
 BUFx2_ASAP7_75t_R input78 (.A(io_ins_left[21]),
    .Y(net78));
 BUFx2_ASAP7_75t_R input79 (.A(io_ins_left[22]),
    .Y(net79));
 BUFx2_ASAP7_75t_R input80 (.A(io_ins_left[23]),
    .Y(net80));
 BUFx2_ASAP7_75t_R input81 (.A(io_ins_left[24]),
    .Y(net81));
 BUFx2_ASAP7_75t_R input82 (.A(io_ins_left[25]),
    .Y(net82));
 BUFx2_ASAP7_75t_R input83 (.A(io_ins_left[26]),
    .Y(net83));
 BUFx2_ASAP7_75t_R input84 (.A(io_ins_left[27]),
    .Y(net84));
 BUFx2_ASAP7_75t_R input85 (.A(io_ins_left[28]),
    .Y(net85));
 BUFx2_ASAP7_75t_R input86 (.A(io_ins_left[29]),
    .Y(net86));
 BUFx2_ASAP7_75t_R input87 (.A(io_ins_left[2]),
    .Y(net87));
 BUFx2_ASAP7_75t_R input88 (.A(io_ins_left[30]),
    .Y(net88));
 BUFx2_ASAP7_75t_R input89 (.A(io_ins_left[31]),
    .Y(net89));
 BUFx2_ASAP7_75t_R input90 (.A(io_ins_left[32]),
    .Y(net90));
 BUFx2_ASAP7_75t_R input91 (.A(io_ins_left[33]),
    .Y(net91));
 BUFx2_ASAP7_75t_R input92 (.A(io_ins_left[34]),
    .Y(net92));
 BUFx2_ASAP7_75t_R input93 (.A(io_ins_left[35]),
    .Y(net93));
 BUFx2_ASAP7_75t_R input94 (.A(io_ins_left[36]),
    .Y(net94));
 BUFx2_ASAP7_75t_R input95 (.A(io_ins_left[37]),
    .Y(net95));
 BUFx2_ASAP7_75t_R input96 (.A(io_ins_left[38]),
    .Y(net96));
 BUFx2_ASAP7_75t_R input97 (.A(io_ins_left[39]),
    .Y(net97));
 BUFx2_ASAP7_75t_R input98 (.A(io_ins_left[3]),
    .Y(net98));
 BUFx2_ASAP7_75t_R input99 (.A(io_ins_left[40]),
    .Y(net99));
 BUFx2_ASAP7_75t_R input100 (.A(io_ins_left[41]),
    .Y(net100));
 BUFx2_ASAP7_75t_R input101 (.A(io_ins_left[42]),
    .Y(net101));
 BUFx2_ASAP7_75t_R input102 (.A(io_ins_left[43]),
    .Y(net102));
 BUFx2_ASAP7_75t_R input103 (.A(io_ins_left[44]),
    .Y(net103));
 BUFx2_ASAP7_75t_R input104 (.A(io_ins_left[45]),
    .Y(net104));
 BUFx2_ASAP7_75t_R input105 (.A(io_ins_left[46]),
    .Y(net105));
 BUFx2_ASAP7_75t_R input106 (.A(io_ins_left[47]),
    .Y(net106));
 BUFx2_ASAP7_75t_R input107 (.A(io_ins_left[48]),
    .Y(net107));
 BUFx2_ASAP7_75t_R input108 (.A(io_ins_left[49]),
    .Y(net108));
 BUFx2_ASAP7_75t_R input109 (.A(io_ins_left[4]),
    .Y(net109));
 BUFx2_ASAP7_75t_R input110 (.A(io_ins_left[50]),
    .Y(net110));
 BUFx2_ASAP7_75t_R input111 (.A(io_ins_left[51]),
    .Y(net111));
 BUFx2_ASAP7_75t_R input112 (.A(io_ins_left[52]),
    .Y(net112));
 BUFx2_ASAP7_75t_R input113 (.A(io_ins_left[53]),
    .Y(net113));
 BUFx2_ASAP7_75t_R input114 (.A(io_ins_left[54]),
    .Y(net114));
 BUFx2_ASAP7_75t_R input115 (.A(io_ins_left[55]),
    .Y(net115));
 BUFx2_ASAP7_75t_R input116 (.A(io_ins_left[56]),
    .Y(net116));
 BUFx2_ASAP7_75t_R input117 (.A(io_ins_left[57]),
    .Y(net117));
 BUFx2_ASAP7_75t_R input118 (.A(io_ins_left[58]),
    .Y(net118));
 BUFx2_ASAP7_75t_R input119 (.A(io_ins_left[59]),
    .Y(net119));
 BUFx2_ASAP7_75t_R input120 (.A(io_ins_left[5]),
    .Y(net120));
 BUFx2_ASAP7_75t_R input121 (.A(io_ins_left[60]),
    .Y(net121));
 BUFx2_ASAP7_75t_R input122 (.A(io_ins_left[61]),
    .Y(net122));
 BUFx2_ASAP7_75t_R input123 (.A(io_ins_left[62]),
    .Y(net123));
 BUFx2_ASAP7_75t_R input124 (.A(io_ins_left[63]),
    .Y(net124));
 BUFx2_ASAP7_75t_R input125 (.A(io_ins_left[6]),
    .Y(net125));
 BUFx2_ASAP7_75t_R input126 (.A(io_ins_left[7]),
    .Y(net126));
 BUFx2_ASAP7_75t_R input127 (.A(io_ins_left[8]),
    .Y(net127));
 BUFx2_ASAP7_75t_R input128 (.A(io_ins_left[9]),
    .Y(net128));
 BUFx2_ASAP7_75t_R input129 (.A(io_ins_right[0]),
    .Y(net129));
 BUFx2_ASAP7_75t_R input130 (.A(io_ins_right[10]),
    .Y(net130));
 BUFx2_ASAP7_75t_R input131 (.A(io_ins_right[11]),
    .Y(net131));
 BUFx2_ASAP7_75t_R input132 (.A(io_ins_right[12]),
    .Y(net132));
 BUFx2_ASAP7_75t_R input133 (.A(io_ins_right[13]),
    .Y(net133));
 BUFx2_ASAP7_75t_R input134 (.A(io_ins_right[14]),
    .Y(net134));
 BUFx2_ASAP7_75t_R input135 (.A(io_ins_right[15]),
    .Y(net135));
 BUFx2_ASAP7_75t_R input136 (.A(io_ins_right[16]),
    .Y(net136));
 BUFx2_ASAP7_75t_R input137 (.A(io_ins_right[17]),
    .Y(net137));
 BUFx2_ASAP7_75t_R input138 (.A(io_ins_right[18]),
    .Y(net138));
 BUFx2_ASAP7_75t_R input139 (.A(io_ins_right[19]),
    .Y(net139));
 BUFx2_ASAP7_75t_R input140 (.A(io_ins_right[1]),
    .Y(net140));
 BUFx2_ASAP7_75t_R input141 (.A(io_ins_right[20]),
    .Y(net141));
 BUFx2_ASAP7_75t_R input142 (.A(io_ins_right[21]),
    .Y(net142));
 BUFx2_ASAP7_75t_R input143 (.A(io_ins_right[22]),
    .Y(net143));
 BUFx2_ASAP7_75t_R input144 (.A(io_ins_right[23]),
    .Y(net144));
 BUFx2_ASAP7_75t_R input145 (.A(io_ins_right[24]),
    .Y(net145));
 BUFx2_ASAP7_75t_R input146 (.A(io_ins_right[25]),
    .Y(net146));
 BUFx2_ASAP7_75t_R input147 (.A(io_ins_right[26]),
    .Y(net147));
 BUFx2_ASAP7_75t_R input148 (.A(io_ins_right[27]),
    .Y(net148));
 BUFx2_ASAP7_75t_R input149 (.A(io_ins_right[28]),
    .Y(net149));
 BUFx2_ASAP7_75t_R input150 (.A(io_ins_right[29]),
    .Y(net150));
 BUFx2_ASAP7_75t_R input151 (.A(io_ins_right[2]),
    .Y(net151));
 BUFx2_ASAP7_75t_R input152 (.A(io_ins_right[30]),
    .Y(net152));
 BUFx2_ASAP7_75t_R input153 (.A(io_ins_right[31]),
    .Y(net153));
 BUFx2_ASAP7_75t_R input154 (.A(io_ins_right[32]),
    .Y(net154));
 BUFx2_ASAP7_75t_R input155 (.A(io_ins_right[33]),
    .Y(net155));
 BUFx2_ASAP7_75t_R input156 (.A(io_ins_right[34]),
    .Y(net156));
 BUFx2_ASAP7_75t_R input157 (.A(io_ins_right[35]),
    .Y(net157));
 BUFx2_ASAP7_75t_R input158 (.A(io_ins_right[36]),
    .Y(net158));
 BUFx2_ASAP7_75t_R input159 (.A(io_ins_right[37]),
    .Y(net159));
 BUFx2_ASAP7_75t_R input160 (.A(io_ins_right[38]),
    .Y(net160));
 BUFx2_ASAP7_75t_R input161 (.A(io_ins_right[39]),
    .Y(net161));
 BUFx2_ASAP7_75t_R input162 (.A(io_ins_right[3]),
    .Y(net162));
 BUFx2_ASAP7_75t_R input163 (.A(io_ins_right[40]),
    .Y(net163));
 BUFx2_ASAP7_75t_R input164 (.A(io_ins_right[41]),
    .Y(net164));
 BUFx2_ASAP7_75t_R input165 (.A(io_ins_right[42]),
    .Y(net165));
 BUFx2_ASAP7_75t_R input166 (.A(io_ins_right[43]),
    .Y(net166));
 BUFx2_ASAP7_75t_R input167 (.A(io_ins_right[44]),
    .Y(net167));
 BUFx2_ASAP7_75t_R input168 (.A(io_ins_right[45]),
    .Y(net168));
 BUFx2_ASAP7_75t_R input169 (.A(io_ins_right[46]),
    .Y(net169));
 BUFx2_ASAP7_75t_R input170 (.A(io_ins_right[47]),
    .Y(net170));
 BUFx2_ASAP7_75t_R input171 (.A(io_ins_right[48]),
    .Y(net171));
 BUFx2_ASAP7_75t_R input172 (.A(io_ins_right[49]),
    .Y(net172));
 BUFx2_ASAP7_75t_R input173 (.A(io_ins_right[4]),
    .Y(net173));
 BUFx2_ASAP7_75t_R input174 (.A(io_ins_right[50]),
    .Y(net174));
 BUFx2_ASAP7_75t_R input175 (.A(io_ins_right[51]),
    .Y(net175));
 BUFx2_ASAP7_75t_R input176 (.A(io_ins_right[52]),
    .Y(net176));
 BUFx2_ASAP7_75t_R input177 (.A(io_ins_right[53]),
    .Y(net177));
 BUFx2_ASAP7_75t_R input178 (.A(io_ins_right[54]),
    .Y(net178));
 BUFx2_ASAP7_75t_R input179 (.A(io_ins_right[55]),
    .Y(net179));
 BUFx2_ASAP7_75t_R input180 (.A(io_ins_right[56]),
    .Y(net180));
 BUFx2_ASAP7_75t_R input181 (.A(io_ins_right[57]),
    .Y(net181));
 BUFx2_ASAP7_75t_R input182 (.A(io_ins_right[58]),
    .Y(net182));
 BUFx2_ASAP7_75t_R input183 (.A(io_ins_right[59]),
    .Y(net183));
 BUFx2_ASAP7_75t_R input184 (.A(io_ins_right[5]),
    .Y(net184));
 BUFx2_ASAP7_75t_R input185 (.A(io_ins_right[60]),
    .Y(net185));
 BUFx2_ASAP7_75t_R input186 (.A(io_ins_right[61]),
    .Y(net186));
 BUFx2_ASAP7_75t_R input187 (.A(io_ins_right[62]),
    .Y(net187));
 BUFx2_ASAP7_75t_R input188 (.A(io_ins_right[63]),
    .Y(net188));
 BUFx2_ASAP7_75t_R input189 (.A(io_ins_right[6]),
    .Y(net189));
 BUFx2_ASAP7_75t_R input190 (.A(io_ins_right[7]),
    .Y(net190));
 BUFx2_ASAP7_75t_R input191 (.A(io_ins_right[8]),
    .Y(net191));
 BUFx2_ASAP7_75t_R input192 (.A(io_ins_right[9]),
    .Y(net192));
 BUFx2_ASAP7_75t_R input193 (.A(io_ins_up[0]),
    .Y(net193));
 BUFx2_ASAP7_75t_R input194 (.A(io_ins_up[10]),
    .Y(net194));
 BUFx2_ASAP7_75t_R input195 (.A(io_ins_up[11]),
    .Y(net195));
 BUFx2_ASAP7_75t_R input196 (.A(io_ins_up[12]),
    .Y(net196));
 BUFx2_ASAP7_75t_R input197 (.A(io_ins_up[13]),
    .Y(net197));
 BUFx2_ASAP7_75t_R input198 (.A(io_ins_up[14]),
    .Y(net198));
 BUFx2_ASAP7_75t_R input199 (.A(io_ins_up[15]),
    .Y(net199));
 BUFx2_ASAP7_75t_R input200 (.A(io_ins_up[16]),
    .Y(net200));
 BUFx2_ASAP7_75t_R input201 (.A(io_ins_up[17]),
    .Y(net201));
 BUFx2_ASAP7_75t_R input202 (.A(io_ins_up[18]),
    .Y(net202));
 BUFx2_ASAP7_75t_R input203 (.A(io_ins_up[19]),
    .Y(net203));
 BUFx2_ASAP7_75t_R input204 (.A(io_ins_up[1]),
    .Y(net204));
 BUFx2_ASAP7_75t_R input205 (.A(io_ins_up[20]),
    .Y(net205));
 BUFx2_ASAP7_75t_R input206 (.A(io_ins_up[21]),
    .Y(net206));
 BUFx2_ASAP7_75t_R input207 (.A(io_ins_up[22]),
    .Y(net207));
 BUFx2_ASAP7_75t_R input208 (.A(io_ins_up[23]),
    .Y(net208));
 BUFx2_ASAP7_75t_R input209 (.A(io_ins_up[24]),
    .Y(net209));
 BUFx2_ASAP7_75t_R input210 (.A(io_ins_up[25]),
    .Y(net210));
 BUFx2_ASAP7_75t_R input211 (.A(io_ins_up[26]),
    .Y(net211));
 BUFx2_ASAP7_75t_R input212 (.A(io_ins_up[27]),
    .Y(net212));
 BUFx2_ASAP7_75t_R input213 (.A(io_ins_up[28]),
    .Y(net213));
 BUFx2_ASAP7_75t_R input214 (.A(io_ins_up[29]),
    .Y(net214));
 BUFx2_ASAP7_75t_R input215 (.A(io_ins_up[2]),
    .Y(net215));
 BUFx2_ASAP7_75t_R input216 (.A(io_ins_up[30]),
    .Y(net216));
 BUFx2_ASAP7_75t_R input217 (.A(io_ins_up[31]),
    .Y(net217));
 BUFx2_ASAP7_75t_R input218 (.A(io_ins_up[32]),
    .Y(net218));
 BUFx2_ASAP7_75t_R input219 (.A(io_ins_up[33]),
    .Y(net219));
 BUFx2_ASAP7_75t_R input220 (.A(io_ins_up[34]),
    .Y(net220));
 BUFx2_ASAP7_75t_R input221 (.A(io_ins_up[35]),
    .Y(net221));
 BUFx2_ASAP7_75t_R input222 (.A(io_ins_up[36]),
    .Y(net222));
 BUFx2_ASAP7_75t_R input223 (.A(io_ins_up[37]),
    .Y(net223));
 BUFx2_ASAP7_75t_R input224 (.A(io_ins_up[38]),
    .Y(net224));
 BUFx2_ASAP7_75t_R input225 (.A(io_ins_up[39]),
    .Y(net225));
 BUFx2_ASAP7_75t_R input226 (.A(io_ins_up[3]),
    .Y(net226));
 BUFx2_ASAP7_75t_R input227 (.A(io_ins_up[40]),
    .Y(net227));
 BUFx2_ASAP7_75t_R input228 (.A(io_ins_up[41]),
    .Y(net228));
 BUFx2_ASAP7_75t_R input229 (.A(io_ins_up[42]),
    .Y(net229));
 BUFx2_ASAP7_75t_R input230 (.A(io_ins_up[43]),
    .Y(net230));
 BUFx2_ASAP7_75t_R input231 (.A(io_ins_up[44]),
    .Y(net231));
 BUFx2_ASAP7_75t_R input232 (.A(io_ins_up[45]),
    .Y(net232));
 BUFx2_ASAP7_75t_R input233 (.A(io_ins_up[46]),
    .Y(net233));
 BUFx2_ASAP7_75t_R input234 (.A(io_ins_up[47]),
    .Y(net234));
 BUFx2_ASAP7_75t_R input235 (.A(io_ins_up[48]),
    .Y(net235));
 BUFx2_ASAP7_75t_R input236 (.A(io_ins_up[49]),
    .Y(net236));
 BUFx2_ASAP7_75t_R input237 (.A(io_ins_up[4]),
    .Y(net237));
 BUFx2_ASAP7_75t_R input238 (.A(io_ins_up[50]),
    .Y(net238));
 BUFx2_ASAP7_75t_R input239 (.A(io_ins_up[51]),
    .Y(net239));
 BUFx2_ASAP7_75t_R input240 (.A(io_ins_up[52]),
    .Y(net240));
 BUFx2_ASAP7_75t_R input241 (.A(io_ins_up[53]),
    .Y(net241));
 BUFx2_ASAP7_75t_R input242 (.A(io_ins_up[54]),
    .Y(net242));
 BUFx2_ASAP7_75t_R input243 (.A(io_ins_up[55]),
    .Y(net243));
 BUFx2_ASAP7_75t_R input244 (.A(io_ins_up[56]),
    .Y(net244));
 BUFx2_ASAP7_75t_R input245 (.A(io_ins_up[57]),
    .Y(net245));
 BUFx2_ASAP7_75t_R input246 (.A(io_ins_up[58]),
    .Y(net246));
 BUFx2_ASAP7_75t_R input247 (.A(io_ins_up[59]),
    .Y(net247));
 BUFx2_ASAP7_75t_R input248 (.A(io_ins_up[5]),
    .Y(net248));
 BUFx2_ASAP7_75t_R input249 (.A(io_ins_up[60]),
    .Y(net249));
 BUFx2_ASAP7_75t_R input250 (.A(io_ins_up[61]),
    .Y(net250));
 BUFx2_ASAP7_75t_R input251 (.A(io_ins_up[62]),
    .Y(net251));
 BUFx2_ASAP7_75t_R input252 (.A(io_ins_up[63]),
    .Y(net252));
 BUFx2_ASAP7_75t_R input253 (.A(io_ins_up[6]),
    .Y(net253));
 BUFx2_ASAP7_75t_R input254 (.A(io_ins_up[7]),
    .Y(net254));
 BUFx2_ASAP7_75t_R input255 (.A(io_ins_up[8]),
    .Y(net255));
 BUFx2_ASAP7_75t_R input256 (.A(io_ins_up[9]),
    .Y(net256));
 BUFx2_ASAP7_75t_R input257 (.A(io_lsbIns_4),
    .Y(net257));
 BUFx2_ASAP7_75t_R output258 (.A(net258),
    .Y(io_lsbOuts_0));
 BUFx2_ASAP7_75t_R output259 (.A(net259),
    .Y(io_lsbOuts_1));
 BUFx2_ASAP7_75t_R output260 (.A(net260),
    .Y(io_lsbOuts_2));
 BUFx2_ASAP7_75t_R output261 (.A(net261),
    .Y(io_lsbOuts_3));
 BUFx2_ASAP7_75t_R output262 (.A(net262),
    .Y(io_lsbOuts_4));
 BUFx2_ASAP7_75t_R output263 (.A(net263),
    .Y(io_lsbOuts_5));
 BUFx2_ASAP7_75t_R output264 (.A(net264),
    .Y(io_lsbOuts_6));
 BUFx2_ASAP7_75t_R output265 (.A(net265),
    .Y(io_lsbOuts_7));
 BUFx2_ASAP7_75t_R output266 (.A(net266),
    .Y(io_outs_down[0]));
 BUFx2_ASAP7_75t_R output267 (.A(net267),
    .Y(io_outs_down[10]));
 BUFx2_ASAP7_75t_R output268 (.A(net268),
    .Y(io_outs_down[11]));
 BUFx2_ASAP7_75t_R output269 (.A(net269),
    .Y(io_outs_down[12]));
 BUFx2_ASAP7_75t_R output270 (.A(net270),
    .Y(io_outs_down[13]));
 BUFx2_ASAP7_75t_R output271 (.A(net271),
    .Y(io_outs_down[14]));
 BUFx2_ASAP7_75t_R output272 (.A(net272),
    .Y(io_outs_down[15]));
 BUFx2_ASAP7_75t_R output273 (.A(net273),
    .Y(io_outs_down[16]));
 BUFx2_ASAP7_75t_R output274 (.A(net274),
    .Y(io_outs_down[17]));
 BUFx2_ASAP7_75t_R output275 (.A(net275),
    .Y(io_outs_down[18]));
 BUFx2_ASAP7_75t_R output276 (.A(net276),
    .Y(io_outs_down[19]));
 BUFx2_ASAP7_75t_R output277 (.A(net277),
    .Y(io_outs_down[1]));
 BUFx2_ASAP7_75t_R output278 (.A(net278),
    .Y(io_outs_down[20]));
 BUFx2_ASAP7_75t_R output279 (.A(net279),
    .Y(io_outs_down[21]));
 BUFx2_ASAP7_75t_R output280 (.A(net280),
    .Y(io_outs_down[22]));
 BUFx2_ASAP7_75t_R output281 (.A(net281),
    .Y(io_outs_down[23]));
 BUFx2_ASAP7_75t_R output282 (.A(net282),
    .Y(io_outs_down[24]));
 BUFx2_ASAP7_75t_R output283 (.A(net283),
    .Y(io_outs_down[25]));
 BUFx2_ASAP7_75t_R output284 (.A(net284),
    .Y(io_outs_down[26]));
 BUFx2_ASAP7_75t_R output285 (.A(net285),
    .Y(io_outs_down[27]));
 BUFx2_ASAP7_75t_R output286 (.A(net286),
    .Y(io_outs_down[28]));
 BUFx2_ASAP7_75t_R output287 (.A(net287),
    .Y(io_outs_down[29]));
 BUFx2_ASAP7_75t_R output288 (.A(net288),
    .Y(io_outs_down[2]));
 BUFx2_ASAP7_75t_R output289 (.A(net289),
    .Y(io_outs_down[30]));
 BUFx2_ASAP7_75t_R output290 (.A(net290),
    .Y(io_outs_down[31]));
 BUFx2_ASAP7_75t_R output291 (.A(net291),
    .Y(io_outs_down[32]));
 BUFx2_ASAP7_75t_R output292 (.A(net292),
    .Y(io_outs_down[33]));
 BUFx2_ASAP7_75t_R output293 (.A(net293),
    .Y(io_outs_down[34]));
 BUFx2_ASAP7_75t_R output294 (.A(net294),
    .Y(io_outs_down[35]));
 BUFx2_ASAP7_75t_R output295 (.A(net295),
    .Y(io_outs_down[36]));
 BUFx2_ASAP7_75t_R output296 (.A(net296),
    .Y(io_outs_down[37]));
 BUFx2_ASAP7_75t_R output297 (.A(net297),
    .Y(io_outs_down[38]));
 BUFx2_ASAP7_75t_R output298 (.A(net298),
    .Y(io_outs_down[39]));
 BUFx2_ASAP7_75t_R output299 (.A(net299),
    .Y(io_outs_down[3]));
 BUFx2_ASAP7_75t_R output300 (.A(net300),
    .Y(io_outs_down[40]));
 BUFx2_ASAP7_75t_R output301 (.A(net301),
    .Y(io_outs_down[41]));
 BUFx2_ASAP7_75t_R output302 (.A(net302),
    .Y(io_outs_down[42]));
 BUFx2_ASAP7_75t_R output303 (.A(net303),
    .Y(io_outs_down[43]));
 BUFx2_ASAP7_75t_R output304 (.A(net304),
    .Y(io_outs_down[44]));
 BUFx2_ASAP7_75t_R output305 (.A(net305),
    .Y(io_outs_down[45]));
 BUFx2_ASAP7_75t_R output306 (.A(net306),
    .Y(io_outs_down[46]));
 BUFx2_ASAP7_75t_R output307 (.A(net307),
    .Y(io_outs_down[47]));
 BUFx2_ASAP7_75t_R output308 (.A(net308),
    .Y(io_outs_down[48]));
 BUFx2_ASAP7_75t_R output309 (.A(net309),
    .Y(io_outs_down[49]));
 BUFx2_ASAP7_75t_R output310 (.A(net310),
    .Y(io_outs_down[4]));
 BUFx2_ASAP7_75t_R output311 (.A(net311),
    .Y(io_outs_down[50]));
 BUFx2_ASAP7_75t_R output312 (.A(net312),
    .Y(io_outs_down[51]));
 BUFx2_ASAP7_75t_R output313 (.A(net313),
    .Y(io_outs_down[52]));
 BUFx2_ASAP7_75t_R output314 (.A(net314),
    .Y(io_outs_down[53]));
 BUFx2_ASAP7_75t_R output315 (.A(net315),
    .Y(io_outs_down[54]));
 BUFx2_ASAP7_75t_R output316 (.A(net316),
    .Y(io_outs_down[55]));
 BUFx2_ASAP7_75t_R output317 (.A(net317),
    .Y(io_outs_down[56]));
 BUFx2_ASAP7_75t_R output318 (.A(net318),
    .Y(io_outs_down[57]));
 BUFx2_ASAP7_75t_R output319 (.A(net319),
    .Y(io_outs_down[58]));
 BUFx2_ASAP7_75t_R output320 (.A(net320),
    .Y(io_outs_down[59]));
 BUFx2_ASAP7_75t_R output321 (.A(net321),
    .Y(io_outs_down[5]));
 BUFx2_ASAP7_75t_R output322 (.A(net322),
    .Y(io_outs_down[60]));
 BUFx2_ASAP7_75t_R output323 (.A(net323),
    .Y(io_outs_down[61]));
 BUFx2_ASAP7_75t_R output324 (.A(net324),
    .Y(io_outs_down[62]));
 BUFx2_ASAP7_75t_R output325 (.A(net325),
    .Y(io_outs_down[63]));
 BUFx2_ASAP7_75t_R output326 (.A(net326),
    .Y(io_outs_down[6]));
 BUFx2_ASAP7_75t_R output327 (.A(net327),
    .Y(io_outs_down[7]));
 BUFx2_ASAP7_75t_R output328 (.A(net328),
    .Y(io_outs_down[8]));
 BUFx2_ASAP7_75t_R output329 (.A(net329),
    .Y(io_outs_down[9]));
 BUFx2_ASAP7_75t_R output330 (.A(net330),
    .Y(io_outs_left[0]));
 BUFx2_ASAP7_75t_R output331 (.A(net331),
    .Y(io_outs_left[10]));
 BUFx2_ASAP7_75t_R output332 (.A(net332),
    .Y(io_outs_left[11]));
 BUFx2_ASAP7_75t_R output333 (.A(net333),
    .Y(io_outs_left[12]));
 BUFx2_ASAP7_75t_R output334 (.A(net334),
    .Y(io_outs_left[13]));
 BUFx2_ASAP7_75t_R output335 (.A(net335),
    .Y(io_outs_left[14]));
 BUFx2_ASAP7_75t_R output336 (.A(net336),
    .Y(io_outs_left[15]));
 BUFx2_ASAP7_75t_R output337 (.A(net337),
    .Y(io_outs_left[16]));
 BUFx2_ASAP7_75t_R output338 (.A(net338),
    .Y(io_outs_left[17]));
 BUFx2_ASAP7_75t_R output339 (.A(net339),
    .Y(io_outs_left[18]));
 BUFx2_ASAP7_75t_R output340 (.A(net340),
    .Y(io_outs_left[19]));
 BUFx2_ASAP7_75t_R output341 (.A(net341),
    .Y(io_outs_left[1]));
 BUFx2_ASAP7_75t_R output342 (.A(net342),
    .Y(io_outs_left[20]));
 BUFx2_ASAP7_75t_R output343 (.A(net343),
    .Y(io_outs_left[21]));
 BUFx2_ASAP7_75t_R output344 (.A(net344),
    .Y(io_outs_left[22]));
 BUFx2_ASAP7_75t_R output345 (.A(net345),
    .Y(io_outs_left[23]));
 BUFx2_ASAP7_75t_R output346 (.A(net346),
    .Y(io_outs_left[24]));
 BUFx2_ASAP7_75t_R output347 (.A(net347),
    .Y(io_outs_left[25]));
 BUFx2_ASAP7_75t_R output348 (.A(net348),
    .Y(io_outs_left[26]));
 BUFx2_ASAP7_75t_R output349 (.A(net349),
    .Y(io_outs_left[27]));
 BUFx2_ASAP7_75t_R output350 (.A(net350),
    .Y(io_outs_left[28]));
 BUFx2_ASAP7_75t_R output351 (.A(net351),
    .Y(io_outs_left[29]));
 BUFx2_ASAP7_75t_R output352 (.A(net352),
    .Y(io_outs_left[2]));
 BUFx2_ASAP7_75t_R output353 (.A(net353),
    .Y(io_outs_left[30]));
 BUFx2_ASAP7_75t_R output354 (.A(net354),
    .Y(io_outs_left[31]));
 BUFx2_ASAP7_75t_R output355 (.A(net355),
    .Y(io_outs_left[32]));
 BUFx2_ASAP7_75t_R output356 (.A(net356),
    .Y(io_outs_left[33]));
 BUFx2_ASAP7_75t_R output357 (.A(net357),
    .Y(io_outs_left[34]));
 BUFx2_ASAP7_75t_R output358 (.A(net358),
    .Y(io_outs_left[35]));
 BUFx2_ASAP7_75t_R output359 (.A(net359),
    .Y(io_outs_left[36]));
 BUFx2_ASAP7_75t_R output360 (.A(net360),
    .Y(io_outs_left[37]));
 BUFx2_ASAP7_75t_R output361 (.A(net361),
    .Y(io_outs_left[38]));
 BUFx2_ASAP7_75t_R output362 (.A(net362),
    .Y(io_outs_left[39]));
 BUFx2_ASAP7_75t_R output363 (.A(net363),
    .Y(io_outs_left[3]));
 BUFx2_ASAP7_75t_R output364 (.A(net364),
    .Y(io_outs_left[40]));
 BUFx2_ASAP7_75t_R output365 (.A(net365),
    .Y(io_outs_left[41]));
 BUFx2_ASAP7_75t_R output366 (.A(net366),
    .Y(io_outs_left[42]));
 BUFx2_ASAP7_75t_R output367 (.A(net367),
    .Y(io_outs_left[43]));
 BUFx2_ASAP7_75t_R output368 (.A(net368),
    .Y(io_outs_left[44]));
 BUFx2_ASAP7_75t_R output369 (.A(net369),
    .Y(io_outs_left[45]));
 BUFx2_ASAP7_75t_R output370 (.A(net370),
    .Y(io_outs_left[46]));
 BUFx2_ASAP7_75t_R output371 (.A(net371),
    .Y(io_outs_left[47]));
 BUFx2_ASAP7_75t_R output372 (.A(net372),
    .Y(io_outs_left[48]));
 BUFx2_ASAP7_75t_R output373 (.A(net373),
    .Y(io_outs_left[49]));
 BUFx2_ASAP7_75t_R output374 (.A(net374),
    .Y(io_outs_left[4]));
 BUFx2_ASAP7_75t_R output375 (.A(net375),
    .Y(io_outs_left[50]));
 BUFx2_ASAP7_75t_R output376 (.A(net376),
    .Y(io_outs_left[51]));
 BUFx2_ASAP7_75t_R output377 (.A(net377),
    .Y(io_outs_left[52]));
 BUFx2_ASAP7_75t_R output378 (.A(net378),
    .Y(io_outs_left[53]));
 BUFx2_ASAP7_75t_R output379 (.A(net379),
    .Y(io_outs_left[54]));
 BUFx2_ASAP7_75t_R output380 (.A(net380),
    .Y(io_outs_left[55]));
 BUFx2_ASAP7_75t_R output381 (.A(net381),
    .Y(io_outs_left[56]));
 BUFx2_ASAP7_75t_R output382 (.A(net382),
    .Y(io_outs_left[57]));
 BUFx2_ASAP7_75t_R output383 (.A(net383),
    .Y(io_outs_left[58]));
 BUFx2_ASAP7_75t_R output384 (.A(net384),
    .Y(io_outs_left[59]));
 BUFx2_ASAP7_75t_R output385 (.A(net385),
    .Y(io_outs_left[5]));
 BUFx2_ASAP7_75t_R output386 (.A(net386),
    .Y(io_outs_left[60]));
 BUFx2_ASAP7_75t_R output387 (.A(net387),
    .Y(io_outs_left[61]));
 BUFx2_ASAP7_75t_R output388 (.A(net388),
    .Y(io_outs_left[62]));
 BUFx2_ASAP7_75t_R output389 (.A(net389),
    .Y(io_outs_left[63]));
 BUFx2_ASAP7_75t_R output390 (.A(net390),
    .Y(io_outs_left[6]));
 BUFx2_ASAP7_75t_R output391 (.A(net391),
    .Y(io_outs_left[7]));
 BUFx2_ASAP7_75t_R output392 (.A(net392),
    .Y(io_outs_left[8]));
 BUFx2_ASAP7_75t_R output393 (.A(net393),
    .Y(io_outs_left[9]));
 BUFx2_ASAP7_75t_R output394 (.A(net394),
    .Y(io_outs_right[0]));
 BUFx2_ASAP7_75t_R output395 (.A(net395),
    .Y(io_outs_right[10]));
 BUFx2_ASAP7_75t_R output396 (.A(net396),
    .Y(io_outs_right[11]));
 BUFx2_ASAP7_75t_R output397 (.A(net397),
    .Y(io_outs_right[12]));
 BUFx2_ASAP7_75t_R output398 (.A(net398),
    .Y(io_outs_right[13]));
 BUFx2_ASAP7_75t_R output399 (.A(net399),
    .Y(io_outs_right[14]));
 BUFx2_ASAP7_75t_R output400 (.A(net400),
    .Y(io_outs_right[15]));
 BUFx2_ASAP7_75t_R output401 (.A(net401),
    .Y(io_outs_right[16]));
 BUFx2_ASAP7_75t_R output402 (.A(net402),
    .Y(io_outs_right[17]));
 BUFx2_ASAP7_75t_R output403 (.A(net403),
    .Y(io_outs_right[18]));
 BUFx2_ASAP7_75t_R output404 (.A(net404),
    .Y(io_outs_right[19]));
 BUFx2_ASAP7_75t_R output405 (.A(net405),
    .Y(io_outs_right[1]));
 BUFx2_ASAP7_75t_R output406 (.A(net406),
    .Y(io_outs_right[20]));
 BUFx2_ASAP7_75t_R output407 (.A(net407),
    .Y(io_outs_right[21]));
 BUFx2_ASAP7_75t_R output408 (.A(net408),
    .Y(io_outs_right[22]));
 BUFx2_ASAP7_75t_R output409 (.A(net409),
    .Y(io_outs_right[23]));
 BUFx2_ASAP7_75t_R output410 (.A(net410),
    .Y(io_outs_right[24]));
 BUFx2_ASAP7_75t_R output411 (.A(net411),
    .Y(io_outs_right[25]));
 BUFx2_ASAP7_75t_R output412 (.A(net412),
    .Y(io_outs_right[26]));
 BUFx2_ASAP7_75t_R output413 (.A(net413),
    .Y(io_outs_right[27]));
 BUFx2_ASAP7_75t_R output414 (.A(net414),
    .Y(io_outs_right[28]));
 BUFx2_ASAP7_75t_R output415 (.A(net415),
    .Y(io_outs_right[29]));
 BUFx2_ASAP7_75t_R output416 (.A(net416),
    .Y(io_outs_right[2]));
 BUFx2_ASAP7_75t_R output417 (.A(net417),
    .Y(io_outs_right[30]));
 BUFx2_ASAP7_75t_R output418 (.A(net418),
    .Y(io_outs_right[31]));
 BUFx2_ASAP7_75t_R output419 (.A(net419),
    .Y(io_outs_right[32]));
 BUFx2_ASAP7_75t_R output420 (.A(net420),
    .Y(io_outs_right[33]));
 BUFx2_ASAP7_75t_R output421 (.A(net421),
    .Y(io_outs_right[34]));
 BUFx2_ASAP7_75t_R output422 (.A(net422),
    .Y(io_outs_right[35]));
 BUFx2_ASAP7_75t_R output423 (.A(net423),
    .Y(io_outs_right[36]));
 BUFx2_ASAP7_75t_R output424 (.A(net424),
    .Y(io_outs_right[37]));
 BUFx2_ASAP7_75t_R output425 (.A(net425),
    .Y(io_outs_right[38]));
 BUFx2_ASAP7_75t_R output426 (.A(net426),
    .Y(io_outs_right[39]));
 BUFx2_ASAP7_75t_R output427 (.A(net427),
    .Y(io_outs_right[3]));
 BUFx2_ASAP7_75t_R output428 (.A(net428),
    .Y(io_outs_right[40]));
 BUFx2_ASAP7_75t_R output429 (.A(net429),
    .Y(io_outs_right[41]));
 BUFx2_ASAP7_75t_R output430 (.A(net430),
    .Y(io_outs_right[42]));
 BUFx2_ASAP7_75t_R output431 (.A(net431),
    .Y(io_outs_right[43]));
 BUFx2_ASAP7_75t_R output432 (.A(net432),
    .Y(io_outs_right[44]));
 BUFx2_ASAP7_75t_R output433 (.A(net433),
    .Y(io_outs_right[45]));
 BUFx2_ASAP7_75t_R output434 (.A(net434),
    .Y(io_outs_right[46]));
 BUFx2_ASAP7_75t_R output435 (.A(net435),
    .Y(io_outs_right[47]));
 BUFx2_ASAP7_75t_R output436 (.A(net436),
    .Y(io_outs_right[48]));
 BUFx2_ASAP7_75t_R output437 (.A(net437),
    .Y(io_outs_right[49]));
 BUFx2_ASAP7_75t_R output438 (.A(net438),
    .Y(io_outs_right[4]));
 BUFx2_ASAP7_75t_R output439 (.A(net439),
    .Y(io_outs_right[50]));
 BUFx2_ASAP7_75t_R output440 (.A(net440),
    .Y(io_outs_right[51]));
 BUFx2_ASAP7_75t_R output441 (.A(net441),
    .Y(io_outs_right[52]));
 BUFx2_ASAP7_75t_R output442 (.A(net442),
    .Y(io_outs_right[53]));
 BUFx2_ASAP7_75t_R output443 (.A(net443),
    .Y(io_outs_right[54]));
 BUFx2_ASAP7_75t_R output444 (.A(net444),
    .Y(io_outs_right[55]));
 BUFx2_ASAP7_75t_R output445 (.A(net445),
    .Y(io_outs_right[56]));
 BUFx2_ASAP7_75t_R output446 (.A(net446),
    .Y(io_outs_right[57]));
 BUFx2_ASAP7_75t_R output447 (.A(net447),
    .Y(io_outs_right[58]));
 BUFx2_ASAP7_75t_R output448 (.A(net448),
    .Y(io_outs_right[59]));
 BUFx2_ASAP7_75t_R output449 (.A(net449),
    .Y(io_outs_right[5]));
 BUFx2_ASAP7_75t_R output450 (.A(net450),
    .Y(io_outs_right[60]));
 BUFx2_ASAP7_75t_R output451 (.A(net451),
    .Y(io_outs_right[61]));
 BUFx2_ASAP7_75t_R output452 (.A(net452),
    .Y(io_outs_right[62]));
 BUFx2_ASAP7_75t_R output453 (.A(net453),
    .Y(io_outs_right[63]));
 BUFx2_ASAP7_75t_R output454 (.A(net454),
    .Y(io_outs_right[6]));
 BUFx2_ASAP7_75t_R output455 (.A(net455),
    .Y(io_outs_right[7]));
 BUFx2_ASAP7_75t_R output456 (.A(net456),
    .Y(io_outs_right[8]));
 BUFx2_ASAP7_75t_R output457 (.A(net457),
    .Y(io_outs_right[9]));
 BUFx2_ASAP7_75t_R output458 (.A(net458),
    .Y(io_outs_up[0]));
 BUFx2_ASAP7_75t_R output459 (.A(net459),
    .Y(io_outs_up[10]));
 BUFx2_ASAP7_75t_R output460 (.A(net460),
    .Y(io_outs_up[11]));
 BUFx2_ASAP7_75t_R output461 (.A(net461),
    .Y(io_outs_up[12]));
 BUFx2_ASAP7_75t_R output462 (.A(net462),
    .Y(io_outs_up[13]));
 BUFx2_ASAP7_75t_R output463 (.A(net463),
    .Y(io_outs_up[14]));
 BUFx2_ASAP7_75t_R output464 (.A(net464),
    .Y(io_outs_up[15]));
 BUFx2_ASAP7_75t_R output465 (.A(net465),
    .Y(io_outs_up[16]));
 BUFx2_ASAP7_75t_R output466 (.A(net466),
    .Y(io_outs_up[17]));
 BUFx2_ASAP7_75t_R output467 (.A(net467),
    .Y(io_outs_up[18]));
 BUFx2_ASAP7_75t_R output468 (.A(net468),
    .Y(io_outs_up[19]));
 BUFx2_ASAP7_75t_R output469 (.A(net469),
    .Y(io_outs_up[1]));
 BUFx2_ASAP7_75t_R output470 (.A(net470),
    .Y(io_outs_up[20]));
 BUFx2_ASAP7_75t_R output471 (.A(net471),
    .Y(io_outs_up[21]));
 BUFx2_ASAP7_75t_R output472 (.A(net472),
    .Y(io_outs_up[22]));
 BUFx2_ASAP7_75t_R output473 (.A(net473),
    .Y(io_outs_up[23]));
 BUFx2_ASAP7_75t_R output474 (.A(net474),
    .Y(io_outs_up[24]));
 BUFx2_ASAP7_75t_R output475 (.A(net475),
    .Y(io_outs_up[25]));
 BUFx2_ASAP7_75t_R output476 (.A(net476),
    .Y(io_outs_up[26]));
 BUFx2_ASAP7_75t_R output477 (.A(net477),
    .Y(io_outs_up[27]));
 BUFx2_ASAP7_75t_R output478 (.A(net478),
    .Y(io_outs_up[28]));
 BUFx2_ASAP7_75t_R output479 (.A(net479),
    .Y(io_outs_up[29]));
 BUFx2_ASAP7_75t_R output480 (.A(net480),
    .Y(io_outs_up[2]));
 BUFx2_ASAP7_75t_R output481 (.A(net481),
    .Y(io_outs_up[30]));
 BUFx2_ASAP7_75t_R output482 (.A(net482),
    .Y(io_outs_up[31]));
 BUFx2_ASAP7_75t_R output483 (.A(net483),
    .Y(io_outs_up[32]));
 BUFx2_ASAP7_75t_R output484 (.A(net484),
    .Y(io_outs_up[33]));
 BUFx2_ASAP7_75t_R output485 (.A(net485),
    .Y(io_outs_up[34]));
 BUFx2_ASAP7_75t_R output486 (.A(net486),
    .Y(io_outs_up[35]));
 BUFx2_ASAP7_75t_R output487 (.A(net487),
    .Y(io_outs_up[36]));
 BUFx2_ASAP7_75t_R output488 (.A(net488),
    .Y(io_outs_up[37]));
 BUFx2_ASAP7_75t_R output489 (.A(net489),
    .Y(io_outs_up[38]));
 BUFx2_ASAP7_75t_R output490 (.A(net490),
    .Y(io_outs_up[39]));
 BUFx2_ASAP7_75t_R output491 (.A(net491),
    .Y(io_outs_up[3]));
 BUFx2_ASAP7_75t_R output492 (.A(net492),
    .Y(io_outs_up[40]));
 BUFx2_ASAP7_75t_R output493 (.A(net493),
    .Y(io_outs_up[41]));
 BUFx2_ASAP7_75t_R output494 (.A(net494),
    .Y(io_outs_up[42]));
 BUFx2_ASAP7_75t_R output495 (.A(net495),
    .Y(io_outs_up[43]));
 BUFx2_ASAP7_75t_R output496 (.A(net496),
    .Y(io_outs_up[44]));
 BUFx2_ASAP7_75t_R output497 (.A(net497),
    .Y(io_outs_up[45]));
 BUFx2_ASAP7_75t_R output498 (.A(net498),
    .Y(io_outs_up[46]));
 BUFx2_ASAP7_75t_R output499 (.A(net499),
    .Y(io_outs_up[47]));
 BUFx2_ASAP7_75t_R output500 (.A(net500),
    .Y(io_outs_up[48]));
 BUFx2_ASAP7_75t_R output501 (.A(net501),
    .Y(io_outs_up[49]));
 BUFx2_ASAP7_75t_R output502 (.A(net502),
    .Y(io_outs_up[4]));
 BUFx2_ASAP7_75t_R output503 (.A(net503),
    .Y(io_outs_up[50]));
 BUFx2_ASAP7_75t_R output504 (.A(net504),
    .Y(io_outs_up[51]));
 BUFx2_ASAP7_75t_R output505 (.A(net505),
    .Y(io_outs_up[52]));
 BUFx2_ASAP7_75t_R output506 (.A(net506),
    .Y(io_outs_up[53]));
 BUFx2_ASAP7_75t_R output507 (.A(net507),
    .Y(io_outs_up[54]));
 BUFx2_ASAP7_75t_R output508 (.A(net508),
    .Y(io_outs_up[55]));
 BUFx2_ASAP7_75t_R output509 (.A(net509),
    .Y(io_outs_up[56]));
 BUFx2_ASAP7_75t_R output510 (.A(net510),
    .Y(io_outs_up[57]));
 BUFx2_ASAP7_75t_R output511 (.A(net511),
    .Y(io_outs_up[58]));
 BUFx2_ASAP7_75t_R output512 (.A(net512),
    .Y(io_outs_up[59]));
 BUFx2_ASAP7_75t_R output513 (.A(net513),
    .Y(io_outs_up[5]));
 BUFx2_ASAP7_75t_R output514 (.A(net514),
    .Y(io_outs_up[60]));
 BUFx2_ASAP7_75t_R output515 (.A(net515),
    .Y(io_outs_up[61]));
 BUFx2_ASAP7_75t_R output516 (.A(net516),
    .Y(io_outs_up[62]));
 BUFx2_ASAP7_75t_R output517 (.A(net517),
    .Y(io_outs_up[63]));
 BUFx2_ASAP7_75t_R output518 (.A(net518),
    .Y(io_outs_up[6]));
 BUFx2_ASAP7_75t_R output519 (.A(net519),
    .Y(io_outs_up[7]));
 BUFx2_ASAP7_75t_R output520 (.A(net520),
    .Y(io_outs_up[8]));
 BUFx2_ASAP7_75t_R output521 (.A(net521),
    .Y(io_outs_up[9]));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_0_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_0_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_1_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_1_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_2_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_2_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_3_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_3_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_4_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_4_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_5_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_5_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_6_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_6_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_7_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_7_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_8_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_8_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_9_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_9_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_10_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_10_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_11_clock (.A(clknet_1_1__leaf_clock),
    .Y(clknet_leaf_11_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_12_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_12_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_13_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_13_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_14_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_14_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_15_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_15_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_16_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_16_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_17_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_17_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_18_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_18_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_19_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_19_clock));
 BUFx16f_ASAP7_75t_R clkbuf_leaf_20_clock (.A(clknet_1_0__leaf_clock),
    .Y(clknet_leaf_20_clock));
 BUFx8_ASAP7_75t_R clkbuf_0_clock (.A(clock),
    .Y(clknet_0_clock));
 BUFx8_ASAP7_75t_R clkbuf_1_0__f_clock (.A(clknet_0_clock),
    .Y(clknet_1_0__leaf_clock));
 BUFx8_ASAP7_75t_R clkbuf_1_1__f_clock (.A(clknet_0_clock),
    .Y(clknet_1_1__leaf_clock));
 BUFx16f_ASAP7_75t_R clkload0 (.A(clknet_1_1__leaf_clock));
 INVxp67_ASAP7_75t_R clkload1 (.A(clknet_leaf_0_clock));
 INVxp33_ASAP7_75t_R clkload2 (.A(clknet_leaf_1_clock));
 BUFx4f_ASAP7_75t_R clkload3 (.A(clknet_leaf_12_clock));
 BUFx12_ASAP7_75t_R clkload4 (.A(clknet_leaf_13_clock));
 CKINVDCx10_ASAP7_75t_R clkload5 (.A(clknet_leaf_14_clock));
 INVxp33_ASAP7_75t_R clkload6 (.A(clknet_leaf_15_clock));
 INVxp67_ASAP7_75t_R clkload7 (.A(clknet_leaf_16_clock));
 BUFx12_ASAP7_75t_R clkload8 (.A(clknet_leaf_17_clock));
 INVxp67_ASAP7_75t_R clkload9 (.A(clknet_leaf_19_clock));
 CKINVDCx12_ASAP7_75t_R clkload10 (.A(clknet_leaf_20_clock));
 BUFx12_ASAP7_75t_R clkload11 (.A(clknet_leaf_2_clock));
 BUFx4f_ASAP7_75t_R clkload12 (.A(clknet_leaf_3_clock));
 INVx13_ASAP7_75t_R clkload13 (.A(clknet_leaf_4_clock));
 INVx6_ASAP7_75t_R clkload14 (.A(clknet_leaf_5_clock));
 INVxp67_ASAP7_75t_R clkload15 (.A(clknet_leaf_6_clock));
 BUFx4f_ASAP7_75t_R clkload16 (.A(clknet_leaf_8_clock));
 CKINVDCx6p67_ASAP7_75t_R clkload17 (.A(clknet_leaf_9_clock));
 INVxp67_ASAP7_75t_R clkload18 (.A(clknet_leaf_10_clock));
 BUFx24_ASAP7_75t_R clkload19 (.A(clknet_leaf_11_clock));
 DECAPx10_ASAP7_75t_R FILLER_0_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_222 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_254 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_304 ();
 FILLER_ASAP7_75t_R FILLER_0_0_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_519 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_541 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_563 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_585 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_607 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_629 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_651 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_673 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_695 ();
 DECAPx10_ASAP7_75t_R FILLER_0_0_717 ();
 DECAPx6_ASAP7_75t_R FILLER_0_0_739 ();
 DECAPx1_ASAP7_75t_R FILLER_0_0_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_0_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_222 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_322 ();
 FILLER_ASAP7_75t_R FILLER_0_1_397 ();
 FILLER_ASAP7_75t_R FILLER_0_1_409 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_438 ();
 DECAPx1_ASAP7_75t_R FILLER_0_1_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_500 ();
 DECAPx2_ASAP7_75t_R FILLER_0_1_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_517 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_523 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_611 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_633 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_677 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_699 ();
 DECAPx10_ASAP7_75t_R FILLER_0_1_721 ();
 DECAPx6_ASAP7_75t_R FILLER_0_1_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_1_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_222 ();
 DECAPx4_ASAP7_75t_R FILLER_0_2_244 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_304 ();
 FILLER_ASAP7_75t_R FILLER_0_2_339 ();
 FILLER_ASAP7_75t_R FILLER_0_2_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_416 ();
 FILLER_ASAP7_75t_R FILLER_0_2_422 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_438 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_454 ();
 FILLER_ASAP7_75t_R FILLER_0_2_460 ();
 DECAPx1_ASAP7_75t_R FILLER_0_2_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_2_468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_2_730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_2_752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_222 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_258 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_272 ();
 FILLER_ASAP7_75t_R FILLER_0_3_278 ();
 DECAPx1_ASAP7_75t_R FILLER_0_3_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_320 ();
 FILLER_ASAP7_75t_R FILLER_0_3_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_331 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_337 ();
 FILLER_ASAP7_75t_R FILLER_0_3_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_357 ();
 DECAPx4_ASAP7_75t_R FILLER_0_3_363 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_396 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_444 ();
 FILLER_ASAP7_75t_R FILLER_0_3_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_3_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_496 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_518 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_540 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_562 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_584 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_606 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_672 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_694 ();
 DECAPx10_ASAP7_75t_R FILLER_0_3_716 ();
 DECAPx6_ASAP7_75t_R FILLER_0_3_738 ();
 DECAPx2_ASAP7_75t_R FILLER_0_3_752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_222 ();
 DECAPx4_ASAP7_75t_R FILLER_0_4_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_254 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_284 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_305 ();
 FILLER_ASAP7_75t_R FILLER_0_4_319 ();
 FILLER_ASAP7_75t_R FILLER_0_4_326 ();
 DECAPx4_ASAP7_75t_R FILLER_0_4_333 ();
 FILLER_ASAP7_75t_R FILLER_0_4_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_4_345 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_370 ();
 FILLER_ASAP7_75t_R FILLER_0_4_376 ();
 FILLER_ASAP7_75t_R FILLER_0_4_388 ();
 DECAPx6_ASAP7_75t_R FILLER_0_4_393 ();
 FILLER_ASAP7_75t_R FILLER_0_4_407 ();
 DECAPx2_ASAP7_75t_R FILLER_0_4_430 ();
 DECAPx1_ASAP7_75t_R FILLER_0_4_464 ();
 FILLER_ASAP7_75t_R FILLER_0_4_471 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_494 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_516 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_560 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_604 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_626 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_648 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_670 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_692 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_714 ();
 DECAPx10_ASAP7_75t_R FILLER_0_4_736 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_244 ();
 DECAPx4_ASAP7_75t_R FILLER_0_5_266 ();
 FILLER_ASAP7_75t_R FILLER_0_5_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_278 ();
 DECAPx4_ASAP7_75t_R FILLER_0_5_287 ();
 FILLER_ASAP7_75t_R FILLER_0_5_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_309 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_335 ();
 FILLER_ASAP7_75t_R FILLER_0_5_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_408 ();
 DECAPx2_ASAP7_75t_R FILLER_0_5_412 ();
 FILLER_ASAP7_75t_R FILLER_0_5_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_5_456 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_5_718 ();
 DECAPx6_ASAP7_75t_R FILLER_0_5_740 ();
 DECAPx1_ASAP7_75t_R FILLER_0_5_754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_266 ();
 DECAPx1_ASAP7_75t_R FILLER_0_6_280 ();
 DECAPx4_ASAP7_75t_R FILLER_0_6_287 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_358 ();
 DECAPx4_ASAP7_75t_R FILLER_0_6_380 ();
 FILLER_ASAP7_75t_R FILLER_0_6_390 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_414 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_441 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_461 ();
 DECAPx6_ASAP7_75t_R FILLER_0_6_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_485 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_507 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_529 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_551 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_573 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_595 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_617 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_639 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_661 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_683 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_705 ();
 DECAPx10_ASAP7_75t_R FILLER_0_6_727 ();
 DECAPx2_ASAP7_75t_R FILLER_0_6_749 ();
 FILLER_ASAP7_75t_R FILLER_0_6_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_6_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_313 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_349 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_356 ();
 FILLER_ASAP7_75t_R FILLER_0_7_370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_378 ();
 DECAPx1_ASAP7_75t_R FILLER_0_7_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_7_411 ();
 FILLER_ASAP7_75t_R FILLER_0_7_417 ();
 DECAPx6_ASAP7_75t_R FILLER_0_7_440 ();
 FILLER_ASAP7_75t_R FILLER_0_7_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_456 ();
 FILLER_ASAP7_75t_R FILLER_0_7_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_483 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_505 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_527 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_549 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_571 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_593 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_615 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_637 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_659 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_681 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_703 ();
 DECAPx10_ASAP7_75t_R FILLER_0_7_725 ();
 DECAPx4_ASAP7_75t_R FILLER_0_7_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_7_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_266 ();
 FILLER_ASAP7_75t_R FILLER_0_8_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_313 ();
 DECAPx1_ASAP7_75t_R FILLER_0_8_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_382 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_402 ();
 DECAPx6_ASAP7_75t_R FILLER_0_8_423 ();
 FILLER_ASAP7_75t_R FILLER_0_8_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_8_439 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_8_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_8_750 ();
 FILLER_ASAP7_75t_R FILLER_0_8_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_288 ();
 DECAPx4_ASAP7_75t_R FILLER_0_9_310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_9_341 ();
 DECAPx1_ASAP7_75t_R FILLER_0_9_355 ();
 DECAPx4_ASAP7_75t_R FILLER_0_9_362 ();
 FILLER_ASAP7_75t_R FILLER_0_9_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_374 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_471 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_493 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_515 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_537 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_559 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_603 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_647 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_669 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_691 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_713 ();
 DECAPx10_ASAP7_75t_R FILLER_0_9_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_9_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_346 ();
 DECAPx6_ASAP7_75t_R FILLER_0_10_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_383 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_405 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_427 ();
 DECAPx4_ASAP7_75t_R FILLER_0_10_449 ();
 FILLER_ASAP7_75t_R FILLER_0_10_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_487 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_509 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_531 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_553 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_575 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_597 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_641 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_663 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_685 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_707 ();
 DECAPx10_ASAP7_75t_R FILLER_0_10_729 ();
 DECAPx2_ASAP7_75t_R FILLER_0_10_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_10_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_244 ();
 DECAPx4_ASAP7_75t_R FILLER_0_11_266 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_279 ();
 FILLER_ASAP7_75t_R FILLER_0_11_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_287 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_321 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_343 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_365 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_389 ();
 FILLER_ASAP7_75t_R FILLER_0_11_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_405 ();
 DECAPx6_ASAP7_75t_R FILLER_0_11_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_441 ();
 DECAPx2_ASAP7_75t_R FILLER_0_11_448 ();
 DECAPx1_ASAP7_75t_R FILLER_0_11_476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_483 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_505 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_527 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_549 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_571 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_593 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_615 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_637 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_659 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_681 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_703 ();
 DECAPx10_ASAP7_75t_R FILLER_0_11_725 ();
 DECAPx4_ASAP7_75t_R FILLER_0_11_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_11_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_266 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_302 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_309 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_344 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_366 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_378 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_406 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_413 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_435 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_12_468 ();
 FILLER_ASAP7_75t_R FILLER_0_12_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_12_476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_12_718 ();
 DECAPx6_ASAP7_75t_R FILLER_0_12_740 ();
 DECAPx1_ASAP7_75t_R FILLER_0_12_754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_332 ();
 DECAPx4_ASAP7_75t_R FILLER_0_13_362 ();
 FILLER_ASAP7_75t_R FILLER_0_13_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_374 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_13_403 ();
 FILLER_ASAP7_75t_R FILLER_0_13_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_419 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_444 ();
 FILLER_ASAP7_75t_R FILLER_0_13_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_491 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_535 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_579 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_601 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_623 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_645 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_667 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_689 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_711 ();
 DECAPx10_ASAP7_75t_R FILLER_0_13_733 ();
 FILLER_ASAP7_75t_R FILLER_0_13_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_13_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_14_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_330 ();
 DECAPx6_ASAP7_75t_R FILLER_0_14_355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_369 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_399 ();
 DECAPx6_ASAP7_75t_R FILLER_0_14_421 ();
 DECAPx1_ASAP7_75t_R FILLER_0_14_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_439 ();
 DECAPx4_ASAP7_75t_R FILLER_0_14_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_495 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_517 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_539 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_561 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_583 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_605 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_627 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_649 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_671 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_693 ();
 DECAPx10_ASAP7_75t_R FILLER_0_14_715 ();
 DECAPx6_ASAP7_75t_R FILLER_0_14_737 ();
 DECAPx2_ASAP7_75t_R FILLER_0_14_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_14_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_288 ();
 FILLER_ASAP7_75t_R FILLER_0_15_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_334 ();
 DECAPx1_ASAP7_75t_R FILLER_0_15_357 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_364 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_386 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_430 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_452 ();
 DECAPx2_ASAP7_75t_R FILLER_0_15_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_472 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_479 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_501 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_523 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_611 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_633 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_677 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_699 ();
 DECAPx10_ASAP7_75t_R FILLER_0_15_721 ();
 DECAPx6_ASAP7_75t_R FILLER_0_15_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_15_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_16_332 ();
 FILLER_ASAP7_75t_R FILLER_0_16_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_350 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_357 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_379 ();
 FILLER_ASAP7_75t_R FILLER_0_16_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_387 ();
 FILLER_ASAP7_75t_R FILLER_0_16_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_16_396 ();
 DECAPx1_ASAP7_75t_R FILLER_0_16_417 ();
 DECAPx6_ASAP7_75t_R FILLER_0_16_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_16_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_16_750 ();
 FILLER_ASAP7_75t_R FILLER_0_16_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_17_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_330 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_352 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_374 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_396 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_429 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_475 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_497 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_519 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_541 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_563 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_585 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_607 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_629 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_651 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_673 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_695 ();
 DECAPx10_ASAP7_75t_R FILLER_0_17_717 ();
 DECAPx6_ASAP7_75t_R FILLER_0_17_739 ();
 DECAPx1_ASAP7_75t_R FILLER_0_17_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_17_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_18_332 ();
 FILLER_ASAP7_75t_R FILLER_0_18_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_18_344 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_370 ();
 DECAPx6_ASAP7_75t_R FILLER_0_18_392 ();
 FILLER_ASAP7_75t_R FILLER_0_18_406 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_414 ();
 DECAPx1_ASAP7_75t_R FILLER_0_18_436 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_18_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_18_750 ();
 FILLER_ASAP7_75t_R FILLER_0_18_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_287 ();
 DECAPx2_ASAP7_75t_R FILLER_0_19_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_307 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_329 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_19_365 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_19_720 ();
 DECAPx6_ASAP7_75t_R FILLER_0_19_742 ();
 FILLER_ASAP7_75t_R FILLER_0_19_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_332 ();
 DECAPx6_ASAP7_75t_R FILLER_0_20_354 ();
 FILLER_ASAP7_75t_R FILLER_0_20_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_404 ();
 DECAPx6_ASAP7_75t_R FILLER_0_20_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_20_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_477 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_499 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_587 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_609 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_631 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_653 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_675 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_697 ();
 DECAPx10_ASAP7_75t_R FILLER_0_20_719 ();
 DECAPx6_ASAP7_75t_R FILLER_0_20_741 ();
 FILLER_ASAP7_75t_R FILLER_0_20_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_20_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_21_332 ();
 FILLER_ASAP7_75t_R FILLER_0_21_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_340 ();
 FILLER_ASAP7_75t_R FILLER_0_21_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_21_346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_21_720 ();
 DECAPx6_ASAP7_75t_R FILLER_0_21_742 ();
 FILLER_ASAP7_75t_R FILLER_0_21_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_22_310 ();
 FILLER_ASAP7_75t_R FILLER_0_22_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_22_326 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_349 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_371 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_398 ();
 FILLER_ASAP7_75t_R FILLER_0_22_404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_22_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_22_750 ();
 FILLER_ASAP7_75t_R FILLER_0_22_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_23_316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_343 ();
 DECAPx6_ASAP7_75t_R FILLER_0_23_365 ();
 DECAPx1_ASAP7_75t_R FILLER_0_23_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_383 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_405 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_427 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_449 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_471 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_493 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_515 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_537 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_559 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_603 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_647 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_669 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_691 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_713 ();
 DECAPx10_ASAP7_75t_R FILLER_0_23_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_23_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_24_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_336 ();
 DECAPx6_ASAP7_75t_R FILLER_0_24_358 ();
 DECAPx1_ASAP7_75t_R FILLER_0_24_372 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_394 ();
 FILLER_ASAP7_75t_R FILLER_0_24_416 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_24_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_24_750 ();
 FILLER_ASAP7_75t_R FILLER_0_24_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_376 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_433 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_455 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_477 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_499 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_587 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_609 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_631 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_653 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_675 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_697 ();
 DECAPx10_ASAP7_75t_R FILLER_0_25_719 ();
 DECAPx6_ASAP7_75t_R FILLER_0_25_741 ();
 FILLER_ASAP7_75t_R FILLER_0_25_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_25_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_332 ();
 DECAPx1_ASAP7_75t_R FILLER_0_26_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_26_350 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_26_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_26_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_26_750 ();
 FILLER_ASAP7_75t_R FILLER_0_26_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_222 ();
 DECAPx6_ASAP7_75t_R FILLER_0_27_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_324 ();
 FILLER_ASAP7_75t_R FILLER_0_27_346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_351 ();
 DECAPx6_ASAP7_75t_R FILLER_0_27_373 ();
 DECAPx2_ASAP7_75t_R FILLER_0_27_387 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_413 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_435 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_457 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_479 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_501 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_523 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_611 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_633 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_677 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_699 ();
 DECAPx10_ASAP7_75t_R FILLER_0_27_721 ();
 DECAPx6_ASAP7_75t_R FILLER_0_27_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_27_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_222 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_284 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_350 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_372 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_394 ();
 FILLER_ASAP7_75t_R FILLER_0_28_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_402 ();
 DECAPx6_ASAP7_75t_R FILLER_0_28_424 ();
 FILLER_ASAP7_75t_R FILLER_0_28_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_28_440 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_28_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_28_750 ();
 FILLER_ASAP7_75t_R FILLER_0_28_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_29_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_29_346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_412 ();
 DECAPx6_ASAP7_75t_R FILLER_0_29_434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_454 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_29_718 ();
 DECAPx6_ASAP7_75t_R FILLER_0_29_740 ();
 DECAPx1_ASAP7_75t_R FILLER_0_29_754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_354 ();
 DECAPx6_ASAP7_75t_R FILLER_0_30_376 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_390 ();
 FILLER_ASAP7_75t_R FILLER_0_30_402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_407 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_429 ();
 DECAPx4_ASAP7_75t_R FILLER_0_30_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_30_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_30_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_30_750 ();
 FILLER_ASAP7_75t_R FILLER_0_30_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_266 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_302 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_324 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_346 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_368 ();
 FILLER_ASAP7_75t_R FILLER_0_31_390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_413 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_435 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_457 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_479 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_501 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_523 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_611 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_633 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_677 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_699 ();
 DECAPx10_ASAP7_75t_R FILLER_0_31_721 ();
 DECAPx6_ASAP7_75t_R FILLER_0_31_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_31_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_288 ();
 DECAPx1_ASAP7_75t_R FILLER_0_32_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_320 ();
 DECAPx4_ASAP7_75t_R FILLER_0_32_342 ();
 FILLER_ASAP7_75t_R FILLER_0_32_352 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_382 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_32_448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_32_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_32_750 ();
 FILLER_ASAP7_75t_R FILLER_0_32_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_354 ();
 DECAPx4_ASAP7_75t_R FILLER_0_33_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_430 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_452 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_474 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_496 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_518 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_540 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_562 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_584 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_606 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_672 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_694 ();
 DECAPx10_ASAP7_75t_R FILLER_0_33_716 ();
 DECAPx6_ASAP7_75t_R FILLER_0_33_738 ();
 DECAPx2_ASAP7_75t_R FILLER_0_33_752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_288 ();
 DECAPx4_ASAP7_75t_R FILLER_0_34_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_323 ();
 FILLER_ASAP7_75t_R FILLER_0_34_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_347 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_369 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_436 ();
 DECAPx1_ASAP7_75t_R FILLER_0_34_458 ();
 DECAPx4_ASAP7_75t_R FILLER_0_34_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_34_474 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_496 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_518 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_540 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_562 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_584 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_606 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_672 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_694 ();
 DECAPx10_ASAP7_75t_R FILLER_0_34_716 ();
 DECAPx6_ASAP7_75t_R FILLER_0_34_738 ();
 DECAPx2_ASAP7_75t_R FILLER_0_34_752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_354 ();
 DECAPx4_ASAP7_75t_R FILLER_0_35_376 ();
 FILLER_ASAP7_75t_R FILLER_0_35_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_35_388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_35_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_35_750 ();
 FILLER_ASAP7_75t_R FILLER_0_35_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_310 ();
 FILLER_ASAP7_75t_R FILLER_0_36_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_318 ();
 DECAPx6_ASAP7_75t_R FILLER_0_36_341 ();
 FILLER_ASAP7_75t_R FILLER_0_36_377 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_385 ();
 DECAPx6_ASAP7_75t_R FILLER_0_36_407 ();
 FILLER_ASAP7_75t_R FILLER_0_36_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_423 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_427 ();
 DECAPx4_ASAP7_75t_R FILLER_0_36_449 ();
 FILLER_ASAP7_75t_R FILLER_0_36_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_36_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_36_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_36_750 ();
 FILLER_ASAP7_75t_R FILLER_0_36_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_37_332 ();
 FILLER_ASAP7_75t_R FILLER_0_37_341 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_436 ();
 DECAPx4_ASAP7_75t_R FILLER_0_37_458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_489 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_511 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_533 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_555 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_577 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_599 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_621 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_643 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_665 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_687 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_709 ();
 DECAPx10_ASAP7_75t_R FILLER_0_37_731 ();
 DECAPx1_ASAP7_75t_R FILLER_0_37_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_37_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_266 ();
 DECAPx6_ASAP7_75t_R FILLER_0_38_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_308 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_334 ();
 DECAPx4_ASAP7_75t_R FILLER_0_38_356 ();
 FILLER_ASAP7_75t_R FILLER_0_38_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_368 ();
 DECAPx4_ASAP7_75t_R FILLER_0_38_372 ();
 DECAPx6_ASAP7_75t_R FILLER_0_38_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_424 ();
 FILLER_ASAP7_75t_R FILLER_0_38_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_38_448 ();
 DECAPx4_ASAP7_75t_R FILLER_0_38_452 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_38_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_38_750 ();
 FILLER_ASAP7_75t_R FILLER_0_38_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_266 ();
 DECAPx6_ASAP7_75t_R FILLER_0_39_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_302 ();
 DECAPx1_ASAP7_75t_R FILLER_0_39_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_315 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_336 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_358 ();
 DECAPx4_ASAP7_75t_R FILLER_0_39_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_39_381 ();
 FILLER_ASAP7_75t_R FILLER_0_39_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_39_730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_39_752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_266 ();
 DECAPx6_ASAP7_75t_R FILLER_0_40_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_324 ();
 DECAPx1_ASAP7_75t_R FILLER_0_40_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_40_350 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_379 ();
 DECAPx2_ASAP7_75t_R FILLER_0_40_401 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_440 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_550 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_594 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_638 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_704 ();
 DECAPx10_ASAP7_75t_R FILLER_0_40_726 ();
 DECAPx4_ASAP7_75t_R FILLER_0_40_748 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_310 ();
 FILLER_ASAP7_75t_R FILLER_0_41_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_318 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_340 ();
 FILLER_ASAP7_75t_R FILLER_0_41_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_41_355 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_387 ();
 DECAPx4_ASAP7_75t_R FILLER_0_41_409 ();
 FILLER_ASAP7_75t_R FILLER_0_41_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_421 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_450 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_457 ();
 FILLER_ASAP7_75t_R FILLER_0_41_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_473 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_495 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_517 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_539 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_561 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_583 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_605 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_627 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_649 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_671 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_693 ();
 DECAPx10_ASAP7_75t_R FILLER_0_41_715 ();
 DECAPx6_ASAP7_75t_R FILLER_0_41_737 ();
 DECAPx2_ASAP7_75t_R FILLER_0_41_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_41_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_332 ();
 FILLER_ASAP7_75t_R FILLER_0_42_342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_353 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_373 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_377 ();
 DECAPx4_ASAP7_75t_R FILLER_0_42_399 ();
 FILLER_ASAP7_75t_R FILLER_0_42_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_42_411 ();
 DECAPx6_ASAP7_75t_R FILLER_0_42_415 ();
 DECAPx1_ASAP7_75t_R FILLER_0_42_429 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_454 ();
 FILLER_ASAP7_75t_R FILLER_0_42_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_42_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_42_750 ();
 FILLER_ASAP7_75t_R FILLER_0_42_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_43_324 ();
 FILLER_ASAP7_75t_R FILLER_0_43_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_352 ();
 FILLER_ASAP7_75t_R FILLER_0_43_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_358 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_365 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_377 ();
 DECAPx2_ASAP7_75t_R FILLER_0_43_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_405 ();
 DECAPx6_ASAP7_75t_R FILLER_0_43_428 ();
 FILLER_ASAP7_75t_R FILLER_0_43_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_493 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_515 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_537 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_559 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_603 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_647 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_669 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_691 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_713 ();
 DECAPx10_ASAP7_75t_R FILLER_0_43_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_43_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_332 ();
 DECAPx1_ASAP7_75t_R FILLER_0_44_354 ();
 DECAPx6_ASAP7_75t_R FILLER_0_44_380 ();
 FILLER_ASAP7_75t_R FILLER_0_44_394 ();
 DECAPx6_ASAP7_75t_R FILLER_0_44_399 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_413 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_425 ();
 DECAPx6_ASAP7_75t_R FILLER_0_44_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_44_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_44_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_44_750 ();
 FILLER_ASAP7_75t_R FILLER_0_44_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_424 ();
 DECAPx2_ASAP7_75t_R FILLER_0_45_467 ();
 FILLER_ASAP7_75t_R FILLER_0_45_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_475 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_497 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_519 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_541 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_563 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_585 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_607 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_629 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_651 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_673 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_695 ();
 DECAPx10_ASAP7_75t_R FILLER_0_45_717 ();
 DECAPx6_ASAP7_75t_R FILLER_0_45_739 ();
 DECAPx1_ASAP7_75t_R FILLER_0_45_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_45_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_46_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_336 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_365 ();
 FILLER_ASAP7_75t_R FILLER_0_46_371 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_379 ();
 FILLER_ASAP7_75t_R FILLER_0_46_389 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_404 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_425 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_461 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_46_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_46_484 ();
 DECAPx4_ASAP7_75t_R FILLER_0_46_491 ();
 FILLER_ASAP7_75t_R FILLER_0_46_501 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46_722 ();
 DECAPx6_ASAP7_75t_R FILLER_0_46_744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_47_332 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_351 ();
 DECAPx6_ASAP7_75t_R FILLER_0_47_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_47_418 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_482 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_504 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_526 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_548 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_570 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_592 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_614 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_636 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_658 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_680 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_702 ();
 DECAPx10_ASAP7_75t_R FILLER_0_47_724 ();
 DECAPx4_ASAP7_75t_R FILLER_0_47_746 ();
 FILLER_ASAP7_75t_R FILLER_0_47_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_310 ();
 FILLER_ASAP7_75t_R FILLER_0_48_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_359 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_397 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_419 ();
 DECAPx1_ASAP7_75t_R FILLER_0_48_429 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_454 ();
 FILLER_ASAP7_75t_R FILLER_0_48_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_485 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_507 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_529 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_551 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_573 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_595 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_617 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_639 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_661 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_683 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_705 ();
 DECAPx10_ASAP7_75t_R FILLER_0_48_727 ();
 DECAPx2_ASAP7_75t_R FILLER_0_48_749 ();
 FILLER_ASAP7_75t_R FILLER_0_48_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_48_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_354 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_376 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_384 ();
 DECAPx6_ASAP7_75t_R FILLER_0_49_406 ();
 FILLER_ASAP7_75t_R FILLER_0_49_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_445 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_467 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_489 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_511 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_533 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_555 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_577 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_599 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_621 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_643 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_665 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_687 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_709 ();
 DECAPx10_ASAP7_75t_R FILLER_0_49_731 ();
 DECAPx1_ASAP7_75t_R FILLER_0_49_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_49_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_328 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_332 ();
 FILLER_ASAP7_75t_R FILLER_0_50_338 ();
 FILLER_ASAP7_75t_R FILLER_0_50_362 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_385 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_401 ();
 DECAPx2_ASAP7_75t_R FILLER_0_50_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_429 ();
 DECAPx4_ASAP7_75t_R FILLER_0_50_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_461 ();
 FILLER_ASAP7_75t_R FILLER_0_50_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_50_476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_50_718 ();
 DECAPx6_ASAP7_75t_R FILLER_0_50_740 ();
 DECAPx1_ASAP7_75t_R FILLER_0_50_754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_288 ();
 DECAPx4_ASAP7_75t_R FILLER_0_51_310 ();
 FILLER_ASAP7_75t_R FILLER_0_51_320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_344 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_366 ();
 FILLER_ASAP7_75t_R FILLER_0_51_380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_388 ();
 DECAPx4_ASAP7_75t_R FILLER_0_51_410 ();
 FILLER_ASAP7_75t_R FILLER_0_51_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_439 ();
 DECAPx6_ASAP7_75t_R FILLER_0_51_461 ();
 DECAPx2_ASAP7_75t_R FILLER_0_51_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_481 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_503 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_525 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_569 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_591 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_613 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_635 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_657 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_679 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_701 ();
 DECAPx10_ASAP7_75t_R FILLER_0_51_723 ();
 DECAPx4_ASAP7_75t_R FILLER_0_51_745 ();
 FILLER_ASAP7_75t_R FILLER_0_51_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_51_757 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_2 ();
 FILLER_ASAP7_75t_R FILLER_0_52_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_45 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_89 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_111 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_133 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_155 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_177 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_199 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_221 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_243 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_265 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_300 ();
 FILLER_ASAP7_75t_R FILLER_0_52_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_314 ();
 DECAPx2_ASAP7_75t_R FILLER_0_52_336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_352 ();
 DECAPx4_ASAP7_75t_R FILLER_0_52_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_384 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_394 ();
 DECAPx6_ASAP7_75t_R FILLER_0_52_416 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_434 ();
 DECAPx1_ASAP7_75t_R FILLER_0_52_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_52_461 ();
 DECAPx4_ASAP7_75t_R FILLER_0_52_464 ();
 FILLER_ASAP7_75t_R FILLER_0_52_474 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_479 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_501 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_523 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_611 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_633 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_677 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_699 ();
 DECAPx4_ASAP7_75t_R FILLER_0_52_721 ();
 DECAPx10_ASAP7_75t_R FILLER_0_52_736 ();
 DECAPx4_ASAP7_75t_R FILLER_0_53_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_12 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_50 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_72 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_94 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_204 ();
 DECAPx1_ASAP7_75t_R FILLER_0_53_226 ();
 DECAPx4_ASAP7_75t_R FILLER_0_53_251 ();
 FILLER_ASAP7_75t_R FILLER_0_53_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_263 ();
 DECAPx6_ASAP7_75t_R FILLER_0_53_285 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_311 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_348 ();
 FILLER_ASAP7_75t_R FILLER_0_53_354 ();
 FILLER_ASAP7_75t_R FILLER_0_53_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_379 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_386 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_430 ();
 DECAPx2_ASAP7_75t_R FILLER_0_53_452 ();
 FILLER_ASAP7_75t_R FILLER_0_53_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_53_708 ();
 DECAPx4_ASAP7_75t_R FILLER_0_53_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_53_740 ();
 FILLER_ASAP7_75t_R FILLER_0_53_751 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_44 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_88 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_132 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_154 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_176 ();
 DECAPx6_ASAP7_75t_R FILLER_0_54_198 ();
 DECAPx2_ASAP7_75t_R FILLER_0_54_212 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_261 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_287 ();
 FILLER_ASAP7_75t_R FILLER_0_54_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_375 ();
 DECAPx6_ASAP7_75t_R FILLER_0_54_380 ();
 FILLER_ASAP7_75t_R FILLER_0_54_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_428 ();
 DECAPx4_ASAP7_75t_R FILLER_0_54_450 ();
 FILLER_ASAP7_75t_R FILLER_0_54_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_550 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_594 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_638 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_54_704 ();
 DECAPx6_ASAP7_75t_R FILLER_0_54_726 ();
 FILLER_ASAP7_75t_R FILLER_0_54_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_742 ();
 DECAPx1_ASAP7_75t_R FILLER_0_54_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_54_757 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_7 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_35 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_57 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_79 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_145 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_167 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_189 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_211 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_233 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_264 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_278 ();
 FILLER_ASAP7_75t_R FILLER_0_55_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_307 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_329 ();
 FILLER_ASAP7_75t_R FILLER_0_55_339 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_384 ();
 FILLER_ASAP7_75t_R FILLER_0_55_390 ();
 DECAPx6_ASAP7_75t_R FILLER_0_55_407 ();
 FILLER_ASAP7_75t_R FILLER_0_55_421 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_445 ();
 FILLER_ASAP7_75t_R FILLER_0_55_455 ();
 DECAPx4_ASAP7_75t_R FILLER_0_55_460 ();
 FILLER_ASAP7_75t_R FILLER_0_55_470 ();
 FILLER_ASAP7_75t_R FILLER_0_55_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_496 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_55_698 ();
 DECAPx2_ASAP7_75t_R FILLER_0_55_720 ();
 FILLER_ASAP7_75t_R FILLER_0_55_736 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_747 ();
 DECAPx1_ASAP7_75t_R FILLER_0_55_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_55_757 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_48 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_70 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_92 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_246 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_296 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_318 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_346 ();
 DECAPx4_ASAP7_75t_R FILLER_0_56_368 ();
 DECAPx4_ASAP7_75t_R FILLER_0_56_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_394 ();
 DECAPx4_ASAP7_75t_R FILLER_0_56_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_417 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_440 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_464 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_485 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_492 ();
 DECAPx2_ASAP7_75t_R FILLER_0_56_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_56_512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_516 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_560 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_604 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_626 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_648 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_670 ();
 DECAPx10_ASAP7_75t_R FILLER_0_56_692 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_714 ();
 DECAPx1_ASAP7_75t_R FILLER_0_56_728 ();
 DECAPx6_ASAP7_75t_R FILLER_0_56_742 ();
 FILLER_ASAP7_75t_R FILLER_0_56_756 ();
 DECAPx4_ASAP7_75t_R FILLER_0_57_2 ();
 FILLER_ASAP7_75t_R FILLER_0_57_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_51 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_73 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_95 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_139 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_161 ();
 DECAPx4_ASAP7_75t_R FILLER_0_57_183 ();
 FILLER_ASAP7_75t_R FILLER_0_57_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_195 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_273 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_317 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_355 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_403 ();
 DECAPx6_ASAP7_75t_R FILLER_0_57_410 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_428 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_432 ();
 DECAPx4_ASAP7_75t_R FILLER_0_57_454 ();
 FILLER_ASAP7_75t_R FILLER_0_57_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_57_706 ();
 FILLER_ASAP7_75t_R FILLER_0_57_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_730 ();
 DECAPx1_ASAP7_75t_R FILLER_0_57_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_740 ();
 DECAPx2_ASAP7_75t_R FILLER_0_57_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_57_752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_8 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_134 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_191 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_213 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_227 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_254 ();
 FILLER_ASAP7_75t_R FILLER_0_58_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_262 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_284 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_306 ();
 FILLER_ASAP7_75t_R FILLER_0_58_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_318 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_361 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_373 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_387 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_413 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_431 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_439 ();
 DECAPx6_ASAP7_75t_R FILLER_0_58_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_482 ();
 DECAPx2_ASAP7_75t_R FILLER_0_58_486 ();
 FILLER_ASAP7_75t_R FILLER_0_58_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_516 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_569 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_591 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_613 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_635 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_657 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_679 ();
 DECAPx10_ASAP7_75t_R FILLER_0_58_701 ();
 DECAPx4_ASAP7_75t_R FILLER_0_58_723 ();
 FILLER_ASAP7_75t_R FILLER_0_58_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_735 ();
 DECAPx1_ASAP7_75t_R FILLER_0_58_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_58_750 ();
 FILLER_ASAP7_75t_R FILLER_0_58_756 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_12 ();
 FILLER_ASAP7_75t_R FILLER_0_59_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_53 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_75 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_97 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_119 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_141 ();
 DECAPx6_ASAP7_75t_R FILLER_0_59_163 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_177 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_204 ();
 FILLER_ASAP7_75t_R FILLER_0_59_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_250 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_325 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_353 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_385 ();
 DECAPx6_ASAP7_75t_R FILLER_0_59_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_421 ();
 DECAPx6_ASAP7_75t_R FILLER_0_59_428 ();
 DECAPx2_ASAP7_75t_R FILLER_0_59_442 ();
 DECAPx1_ASAP7_75t_R FILLER_0_59_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_474 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_59_698 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_720 ();
 FILLER_ASAP7_75t_R FILLER_0_59_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_59_732 ();
 DECAPx4_ASAP7_75t_R FILLER_0_59_748 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_12 ();
 FILLER_ASAP7_75t_R FILLER_0_60_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_51 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_73 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_95 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_139 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_161 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_186 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_208 ();
 FILLER_ASAP7_75t_R FILLER_0_60_214 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_237 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_259 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_303 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_325 ();
 FILLER_ASAP7_75t_R FILLER_0_60_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_359 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_381 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_395 ();
 DECAPx1_ASAP7_75t_R FILLER_0_60_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_415 ();
 FILLER_ASAP7_75t_R FILLER_0_60_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_424 ();
 DECAPx4_ASAP7_75t_R FILLER_0_60_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_438 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_456 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_478 ();
 FILLER_ASAP7_75t_R FILLER_0_60_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_503 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_507 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_549 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_571 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_593 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_615 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_637 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_659 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_681 ();
 DECAPx10_ASAP7_75t_R FILLER_0_60_703 ();
 DECAPx6_ASAP7_75t_R FILLER_0_60_725 ();
 FILLER_ASAP7_75t_R FILLER_0_60_739 ();
 DECAPx2_ASAP7_75t_R FILLER_0_60_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_60_752 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_49 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_71 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_93 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_115 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_137 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_159 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_181 ();
 DECAPx6_ASAP7_75t_R FILLER_0_61_203 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_242 ();
 FILLER_ASAP7_75t_R FILLER_0_61_264 ();
 DECAPx6_ASAP7_75t_R FILLER_0_61_287 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_307 ();
 FILLER_ASAP7_75t_R FILLER_0_61_329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_61_358 ();
 FILLER_ASAP7_75t_R FILLER_0_61_364 ();
 DECAPx6_ASAP7_75t_R FILLER_0_61_370 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_446 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_497 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_504 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_517 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_551 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_573 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_595 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_617 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_639 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_661 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_683 ();
 DECAPx10_ASAP7_75t_R FILLER_0_61_705 ();
 DECAPx4_ASAP7_75t_R FILLER_0_61_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_737 ();
 DECAPx1_ASAP7_75t_R FILLER_0_61_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_61_757 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_2 ();
 FILLER_ASAP7_75t_R FILLER_0_62_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_50 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_72 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_94 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_138 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_170 ();
 DECAPx2_ASAP7_75t_R FILLER_0_62_213 ();
 FILLER_ASAP7_75t_R FILLER_0_62_219 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_268 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_290 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_334 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_372 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_398 ();
 DECAPx4_ASAP7_75t_R FILLER_0_62_402 ();
 FILLER_ASAP7_75t_R FILLER_0_62_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_437 ();
 FILLER_ASAP7_75t_R FILLER_0_62_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_461 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_482 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_62_684 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_720 ();
 DECAPx1_ASAP7_75t_R FILLER_0_62_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_735 ();
 DECAPx6_ASAP7_75t_R FILLER_0_62_741 ();
 FILLER_ASAP7_75t_R FILLER_0_62_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_62_757 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_11 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_44 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_88 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_132 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_154 ();
 DECAPx4_ASAP7_75t_R FILLER_0_63_176 ();
 FILLER_ASAP7_75t_R FILLER_0_63_186 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_209 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_231 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_253 ();
 FILLER_ASAP7_75t_R FILLER_0_63_259 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_304 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_326 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_363 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_386 ();
 DECAPx6_ASAP7_75t_R FILLER_0_63_408 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_428 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_435 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_457 ();
 DECAPx1_ASAP7_75t_R FILLER_0_63_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_483 ();
 FILLER_ASAP7_75t_R FILLER_0_63_506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_511 ();
 DECAPx4_ASAP7_75t_R FILLER_0_63_533 ();
 FILLER_ASAP7_75t_R FILLER_0_63_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_63_545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_571 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_593 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_615 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_637 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_659 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_681 ();
 DECAPx10_ASAP7_75t_R FILLER_0_63_703 ();
 FILLER_ASAP7_75t_R FILLER_0_63_725 ();
 DECAPx4_ASAP7_75t_R FILLER_0_63_732 ();
 DECAPx2_ASAP7_75t_R FILLER_0_63_752 ();
 DECAPx4_ASAP7_75t_R FILLER_0_64_2 ();
 FILLER_ASAP7_75t_R FILLER_0_64_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_51 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_73 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_95 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_139 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_161 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_189 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_211 ();
 DECAPx1_ASAP7_75t_R FILLER_0_64_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_251 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_273 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_293 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_315 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_337 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_359 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_373 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_407 ();
 FILLER_ASAP7_75t_R FILLER_0_64_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_415 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_422 ();
 DECAPx2_ASAP7_75t_R FILLER_0_64_431 ();
 FILLER_ASAP7_75t_R FILLER_0_64_437 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_439 ();
 DECAPx4_ASAP7_75t_R FILLER_0_64_446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_508 ();
 FILLER_ASAP7_75t_R FILLER_0_64_530 ();
 DECAPx6_ASAP7_75t_R FILLER_0_64_554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_571 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_593 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_615 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_637 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_659 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_681 ();
 DECAPx10_ASAP7_75t_R FILLER_0_64_703 ();
 FILLER_ASAP7_75t_R FILLER_0_64_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_64_727 ();
 DECAPx4_ASAP7_75t_R FILLER_0_64_733 ();
 DECAPx4_ASAP7_75t_R FILLER_0_64_748 ();
 DECAPx4_ASAP7_75t_R FILLER_0_65_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_17 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_35 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_57 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_79 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_145 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_167 ();
 FILLER_ASAP7_75t_R FILLER_0_65_173 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_196 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_266 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_280 ();
 FILLER_ASAP7_75t_R FILLER_0_65_307 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_331 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_353 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_375 ();
 FILLER_ASAP7_75t_R FILLER_0_65_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_391 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_398 ();
 DECAPx2_ASAP7_75t_R FILLER_0_65_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_418 ();
 FILLER_ASAP7_75t_R FILLER_0_65_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_449 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_459 ();
 DECAPx4_ASAP7_75t_R FILLER_0_65_481 ();
 FILLER_ASAP7_75t_R FILLER_0_65_491 ();
 DECAPx6_ASAP7_75t_R FILLER_0_65_518 ();
 DECAPx1_ASAP7_75t_R FILLER_0_65_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_562 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_584 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_606 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_672 ();
 DECAPx10_ASAP7_75t_R FILLER_0_65_694 ();
 DECAPx4_ASAP7_75t_R FILLER_0_65_716 ();
 FILLER_ASAP7_75t_R FILLER_0_65_726 ();
 DECAPx4_ASAP7_75t_R FILLER_0_65_733 ();
 FILLER_ASAP7_75t_R FILLER_0_65_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_65_745 ();
 FILLER_ASAP7_75t_R FILLER_0_65_756 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_7 ();
 FILLER_ASAP7_75t_R FILLER_0_66_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_51 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_73 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_95 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_139 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_161 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_183 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_203 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_225 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_247 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_269 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_291 ();
 DECAPx1_ASAP7_75t_R FILLER_0_66_305 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_312 ();
 FILLER_ASAP7_75t_R FILLER_0_66_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_341 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_369 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_401 ();
 DECAPx6_ASAP7_75t_R FILLER_0_66_430 ();
 FILLER_ASAP7_75t_R FILLER_0_66_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_452 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_486 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_561 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_66_700 ();
 DECAPx2_ASAP7_75t_R FILLER_0_66_722 ();
 FILLER_ASAP7_75t_R FILLER_0_66_728 ();
 DECAPx4_ASAP7_75t_R FILLER_0_66_735 ();
 FILLER_ASAP7_75t_R FILLER_0_66_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_66_747 ();
 DECAPx6_ASAP7_75t_R FILLER_0_67_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_67_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_53 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_75 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_97 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_119 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_141 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_163 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_293 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_315 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_359 ();
 DECAPx6_ASAP7_75t_R FILLER_0_67_381 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_395 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_404 ();
 DECAPx6_ASAP7_75t_R FILLER_0_67_416 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_430 ();
 DECAPx4_ASAP7_75t_R FILLER_0_67_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_474 ();
 DECAPx4_ASAP7_75t_R FILLER_0_67_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_513 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_67_700 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_722 ();
 FILLER_ASAP7_75t_R FILLER_0_67_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_67_741 ();
 FILLER_ASAP7_75t_R FILLER_0_67_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_749 ();
 FILLER_ASAP7_75t_R FILLER_0_67_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_67_757 ();
 DECAPx4_ASAP7_75t_R FILLER_0_68_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_45 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_67 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_89 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_111 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_133 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_155 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_177 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_199 ();
 FILLER_ASAP7_75t_R FILLER_0_68_221 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_266 ();
 DECAPx6_ASAP7_75t_R FILLER_0_68_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_308 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_330 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_358 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_387 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_394 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_429 ();
 DECAPx4_ASAP7_75t_R FILLER_0_68_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_461 ();
 FILLER_ASAP7_75t_R FILLER_0_68_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_466 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_473 ();
 FILLER_ASAP7_75t_R FILLER_0_68_501 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_506 ();
 FILLER_ASAP7_75t_R FILLER_0_68_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_530 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_553 ();
 FILLER_ASAP7_75t_R FILLER_0_68_559 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68_696 ();
 DECAPx4_ASAP7_75t_R FILLER_0_68_718 ();
 FILLER_ASAP7_75t_R FILLER_0_68_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_730 ();
 DECAPx1_ASAP7_75t_R FILLER_0_68_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_740 ();
 DECAPx2_ASAP7_75t_R FILLER_0_68_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_68_757 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_6 ();
 FILLER_ASAP7_75t_R FILLER_0_69_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_51 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_73 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_95 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_139 ();
 DECAPx6_ASAP7_75t_R FILLER_0_69_161 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_175 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_200 ();
 DECAPx6_ASAP7_75t_R FILLER_0_69_222 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_236 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_305 ();
 DECAPx6_ASAP7_75t_R FILLER_0_69_327 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_341 ();
 DECAPx6_ASAP7_75t_R FILLER_0_69_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_380 ();
 DECAPx4_ASAP7_75t_R FILLER_0_69_409 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_428 ();
 DECAPx6_ASAP7_75t_R FILLER_0_69_449 ();
 FILLER_ASAP7_75t_R FILLER_0_69_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_465 ();
 FILLER_ASAP7_75t_R FILLER_0_69_478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_501 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_523 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_611 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_633 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_677 ();
 DECAPx10_ASAP7_75t_R FILLER_0_69_699 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_721 ();
 FILLER_ASAP7_75t_R FILLER_0_69_727 ();
 DECAPx2_ASAP7_75t_R FILLER_0_69_732 ();
 DECAPx1_ASAP7_75t_R FILLER_0_69_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_69_747 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_47 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_69 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_91 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_113 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_135 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_157 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_179 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_201 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_223 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_245 ();
 DECAPx6_ASAP7_75t_R FILLER_0_70_267 ();
 FILLER_ASAP7_75t_R FILLER_0_70_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_283 ();
 DECAPx4_ASAP7_75t_R FILLER_0_70_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_315 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_337 ();
 DECAPx6_ASAP7_75t_R FILLER_0_70_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_373 ();
 DECAPx4_ASAP7_75t_R FILLER_0_70_401 ();
 FILLER_ASAP7_75t_R FILLER_0_70_411 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_512 ();
 FILLER_ASAP7_75t_R FILLER_0_70_518 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_541 ();
 FILLER_ASAP7_75t_R FILLER_0_70_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_549 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_571 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_593 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_615 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_637 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_659 ();
 DECAPx10_ASAP7_75t_R FILLER_0_70_681 ();
 DECAPx4_ASAP7_75t_R FILLER_0_70_703 ();
 FILLER_ASAP7_75t_R FILLER_0_70_713 ();
 DECAPx2_ASAP7_75t_R FILLER_0_70_718 ();
 FILLER_ASAP7_75t_R FILLER_0_70_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_726 ();
 FILLER_ASAP7_75t_R FILLER_0_70_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_736 ();
 FILLER_ASAP7_75t_R FILLER_0_70_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_70_752 ();
 FILLER_ASAP7_75t_R FILLER_0_71_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_4 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_47 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_69 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_91 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_113 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_135 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_157 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_179 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_201 ();
 DECAPx6_ASAP7_75t_R FILLER_0_71_223 ();
 FILLER_ASAP7_75t_R FILLER_0_71_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_261 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_283 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_309 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_359 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_403 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_425 ();
 FILLER_ASAP7_75t_R FILLER_0_71_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_433 ();
 DECAPx6_ASAP7_75t_R FILLER_0_71_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_468 ();
 DECAPx6_ASAP7_75t_R FILLER_0_71_490 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_71_706 ();
 DECAPx2_ASAP7_75t_R FILLER_0_71_728 ();
 FILLER_ASAP7_75t_R FILLER_0_71_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_736 ();
 FILLER_ASAP7_75t_R FILLER_0_71_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_742 ();
 DECAPx1_ASAP7_75t_R FILLER_0_71_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_71_752 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_7 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_53 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_75 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_97 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_119 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_141 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_163 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_185 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_207 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_229 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_251 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_273 ();
 DECAPx4_ASAP7_75t_R FILLER_0_72_295 ();
 FILLER_ASAP7_75t_R FILLER_0_72_305 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_349 ();
 DECAPx1_ASAP7_75t_R FILLER_0_72_371 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_423 ();
 DECAPx4_ASAP7_75t_R FILLER_0_72_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_461 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_490 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_512 ();
 DECAPx6_ASAP7_75t_R FILLER_0_72_539 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_559 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_603 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_647 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_669 ();
 DECAPx10_ASAP7_75t_R FILLER_0_72_691 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_713 ();
 DECAPx2_ASAP7_75t_R FILLER_0_72_722 ();
 FILLER_ASAP7_75t_R FILLER_0_72_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_72_742 ();
 FILLER_ASAP7_75t_R FILLER_0_72_746 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_6 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_16 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_44 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_88 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_132 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_154 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_176 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_198 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_220 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_242 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_264 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_286 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_308 ();
 DECAPx2_ASAP7_75t_R FILLER_0_73_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_336 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_358 ();
 DECAPx4_ASAP7_75t_R FILLER_0_73_380 ();
 FILLER_ASAP7_75t_R FILLER_0_73_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_392 ();
 FILLER_ASAP7_75t_R FILLER_0_73_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_422 ();
 DECAPx6_ASAP7_75t_R FILLER_0_73_450 ();
 FILLER_ASAP7_75t_R FILLER_0_73_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_493 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_515 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_537 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_559 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_603 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_647 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_669 ();
 DECAPx10_ASAP7_75t_R FILLER_0_73_691 ();
 DECAPx4_ASAP7_75t_R FILLER_0_73_713 ();
 FILLER_ASAP7_75t_R FILLER_0_73_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_73_725 ();
 DECAPx1_ASAP7_75t_R FILLER_0_73_729 ();
 FILLER_ASAP7_75t_R FILLER_0_73_741 ();
 FILLER_ASAP7_75t_R FILLER_0_73_751 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_7 ();
 FILLER_ASAP7_75t_R FILLER_0_74_21 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_23 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_51 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_73 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_95 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_139 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_161 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_183 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_205 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_227 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_249 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_271 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_293 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_315 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_337 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_381 ();
 DECAPx6_ASAP7_75t_R FILLER_0_74_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_417 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_587 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_609 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_631 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_653 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_675 ();
 DECAPx10_ASAP7_75t_R FILLER_0_74_697 ();
 DECAPx4_ASAP7_75t_R FILLER_0_74_719 ();
 FILLER_ASAP7_75t_R FILLER_0_74_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_734 ();
 DECAPx1_ASAP7_75t_R FILLER_0_74_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_74_747 ();
 DECAPx4_ASAP7_75t_R FILLER_0_75_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_50 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_72 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_94 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_182 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_226 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_248 ();
 FILLER_ASAP7_75t_R FILLER_0_75_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_279 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_301 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_336 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_358 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_378 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_391 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_416 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_438 ();
 FILLER_ASAP7_75t_R FILLER_0_75_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_465 ();
 DECAPx6_ASAP7_75t_R FILLER_0_75_472 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_558 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_580 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_602 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_624 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_646 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_668 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_75_712 ();
 DECAPx2_ASAP7_75t_R FILLER_0_75_734 ();
 DECAPx1_ASAP7_75t_R FILLER_0_75_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_75_757 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_50 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_72 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_94 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_160 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_182 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_218 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_222 ();
 FILLER_ASAP7_75t_R FILLER_0_76_239 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_266 ();
 FILLER_ASAP7_75t_R FILLER_0_76_280 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_324 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_344 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_366 ();
 FILLER_ASAP7_75t_R FILLER_0_76_372 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_417 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_464 ();
 DECAPx1_ASAP7_75t_R FILLER_0_76_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_496 ();
 DECAPx2_ASAP7_75t_R FILLER_0_76_518 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_567 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_589 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_611 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_633 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_655 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_677 ();
 DECAPx10_ASAP7_75t_R FILLER_0_76_699 ();
 DECAPx6_ASAP7_75t_R FILLER_0_76_721 ();
 FILLER_ASAP7_75t_R FILLER_0_76_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_76_737 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_6 ();
 DECAPx6_ASAP7_75t_R FILLER_0_77_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_32 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_54 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_76 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_98 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_120 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_142 ();
 DECAPx4_ASAP7_75t_R FILLER_0_77_164 ();
 FILLER_ASAP7_75t_R FILLER_0_77_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_199 ();
 DECAPx6_ASAP7_75t_R FILLER_0_77_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_283 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_290 ();
 DECAPx4_ASAP7_75t_R FILLER_0_77_308 ();
 FILLER_ASAP7_75t_R FILLER_0_77_318 ();
 DECAPx2_ASAP7_75t_R FILLER_0_77_323 ();
 FILLER_ASAP7_75t_R FILLER_0_77_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_331 ();
 DECAPx4_ASAP7_75t_R FILLER_0_77_353 ();
 FILLER_ASAP7_75t_R FILLER_0_77_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_365 ();
 FILLER_ASAP7_75t_R FILLER_0_77_414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_437 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_459 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_481 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_503 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_525 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_569 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_591 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_613 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_635 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_657 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_679 ();
 DECAPx10_ASAP7_75t_R FILLER_0_77_701 ();
 DECAPx6_ASAP7_75t_R FILLER_0_77_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_737 ();
 DECAPx1_ASAP7_75t_R FILLER_0_77_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_77_757 ();
 DECAPx1_ASAP7_75t_R FILLER_0_78_7 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_11 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_50 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_72 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_94 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_138 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_160 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_174 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_197 ();
 FILLER_ASAP7_75t_R FILLER_0_78_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_203 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_207 ();
 FILLER_ASAP7_75t_R FILLER_0_78_221 ();
 DECAPx4_ASAP7_75t_R FILLER_0_78_245 ();
 FILLER_ASAP7_75t_R FILLER_0_78_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_257 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_261 ();
 FILLER_ASAP7_75t_R FILLER_0_78_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_311 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_340 ();
 FILLER_ASAP7_75t_R FILLER_0_78_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_356 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_363 ();
 DECAPx2_ASAP7_75t_R FILLER_0_78_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_391 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_418 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_440 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_78_706 ();
 DECAPx6_ASAP7_75t_R FILLER_0_78_728 ();
 FILLER_ASAP7_75t_R FILLER_0_78_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_744 ();
 FILLER_ASAP7_75t_R FILLER_0_78_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_78_752 ();
 DECAPx4_ASAP7_75t_R FILLER_0_79_2 ();
 FILLER_ASAP7_75t_R FILLER_0_79_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_47 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_69 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_91 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_113 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_135 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_157 ();
 DECAPx6_ASAP7_75t_R FILLER_0_79_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_218 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_222 ();
 FILLER_ASAP7_75t_R FILLER_0_79_228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_252 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_296 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_318 ();
 DECAPx1_ASAP7_75t_R FILLER_0_79_340 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_350 ();
 DECAPx4_ASAP7_75t_R FILLER_0_79_362 ();
 FILLER_ASAP7_75t_R FILLER_0_79_372 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_395 ();
 DECAPx4_ASAP7_75t_R FILLER_0_79_417 ();
 FILLER_ASAP7_75t_R FILLER_0_79_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_429 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_472 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_494 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_516 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_560 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_604 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_626 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_648 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_670 ();
 DECAPx10_ASAP7_75t_R FILLER_0_79_692 ();
 DECAPx6_ASAP7_75t_R FILLER_0_79_714 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_79_739 ();
 FILLER_ASAP7_75t_R FILLER_0_79_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_79_752 ();
 FILLER_ASAP7_75t_R FILLER_0_80_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_4 ();
 DECAPx6_ASAP7_75t_R FILLER_0_80_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_35 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_57 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_79 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_145 ();
 DECAPx6_ASAP7_75t_R FILLER_0_80_167 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_181 ();
 DECAPx4_ASAP7_75t_R FILLER_0_80_207 ();
 FILLER_ASAP7_75t_R FILLER_0_80_217 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_241 ();
 DECAPx6_ASAP7_75t_R FILLER_0_80_263 ();
 FILLER_ASAP7_75t_R FILLER_0_80_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_80_279 ();
 DECAPx1_ASAP7_75t_R FILLER_0_80_311 ();
 FILLER_ASAP7_75t_R FILLER_0_80_342 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_390 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_684 ();
 DECAPx6_ASAP7_75t_R FILLER_0_80_706 ();
 DECAPx2_ASAP7_75t_R FILLER_0_80_720 ();
 DECAPx10_ASAP7_75t_R FILLER_0_80_736 ();
 FILLER_ASAP7_75t_R FILLER_0_81_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_9 ();
 FILLER_ASAP7_75t_R FILLER_0_81_15 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_44 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_66 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_88 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_110 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_132 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_154 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_176 ();
 DECAPx6_ASAP7_75t_R FILLER_0_81_198 ();
 FILLER_ASAP7_75t_R FILLER_0_81_212 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_220 ();
 FILLER_ASAP7_75t_R FILLER_0_81_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_228 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_251 ();
 FILLER_ASAP7_75t_R FILLER_0_81_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_259 ();
 DECAPx4_ASAP7_75t_R FILLER_0_81_285 ();
 FILLER_ASAP7_75t_R FILLER_0_81_295 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_303 ();
 FILLER_ASAP7_75t_R FILLER_0_81_309 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_323 ();
 FILLER_ASAP7_75t_R FILLER_0_81_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_332 ();
 DECAPx6_ASAP7_75t_R FILLER_0_81_354 ();
 FILLER_ASAP7_75t_R FILLER_0_81_368 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_81_706 ();
 DECAPx4_ASAP7_75t_R FILLER_0_81_728 ();
 FILLER_ASAP7_75t_R FILLER_0_81_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_740 ();
 DECAPx2_ASAP7_75t_R FILLER_0_81_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_81_757 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_2 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_25 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_53 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_75 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_97 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_119 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_141 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_163 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_185 ();
 FILLER_ASAP7_75t_R FILLER_0_82_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_201 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_231 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_235 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_273 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_335 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_353 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_375 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_397 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_419 ();
 DECAPx6_ASAP7_75t_R FILLER_0_82_441 ();
 DECAPx2_ASAP7_75t_R FILLER_0_82_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_82_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_82_708 ();
 DECAPx4_ASAP7_75t_R FILLER_0_82_730 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_745 ();
 DECAPx1_ASAP7_75t_R FILLER_0_82_754 ();
 DECAPx4_ASAP7_75t_R FILLER_0_83_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_40 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_62 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_84 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_106 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_128 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_150 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_172 ();
 FILLER_ASAP7_75t_R FILLER_0_83_194 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_199 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_227 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_272 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_294 ();
 FILLER_ASAP7_75t_R FILLER_0_83_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_339 ();
 FILLER_ASAP7_75t_R FILLER_0_83_345 ();
 DECAPx6_ASAP7_75t_R FILLER_0_83_359 ();
 FILLER_ASAP7_75t_R FILLER_0_83_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_375 ();
 FILLER_ASAP7_75t_R FILLER_0_83_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_384 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_83_412 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_434 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_500 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_698 ();
 DECAPx10_ASAP7_75t_R FILLER_0_83_720 ();
 DECAPx2_ASAP7_75t_R FILLER_0_83_742 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_17 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_50 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_72 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_94 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_116 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_138 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_160 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_186 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_190 ();
 FILLER_ASAP7_75t_R FILLER_0_84_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_198 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_225 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_233 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_247 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_276 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_312 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_341 ();
 DECAPx2_ASAP7_75t_R FILLER_0_84_363 ();
 FILLER_ASAP7_75t_R FILLER_0_84_369 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_377 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_393 ();
 DECAPx1_ASAP7_75t_R FILLER_0_84_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_419 ();
 DECAPx6_ASAP7_75t_R FILLER_0_84_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_478 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_587 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_609 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_631 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_653 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_675 ();
 DECAPx10_ASAP7_75t_R FILLER_0_84_697 ();
 DECAPx6_ASAP7_75t_R FILLER_0_84_719 ();
 FILLER_ASAP7_75t_R FILLER_0_84_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_84_735 ();
 DECAPx4_ASAP7_75t_R FILLER_0_84_746 ();
 FILLER_ASAP7_75t_R FILLER_0_84_756 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_6 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_12 ();
 DECAPx4_ASAP7_75t_R FILLER_0_85_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_33 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_55 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_77 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_99 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_121 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_143 ();
 DECAPx1_ASAP7_75t_R FILLER_0_85_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_169 ();
 FILLER_ASAP7_75t_R FILLER_0_85_192 ();
 DECAPx6_ASAP7_75t_R FILLER_0_85_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_211 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_256 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_278 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_300 ();
 FILLER_ASAP7_75t_R FILLER_0_85_306 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_351 ();
 DECAPx6_ASAP7_75t_R FILLER_0_85_373 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_430 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_452 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_474 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_496 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_518 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_540 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_562 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_584 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_606 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_672 ();
 DECAPx10_ASAP7_75t_R FILLER_0_85_694 ();
 DECAPx4_ASAP7_75t_R FILLER_0_85_716 ();
 FILLER_ASAP7_75t_R FILLER_0_85_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_733 ();
 FILLER_ASAP7_75t_R FILLER_0_85_744 ();
 DECAPx2_ASAP7_75t_R FILLER_0_85_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_85_757 ();
 DECAPx6_ASAP7_75t_R FILLER_0_86_2 ();
 FILLER_ASAP7_75t_R FILLER_0_86_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_33 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_55 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_77 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_99 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_121 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_143 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_165 ();
 FILLER_ASAP7_75t_R FILLER_0_86_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_173 ();
 FILLER_ASAP7_75t_R FILLER_0_86_177 ();
 DECAPx6_ASAP7_75t_R FILLER_0_86_182 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_218 ();
 FILLER_ASAP7_75t_R FILLER_0_86_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_252 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_262 ();
 FILLER_ASAP7_75t_R FILLER_0_86_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_287 ();
 DECAPx6_ASAP7_75t_R FILLER_0_86_313 ();
 FILLER_ASAP7_75t_R FILLER_0_86_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_329 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_336 ();
 FILLER_ASAP7_75t_R FILLER_0_86_342 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_360 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_367 ();
 FILLER_ASAP7_75t_R FILLER_0_86_373 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_381 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_403 ();
 DECAPx6_ASAP7_75t_R FILLER_0_86_425 ();
 FILLER_ASAP7_75t_R FILLER_0_86_439 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_464 ();
 FILLER_ASAP7_75t_R FILLER_0_86_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_498 ();
 FILLER_ASAP7_75t_R FILLER_0_86_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_522 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_544 ();
 FILLER_ASAP7_75t_R FILLER_0_86_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_86_700 ();
 DECAPx4_ASAP7_75t_R FILLER_0_86_722 ();
 FILLER_ASAP7_75t_R FILLER_0_86_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_86_734 ();
 DECAPx2_ASAP7_75t_R FILLER_0_86_740 ();
 FILLER_ASAP7_75t_R FILLER_0_86_746 ();
 DECAPx1_ASAP7_75t_R FILLER_0_87_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_6 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_51 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_73 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_95 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_139 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_161 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_183 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_205 ();
 FILLER_ASAP7_75t_R FILLER_0_87_211 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_260 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_282 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_304 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_348 ();
 DECAPx4_ASAP7_75t_R FILLER_0_87_355 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_371 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_393 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_415 ();
 DECAPx6_ASAP7_75t_R FILLER_0_87_437 ();
 FILLER_ASAP7_75t_R FILLER_0_87_451 ();
 DECAPx6_ASAP7_75t_R FILLER_0_87_483 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_497 ();
 DECAPx6_ASAP7_75t_R FILLER_0_87_524 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_87_544 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_87_698 ();
 DECAPx2_ASAP7_75t_R FILLER_0_87_720 ();
 DECAPx4_ASAP7_75t_R FILLER_0_87_736 ();
 FILLER_ASAP7_75t_R FILLER_0_87_746 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_2 ();
 FILLER_ASAP7_75t_R FILLER_0_88_8 ();
 DECAPx6_ASAP7_75t_R FILLER_0_88_20 ();
 FILLER_ASAP7_75t_R FILLER_0_88_34 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_41 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_63 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_85 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_107 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_129 ();
 DECAPx6_ASAP7_75t_R FILLER_0_88_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_165 ();
 DECAPx6_ASAP7_75t_R FILLER_0_88_194 ();
 FILLER_ASAP7_75t_R FILLER_0_88_208 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_257 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_279 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_301 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_323 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_351 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_361 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_373 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_395 ();
 FILLER_ASAP7_75t_R FILLER_0_88_401 ();
 DECAPx1_ASAP7_75t_R FILLER_0_88_409 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_434 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_486 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_518 ();
 DECAPx6_ASAP7_75t_R FILLER_0_88_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_88_554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_88_708 ();
 DECAPx2_ASAP7_75t_R FILLER_0_88_730 ();
 FILLER_ASAP7_75t_R FILLER_0_88_736 ();
 DECAPx4_ASAP7_75t_R FILLER_0_88_743 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_6 ();
 DECAPx4_ASAP7_75t_R FILLER_0_89_12 ();
 FILLER_ASAP7_75t_R FILLER_0_89_22 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_29 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_51 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_73 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_95 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_117 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_139 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_161 ();
 DECAPx4_ASAP7_75t_R FILLER_0_89_183 ();
 FILLER_ASAP7_75t_R FILLER_0_89_193 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_198 ();
 FILLER_ASAP7_75t_R FILLER_0_89_204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_228 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_250 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_265 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_283 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_336 ();
 FILLER_ASAP7_75t_R FILLER_0_89_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_342 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_375 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_393 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_415 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_437 ();
 FILLER_ASAP7_75t_R FILLER_0_89_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_475 ();
 DECAPx6_ASAP7_75t_R FILLER_0_89_497 ();
 FILLER_ASAP7_75t_R FILLER_0_89_511 ();
 DECAPx4_ASAP7_75t_R FILLER_0_89_534 ();
 FILLER_ASAP7_75t_R FILLER_0_89_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_89_700 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_728 ();
 DECAPx1_ASAP7_75t_R FILLER_0_89_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_738 ();
 DECAPx2_ASAP7_75t_R FILLER_0_89_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_89_750 ();
 FILLER_ASAP7_75t_R FILLER_0_89_756 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_7 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_22 ();
 FILLER_ASAP7_75t_R FILLER_0_90_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_35 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_57 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_79 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_123 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_145 ();
 FILLER_ASAP7_75t_R FILLER_0_90_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_161 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_165 ();
 FILLER_ASAP7_75t_R FILLER_0_90_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_181 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_204 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_226 ();
 DECAPx2_ASAP7_75t_R FILLER_0_90_248 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_276 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_290 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_341 ();
 FILLER_ASAP7_75t_R FILLER_0_90_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_359 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_370 ();
 FILLER_ASAP7_75t_R FILLER_0_90_392 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_400 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_424 ();
 DECAPx6_ASAP7_75t_R FILLER_0_90_446 ();
 FILLER_ASAP7_75t_R FILLER_0_90_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_555 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_577 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_599 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_621 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_643 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_665 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_687 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90_709 ();
 DECAPx4_ASAP7_75t_R FILLER_0_90_731 ();
 FILLER_ASAP7_75t_R FILLER_0_90_741 ();
 DECAPx1_ASAP7_75t_R FILLER_0_90_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_90_757 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_7 ();
 FILLER_ASAP7_75t_R FILLER_0_91_17 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_19 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_25 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_31 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_37 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_59 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_81 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_103 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_125 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_147 ();
 DECAPx1_ASAP7_75t_R FILLER_0_91_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_173 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_177 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_199 ();
 DECAPx6_ASAP7_75t_R FILLER_0_91_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_245 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_274 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_296 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_318 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_340 ();
 FILLER_ASAP7_75t_R FILLER_0_91_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_358 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_365 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_377 ();
 FILLER_ASAP7_75t_R FILLER_0_91_383 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_416 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_438 ();
 FILLER_ASAP7_75t_R FILLER_0_91_448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_513 ();
 DECAPx4_ASAP7_75t_R FILLER_0_91_535 ();
 FILLER_ASAP7_75t_R FILLER_0_91_545 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_91_678 ();
 DECAPx6_ASAP7_75t_R FILLER_0_91_700 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_714 ();
 FILLER_ASAP7_75t_R FILLER_0_91_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_727 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_733 ();
 FILLER_ASAP7_75t_R FILLER_0_91_739 ();
 DECAPx2_ASAP7_75t_R FILLER_0_91_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_91_757 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_7 ();
 FILLER_ASAP7_75t_R FILLER_0_92_13 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_20 ();
 FILLER_ASAP7_75t_R FILLER_0_92_26 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_34 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_56 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_78 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_100 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_122 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_144 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_166 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_188 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_210 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_228 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_238 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_283 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_305 ();
 DECAPx2_ASAP7_75t_R FILLER_0_92_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_373 ();
 FILLER_ASAP7_75t_R FILLER_0_92_399 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_407 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_427 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_449 ();
 FILLER_ASAP7_75t_R FILLER_0_92_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_486 ();
 FILLER_ASAP7_75t_R FILLER_0_92_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_532 ();
 DECAPx4_ASAP7_75t_R FILLER_0_92_554 ();
 FILLER_ASAP7_75t_R FILLER_0_92_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_566 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_588 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_610 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_632 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_654 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_676 ();
 DECAPx10_ASAP7_75t_R FILLER_0_92_698 ();
 DECAPx6_ASAP7_75t_R FILLER_0_92_720 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_734 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_92_738 ();
 DECAPx1_ASAP7_75t_R FILLER_0_92_749 ();
 DECAPx4_ASAP7_75t_R FILLER_0_93_2 ();
 FILLER_ASAP7_75t_R FILLER_0_93_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_14 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_30 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_52 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_74 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_96 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_206 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_228 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_250 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_294 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_316 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_352 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_374 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_388 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_402 ();
 DECAPx4_ASAP7_75t_R FILLER_0_93_424 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_438 ();
 FILLER_ASAP7_75t_R FILLER_0_93_448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_471 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_493 ();
 DECAPx6_ASAP7_75t_R FILLER_0_93_518 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_558 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_580 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_602 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_624 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_646 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_668 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_93_712 ();
 DECAPx2_ASAP7_75t_R FILLER_0_93_734 ();
 FILLER_ASAP7_75t_R FILLER_0_93_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_742 ();
 DECAPx1_ASAP7_75t_R FILLER_0_93_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_93_757 ();
 FILLER_ASAP7_75t_R FILLER_0_94_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_4 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_10 ();
 FILLER_ASAP7_75t_R FILLER_0_94_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_18 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_178 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_200 ();
 FILLER_ASAP7_75t_R FILLER_0_94_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_216 ();
 FILLER_ASAP7_75t_R FILLER_0_94_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_245 ();
 DECAPx4_ASAP7_75t_R FILLER_0_94_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_277 ();
 FILLER_ASAP7_75t_R FILLER_0_94_281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_327 ();
 DECAPx4_ASAP7_75t_R FILLER_0_94_331 ();
 DECAPx4_ASAP7_75t_R FILLER_0_94_363 ();
 FILLER_ASAP7_75t_R FILLER_0_94_373 ();
 FILLER_ASAP7_75t_R FILLER_0_94_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_395 ();
 FILLER_ASAP7_75t_R FILLER_0_94_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_426 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_433 ();
 FILLER_ASAP7_75t_R FILLER_0_94_439 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_486 ();
 FILLER_ASAP7_75t_R FILLER_0_94_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_494 ();
 DECAPx2_ASAP7_75t_R FILLER_0_94_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_587 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_609 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_631 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_653 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_675 ();
 DECAPx10_ASAP7_75t_R FILLER_0_94_697 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_723 ();
 DECAPx6_ASAP7_75t_R FILLER_0_94_729 ();
 DECAPx1_ASAP7_75t_R FILLER_0_94_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_94_752 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_7 ();
 DECAPx1_ASAP7_75t_R FILLER_0_95_21 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_35 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_57 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_79 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_101 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_123 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_145 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_167 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_189 ();
 FILLER_ASAP7_75t_R FILLER_0_95_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_197 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_201 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_223 ();
 FILLER_ASAP7_75t_R FILLER_0_95_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_231 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_254 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_276 ();
 DECAPx4_ASAP7_75t_R FILLER_0_95_298 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_314 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_336 ();
 DECAPx4_ASAP7_75t_R FILLER_0_95_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_368 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_396 ();
 FILLER_ASAP7_75t_R FILLER_0_95_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_404 ();
 FILLER_ASAP7_75t_R FILLER_0_95_409 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_421 ();
 DECAPx6_ASAP7_75t_R FILLER_0_95_506 ();
 DECAPx2_ASAP7_75t_R FILLER_0_95_520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_547 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_569 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_591 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_613 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_635 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_657 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_679 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_701 ();
 DECAPx10_ASAP7_75t_R FILLER_0_95_723 ();
 FILLER_ASAP7_75t_R FILLER_0_95_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_95_752 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_2 ();
 FILLER_ASAP7_75t_R FILLER_0_96_8 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_15 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_19 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_30 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_52 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_74 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_96 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_118 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_140 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_162 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_184 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_206 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_228 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_246 ();
 DECAPx4_ASAP7_75t_R FILLER_0_96_250 ();
 FILLER_ASAP7_75t_R FILLER_0_96_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_262 ();
 DECAPx4_ASAP7_75t_R FILLER_0_96_285 ();
 FILLER_ASAP7_75t_R FILLER_0_96_295 ();
 DECAPx4_ASAP7_75t_R FILLER_0_96_300 ();
 FILLER_ASAP7_75t_R FILLER_0_96_332 ();
 FILLER_ASAP7_75t_R FILLER_0_96_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_376 ();
 FILLER_ASAP7_75t_R FILLER_0_96_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_403 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_486 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_508 ();
 FILLER_ASAP7_75t_R FILLER_0_96_514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_537 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_559 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_603 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_647 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_669 ();
 DECAPx10_ASAP7_75t_R FILLER_0_96_691 ();
 DECAPx6_ASAP7_75t_R FILLER_0_96_713 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_727 ();
 DECAPx1_ASAP7_75t_R FILLER_0_96_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_745 ();
 DECAPx2_ASAP7_75t_R FILLER_0_96_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_96_757 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_12 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_49 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_71 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_93 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_115 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_137 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_159 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_181 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_203 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_225 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_247 ();
 DECAPx2_ASAP7_75t_R FILLER_0_97_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_275 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_297 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_319 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_341 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_377 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_400 ();
 FILLER_ASAP7_75t_R FILLER_0_97_410 ();
 DECAPx4_ASAP7_75t_R FILLER_0_97_416 ();
 FILLER_ASAP7_75t_R FILLER_0_97_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_428 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_433 ();
 FILLER_ASAP7_75t_R FILLER_0_97_447 ();
 DECAPx6_ASAP7_75t_R FILLER_0_97_470 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_484 ();
 FILLER_ASAP7_75t_R FILLER_0_97_509 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_97_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_730 ();
 DECAPx1_ASAP7_75t_R FILLER_0_97_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_97_750 ();
 FILLER_ASAP7_75t_R FILLER_0_97_756 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_26 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_48 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_70 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_92 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_114 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_136 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_158 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_180 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_202 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_224 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_246 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_268 ();
 DECAPx4_ASAP7_75t_R FILLER_0_98_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_300 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_332 ();
 DECAPx1_ASAP7_75t_R FILLER_0_98_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_369 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_388 ();
 DECAPx4_ASAP7_75t_R FILLER_0_98_395 ();
 FILLER_ASAP7_75t_R FILLER_0_98_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_461 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_464 ();
 DECAPx2_ASAP7_75t_R FILLER_0_98_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_484 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_550 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_594 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_638 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_98_704 ();
 DECAPx4_ASAP7_75t_R FILLER_0_98_726 ();
 FILLER_ASAP7_75t_R FILLER_0_98_736 ();
 DECAPx6_ASAP7_75t_R FILLER_0_98_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_98_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_2 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_8 ();
 FILLER_ASAP7_75t_R FILLER_0_99_18 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_20 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_27 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_49 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_71 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_93 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_115 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_137 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_159 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_181 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_203 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_225 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_247 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_269 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_291 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_335 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_357 ();
 DECAPx4_ASAP7_75t_R FILLER_0_99_402 ();
 FILLER_ASAP7_75t_R FILLER_0_99_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_471 ();
 DECAPx6_ASAP7_75t_R FILLER_0_99_493 ();
 FILLER_ASAP7_75t_R FILLER_0_99_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_509 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_531 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_553 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_575 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_597 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_641 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_663 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_685 ();
 DECAPx10_ASAP7_75t_R FILLER_0_99_707 ();
 DECAPx2_ASAP7_75t_R FILLER_0_99_749 ();
 FILLER_ASAP7_75t_R FILLER_0_99_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_99_757 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_2 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_16 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_28 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_39 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_61 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_83 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_105 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_127 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_149 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_171 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_193 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_215 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_237 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_259 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_281 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_303 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_325 ();
 DECAPx4_ASAP7_75t_R FILLER_0_100_361 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_406 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_432 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_454 ();
 FILLER_ASAP7_75t_R FILLER_0_100_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_558 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_580 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_602 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_624 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_646 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_668 ();
 DECAPx10_ASAP7_75t_R FILLER_0_100_690 ();
 DECAPx6_ASAP7_75t_R FILLER_0_100_712 ();
 DECAPx2_ASAP7_75t_R FILLER_0_100_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_737 ();
 DECAPx1_ASAP7_75t_R FILLER_0_100_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_100_747 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_244 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_266 ();
 FILLER_ASAP7_75t_R FILLER_0_101_276 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_309 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_352 ();
 FILLER_ASAP7_75t_R FILLER_0_101_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_376 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_399 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_430 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_452 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_474 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_496 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_518 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_540 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_562 ();
 DECAPx2_ASAP7_75t_R FILLER_0_101_584 ();
 FILLER_ASAP7_75t_R FILLER_0_101_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_101_592 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_101_686 ();
 DECAPx6_ASAP7_75t_R FILLER_0_101_708 ();
 FILLER_ASAP7_75t_R FILLER_0_101_722 ();
 DECAPx4_ASAP7_75t_R FILLER_0_101_729 ();
 DECAPx1_ASAP7_75t_R FILLER_0_101_749 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_266 ();
 DECAPx6_ASAP7_75t_R FILLER_0_102_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_308 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_341 ();
 DECAPx4_ASAP7_75t_R FILLER_0_102_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_396 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_400 ();
 DECAPx6_ASAP7_75t_R FILLER_0_102_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_102_436 ();
 DECAPx1_ASAP7_75t_R FILLER_0_102_458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_102_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_102_750 ();
 FILLER_ASAP7_75t_R FILLER_0_102_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_266 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_292 ();
 DECAPx6_ASAP7_75t_R FILLER_0_103_314 ();
 DECAPx2_ASAP7_75t_R FILLER_0_103_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_341 ();
 DECAPx1_ASAP7_75t_R FILLER_0_103_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_367 ();
 DECAPx6_ASAP7_75t_R FILLER_0_103_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_103_426 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_558 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_580 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_602 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_624 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_646 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_668 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_712 ();
 DECAPx10_ASAP7_75t_R FILLER_0_103_734 ();
 FILLER_ASAP7_75t_R FILLER_0_103_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_104_266 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_286 ();
 DECAPx6_ASAP7_75t_R FILLER_0_104_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_322 ();
 DECAPx4_ASAP7_75t_R FILLER_0_104_344 ();
 FILLER_ASAP7_75t_R FILLER_0_104_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_356 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_363 ();
 FILLER_ASAP7_75t_R FILLER_0_104_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_415 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_437 ();
 FILLER_ASAP7_75t_R FILLER_0_104_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_104_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_104_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_104_750 ();
 FILLER_ASAP7_75t_R FILLER_0_104_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_288 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_310 ();
 FILLER_ASAP7_75t_R FILLER_0_105_320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_388 ();
 DECAPx4_ASAP7_75t_R FILLER_0_105_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_105_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_446 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_512 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_534 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_556 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_578 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_600 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_622 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_644 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_666 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_688 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_710 ();
 DECAPx10_ASAP7_75t_R FILLER_0_105_732 ();
 DECAPx1_ASAP7_75t_R FILLER_0_105_754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_266 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_288 ();
 FILLER_ASAP7_75t_R FILLER_0_106_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_296 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_318 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_340 ();
 DECAPx1_ASAP7_75t_R FILLER_0_106_362 ();
 DECAPx4_ASAP7_75t_R FILLER_0_106_397 ();
 FILLER_ASAP7_75t_R FILLER_0_106_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_409 ();
 FILLER_ASAP7_75t_R FILLER_0_106_416 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_427 ();
 DECAPx4_ASAP7_75t_R FILLER_0_106_449 ();
 FILLER_ASAP7_75t_R FILLER_0_106_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_106_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_106_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_106_750 ();
 FILLER_ASAP7_75t_R FILLER_0_106_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_200 ();
 DECAPx4_ASAP7_75t_R FILLER_0_107_222 ();
 FILLER_ASAP7_75t_R FILLER_0_107_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_250 ();
 DECAPx1_ASAP7_75t_R FILLER_0_107_272 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_297 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_341 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_362 ();
 DECAPx4_ASAP7_75t_R FILLER_0_107_384 ();
 FILLER_ASAP7_75t_R FILLER_0_107_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_107_396 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_418 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_440 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_484 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_550 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_594 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_638 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_704 ();
 DECAPx10_ASAP7_75t_R FILLER_0_107_726 ();
 DECAPx4_ASAP7_75t_R FILLER_0_107_748 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_200 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_222 ();
 FILLER_ASAP7_75t_R FILLER_0_108_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_234 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_257 ();
 DECAPx6_ASAP7_75t_R FILLER_0_108_279 ();
 DECAPx1_ASAP7_75t_R FILLER_0_108_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_304 ();
 DECAPx4_ASAP7_75t_R FILLER_0_108_331 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_368 ();
 FILLER_ASAP7_75t_R FILLER_0_108_390 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_426 ();
 FILLER_ASAP7_75t_R FILLER_0_108_432 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_108_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_108_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_108_750 ();
 FILLER_ASAP7_75t_R FILLER_0_108_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_222 ();
 DECAPx6_ASAP7_75t_R FILLER_0_109_244 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_258 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_285 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_311 ();
 DECAPx1_ASAP7_75t_R FILLER_0_109_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_357 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_379 ();
 FILLER_ASAP7_75t_R FILLER_0_109_385 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_399 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_421 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_443 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_465 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_487 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_509 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_531 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_553 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_575 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_597 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_641 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_663 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_685 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_707 ();
 DECAPx10_ASAP7_75t_R FILLER_0_109_729 ();
 DECAPx2_ASAP7_75t_R FILLER_0_109_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_109_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_266 ();
 FILLER_ASAP7_75t_R FILLER_0_110_280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_324 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_352 ();
 DECAPx4_ASAP7_75t_R FILLER_0_110_382 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_414 ();
 FILLER_ASAP7_75t_R FILLER_0_110_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_110_422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_426 ();
 DECAPx6_ASAP7_75t_R FILLER_0_110_448 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_110_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_110_750 ();
 FILLER_ASAP7_75t_R FILLER_0_110_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_111_332 ();
 DECAPx4_ASAP7_75t_R FILLER_0_111_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_383 ();
 DECAPx1_ASAP7_75t_R FILLER_0_111_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_433 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_455 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_477 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_499 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_587 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_609 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_631 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_653 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_675 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_697 ();
 DECAPx10_ASAP7_75t_R FILLER_0_111_719 ();
 DECAPx6_ASAP7_75t_R FILLER_0_111_741 ();
 FILLER_ASAP7_75t_R FILLER_0_111_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_111_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_112_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_112_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_359 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_363 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_385 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_407 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_429 ();
 DECAPx4_ASAP7_75t_R FILLER_0_112_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_112_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_112_750 ();
 FILLER_ASAP7_75t_R FILLER_0_112_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_310 ();
 FILLER_ASAP7_75t_R FILLER_0_113_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_334 ();
 DECAPx6_ASAP7_75t_R FILLER_0_113_341 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_113_367 ();
 DECAPx6_ASAP7_75t_R FILLER_0_113_393 ();
 FILLER_ASAP7_75t_R FILLER_0_113_407 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_430 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_452 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_474 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_496 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_518 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_540 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_562 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_584 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_606 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_672 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_694 ();
 DECAPx10_ASAP7_75t_R FILLER_0_113_716 ();
 DECAPx6_ASAP7_75t_R FILLER_0_113_738 ();
 DECAPx2_ASAP7_75t_R FILLER_0_113_752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_266 ();
 DECAPx1_ASAP7_75t_R FILLER_0_114_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_292 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_342 ();
 FILLER_ASAP7_75t_R FILLER_0_114_348 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_377 ();
 FILLER_ASAP7_75t_R FILLER_0_114_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_385 ();
 FILLER_ASAP7_75t_R FILLER_0_114_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_394 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_401 ();
 FILLER_ASAP7_75t_R FILLER_0_114_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_114_409 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_432 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_454 ();
 FILLER_ASAP7_75t_R FILLER_0_114_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_114_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_114_750 ();
 FILLER_ASAP7_75t_R FILLER_0_114_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_266 ();
 DECAPx6_ASAP7_75t_R FILLER_0_115_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_115_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_308 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_376 ();
 DECAPx1_ASAP7_75t_R FILLER_0_115_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_403 ();
 DECAPx4_ASAP7_75t_R FILLER_0_115_424 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_455 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_477 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_499 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_587 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_609 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_631 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_653 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_675 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_697 ();
 DECAPx10_ASAP7_75t_R FILLER_0_115_719 ();
 DECAPx6_ASAP7_75t_R FILLER_0_115_741 ();
 FILLER_ASAP7_75t_R FILLER_0_115_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_115_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_288 ();
 DECAPx4_ASAP7_75t_R FILLER_0_116_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_326 ();
 FILLER_ASAP7_75t_R FILLER_0_116_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_334 ();
 FILLER_ASAP7_75t_R FILLER_0_116_358 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_116_388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_438 ();
 FILLER_ASAP7_75t_R FILLER_0_116_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_116_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_116_750 ();
 FILLER_ASAP7_75t_R FILLER_0_116_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_266 ();
 DECAPx6_ASAP7_75t_R FILLER_0_117_288 ();
 FILLER_ASAP7_75t_R FILLER_0_117_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_304 ();
 DECAPx6_ASAP7_75t_R FILLER_0_117_347 ();
 FILLER_ASAP7_75t_R FILLER_0_117_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_363 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_385 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_407 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_451 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_473 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_495 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_517 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_539 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_561 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_583 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_605 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_627 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_649 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_671 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_693 ();
 DECAPx10_ASAP7_75t_R FILLER_0_117_715 ();
 DECAPx6_ASAP7_75t_R FILLER_0_117_737 ();
 DECAPx2_ASAP7_75t_R FILLER_0_117_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_117_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_266 ();
 FILLER_ASAP7_75t_R FILLER_0_118_280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_303 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_325 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_347 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_367 ();
 DECAPx4_ASAP7_75t_R FILLER_0_118_390 ();
 FILLER_ASAP7_75t_R FILLER_0_118_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_402 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_118_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_424 ();
 DECAPx6_ASAP7_75t_R FILLER_0_118_446 ();
 FILLER_ASAP7_75t_R FILLER_0_118_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_118_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_118_750 ();
 FILLER_ASAP7_75t_R FILLER_0_118_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_310 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_332 ();
 FILLER_ASAP7_75t_R FILLER_0_119_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_344 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_351 ();
 DECAPx4_ASAP7_75t_R FILLER_0_119_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_374 ();
 FILLER_ASAP7_75t_R FILLER_0_119_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_383 ();
 FILLER_ASAP7_75t_R FILLER_0_119_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_418 ();
 FILLER_ASAP7_75t_R FILLER_0_119_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_449 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_471 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_493 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_515 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_537 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_559 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_603 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_647 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_669 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_691 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_713 ();
 DECAPx10_ASAP7_75t_R FILLER_0_119_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_119_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_120_332 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_120_352 ();
 DECAPx4_ASAP7_75t_R FILLER_0_120_365 ();
 FILLER_ASAP7_75t_R FILLER_0_120_375 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_120_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_120_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_120_750 ();
 FILLER_ASAP7_75t_R FILLER_0_120_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_310 ();
 FILLER_ASAP7_75t_R FILLER_0_121_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_355 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_121_383 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_406 ();
 FILLER_ASAP7_75t_R FILLER_0_121_412 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_435 ();
 FILLER_ASAP7_75t_R FILLER_0_121_441 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_121_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_121_750 ();
 FILLER_ASAP7_75t_R FILLER_0_121_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_316 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_323 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_345 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_122_373 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_380 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_402 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_424 ();
 DECAPx6_ASAP7_75t_R FILLER_0_122_446 ();
 FILLER_ASAP7_75t_R FILLER_0_122_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_122_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_122_750 ();
 FILLER_ASAP7_75t_R FILLER_0_122_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_244 ();
 DECAPx6_ASAP7_75t_R FILLER_0_123_266 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_280 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_307 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_333 ();
 DECAPx2_ASAP7_75t_R FILLER_0_123_378 ();
 FILLER_ASAP7_75t_R FILLER_0_123_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_386 ();
 DECAPx1_ASAP7_75t_R FILLER_0_123_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_123_397 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_419 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_462 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_484 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_550 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_594 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_638 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_704 ();
 DECAPx10_ASAP7_75t_R FILLER_0_123_726 ();
 DECAPx4_ASAP7_75t_R FILLER_0_123_748 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_310 ();
 FILLER_ASAP7_75t_R FILLER_0_124_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_334 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_359 ();
 FILLER_ASAP7_75t_R FILLER_0_124_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_383 ();
 DECAPx6_ASAP7_75t_R FILLER_0_124_387 ();
 DECAPx1_ASAP7_75t_R FILLER_0_124_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_405 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_409 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_431 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_453 ();
 FILLER_ASAP7_75t_R FILLER_0_124_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_124_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_124_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_124_750 ();
 FILLER_ASAP7_75t_R FILLER_0_124_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_332 ();
 FILLER_ASAP7_75t_R FILLER_0_125_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_377 ();
 DECAPx2_ASAP7_75t_R FILLER_0_125_399 ();
 FILLER_ASAP7_75t_R FILLER_0_125_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_407 ();
 DECAPx1_ASAP7_75t_R FILLER_0_125_429 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_439 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_483 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_505 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_527 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_549 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_571 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_593 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_615 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_637 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_659 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_681 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_703 ();
 DECAPx10_ASAP7_75t_R FILLER_0_125_725 ();
 DECAPx4_ASAP7_75t_R FILLER_0_125_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_125_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_420 ();
 DECAPx6_ASAP7_75t_R FILLER_0_126_442 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_456 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_126_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_126_750 ();
 FILLER_ASAP7_75t_R FILLER_0_126_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_354 ();
 FILLER_ASAP7_75t_R FILLER_0_127_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_384 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_406 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_428 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_450 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_472 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_494 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_516 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_560 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_604 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_626 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_648 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_670 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_692 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_714 ();
 DECAPx10_ASAP7_75t_R FILLER_0_127_736 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_354 ();
 DECAPx6_ASAP7_75t_R FILLER_0_128_376 ();
 DECAPx1_ASAP7_75t_R FILLER_0_128_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_394 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_416 ();
 FILLER_ASAP7_75t_R FILLER_0_128_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_128_440 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_128_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_128_750 ();
 FILLER_ASAP7_75t_R FILLER_0_128_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_310 ();
 DECAPx6_ASAP7_75t_R FILLER_0_129_332 ();
 FILLER_ASAP7_75t_R FILLER_0_129_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_348 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_370 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_392 ();
 FILLER_ASAP7_75t_R FILLER_0_129_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_129_400 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_444 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_466 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_488 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_510 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_532 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_554 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_576 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_598 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_620 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_642 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_664 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_686 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_708 ();
 DECAPx10_ASAP7_75t_R FILLER_0_129_730 ();
 DECAPx2_ASAP7_75t_R FILLER_0_129_752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_376 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_130_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_411 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_438 ();
 FILLER_ASAP7_75t_R FILLER_0_130_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_130_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_130_750 ();
 FILLER_ASAP7_75t_R FILLER_0_130_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_131_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_131_750 ();
 FILLER_ASAP7_75t_R FILLER_0_131_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_332 ();
 DECAPx6_ASAP7_75t_R FILLER_0_132_354 ();
 FILLER_ASAP7_75t_R FILLER_0_132_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_132_370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_392 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_414 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_436 ();
 DECAPx1_ASAP7_75t_R FILLER_0_132_458 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_470 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_514 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_536 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_558 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_580 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_602 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_624 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_646 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_668 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_690 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_712 ();
 DECAPx10_ASAP7_75t_R FILLER_0_132_734 ();
 FILLER_ASAP7_75t_R FILLER_0_132_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_420 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_442 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_133_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_133_750 ();
 FILLER_ASAP7_75t_R FILLER_0_133_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_288 ();
 DECAPx4_ASAP7_75t_R FILLER_0_134_310 ();
 FILLER_ASAP7_75t_R FILLER_0_134_320 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_343 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_365 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_387 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_409 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_431 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_453 ();
 FILLER_ASAP7_75t_R FILLER_0_134_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_134_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_134_750 ();
 FILLER_ASAP7_75t_R FILLER_0_134_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_354 ();
 DECAPx4_ASAP7_75t_R FILLER_0_135_376 ();
 FILLER_ASAP7_75t_R FILLER_0_135_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_388 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_410 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_432 ();
 DECAPx6_ASAP7_75t_R FILLER_0_135_454 ();
 FILLER_ASAP7_75t_R FILLER_0_135_468 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_491 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_535 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_579 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_601 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_623 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_645 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_667 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_689 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_711 ();
 DECAPx10_ASAP7_75t_R FILLER_0_135_733 ();
 FILLER_ASAP7_75t_R FILLER_0_135_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_135_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_398 ();
 DECAPx6_ASAP7_75t_R FILLER_0_136_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_434 ();
 DECAPx6_ASAP7_75t_R FILLER_0_136_441 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_136_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_136_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_136_750 ();
 FILLER_ASAP7_75t_R FILLER_0_136_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_354 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_376 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_398 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_420 ();
 DECAPx4_ASAP7_75t_R FILLER_0_137_442 ();
 FILLER_ASAP7_75t_R FILLER_0_137_452 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_476 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_498 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_520 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_542 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_564 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_586 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_608 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_630 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_652 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_674 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_696 ();
 DECAPx10_ASAP7_75t_R FILLER_0_137_718 ();
 DECAPx6_ASAP7_75t_R FILLER_0_137_740 ();
 DECAPx1_ASAP7_75t_R FILLER_0_137_754 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_332 ();
 DECAPx6_ASAP7_75t_R FILLER_0_138_354 ();
 FILLER_ASAP7_75t_R FILLER_0_138_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_370 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_397 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_413 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_435 ();
 DECAPx1_ASAP7_75t_R FILLER_0_138_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_461 ();
 DECAPx6_ASAP7_75t_R FILLER_0_138_464 ();
 FILLER_ASAP7_75t_R FILLER_0_138_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_138_480 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_484 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_506 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_528 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_550 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_572 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_594 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_616 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_638 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_660 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_682 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_704 ();
 DECAPx10_ASAP7_75t_R FILLER_0_138_726 ();
 DECAPx4_ASAP7_75t_R FILLER_0_138_748 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_288 ();
 DECAPx6_ASAP7_75t_R FILLER_0_139_310 ();
 DECAPx1_ASAP7_75t_R FILLER_0_139_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_139_328 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_350 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_372 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_394 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_416 ();
 FILLER_ASAP7_75t_R FILLER_0_139_422 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_452 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_474 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_496 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_518 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_540 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_562 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_584 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_606 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_628 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_650 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_672 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_694 ();
 DECAPx10_ASAP7_75t_R FILLER_0_139_716 ();
 DECAPx6_ASAP7_75t_R FILLER_0_139_738 ();
 DECAPx2_ASAP7_75t_R FILLER_0_139_752 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_310 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_140_338 ();
 DECAPx4_ASAP7_75t_R FILLER_0_140_369 ();
 FILLER_ASAP7_75t_R FILLER_0_140_379 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_408 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_430 ();
 DECAPx4_ASAP7_75t_R FILLER_0_140_452 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_140_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_140_750 ();
 FILLER_ASAP7_75t_R FILLER_0_140_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_288 ();
 FILLER_ASAP7_75t_R FILLER_0_141_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_312 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_141_364 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_386 ();
 FILLER_ASAP7_75t_R FILLER_0_141_392 ();
 DECAPx1_ASAP7_75t_R FILLER_0_141_415 ();
 DECAPx2_ASAP7_75t_R FILLER_0_141_441 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_472 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_494 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_516 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_538 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_560 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_582 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_604 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_626 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_648 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_670 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_692 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_714 ();
 DECAPx10_ASAP7_75t_R FILLER_0_141_736 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_244 ();
 DECAPx4_ASAP7_75t_R FILLER_0_142_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_297 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_319 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_341 ();
 DECAPx4_ASAP7_75t_R FILLER_0_142_363 ();
 DECAPx6_ASAP7_75t_R FILLER_0_142_401 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_415 ();
 DECAPx6_ASAP7_75t_R FILLER_0_142_443 ();
 DECAPx1_ASAP7_75t_R FILLER_0_142_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_142_461 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_486 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_508 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_530 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_552 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_574 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_596 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_618 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_640 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_662 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_684 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_706 ();
 DECAPx10_ASAP7_75t_R FILLER_0_142_728 ();
 DECAPx2_ASAP7_75t_R FILLER_0_142_750 ();
 FILLER_ASAP7_75t_R FILLER_0_142_756 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_310 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_332 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_354 ();
 DECAPx6_ASAP7_75t_R FILLER_0_143_376 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_390 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_401 ();
 FILLER_ASAP7_75t_R FILLER_0_143_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_410 ();
 DECAPx1_ASAP7_75t_R FILLER_0_143_440 ();
 DECAPx2_ASAP7_75t_R FILLER_0_143_466 ();
 FILLER_ASAP7_75t_R FILLER_0_143_472 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_477 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_499 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_587 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_609 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_631 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_653 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_675 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_697 ();
 DECAPx10_ASAP7_75t_R FILLER_0_143_719 ();
 DECAPx6_ASAP7_75t_R FILLER_0_143_741 ();
 FILLER_ASAP7_75t_R FILLER_0_143_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_143_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_310 ();
 FILLER_ASAP7_75t_R FILLER_0_144_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_318 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_382 ();
 DECAPx4_ASAP7_75t_R FILLER_0_144_404 ();
 DECAPx2_ASAP7_75t_R FILLER_0_144_434 ();
 DECAPx6_ASAP7_75t_R FILLER_0_144_443 ();
 DECAPx1_ASAP7_75t_R FILLER_0_144_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_461 ();
 FILLER_ASAP7_75t_R FILLER_0_144_464 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_469 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_491 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_535 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_579 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_601 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_623 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_645 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_667 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_689 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_711 ();
 DECAPx10_ASAP7_75t_R FILLER_0_144_733 ();
 FILLER_ASAP7_75t_R FILLER_0_144_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_288 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_332 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_360 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_367 ();
 DECAPx2_ASAP7_75t_R FILLER_0_145_389 ();
 FILLER_ASAP7_75t_R FILLER_0_145_395 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_418 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_444 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_465 ();
 FILLER_ASAP7_75t_R FILLER_0_145_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_471 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_475 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_497 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_519 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_541 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_563 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_585 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_607 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_629 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_651 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_673 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_695 ();
 DECAPx10_ASAP7_75t_R FILLER_0_145_717 ();
 DECAPx6_ASAP7_75t_R FILLER_0_145_739 ();
 DECAPx1_ASAP7_75t_R FILLER_0_145_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_145_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_244 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_288 ();
 DECAPx2_ASAP7_75t_R FILLER_0_146_310 ();
 FILLER_ASAP7_75t_R FILLER_0_146_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_318 ();
 DECAPx1_ASAP7_75t_R FILLER_0_146_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_328 ();
 FILLER_ASAP7_75t_R FILLER_0_146_339 ();
 DECAPx6_ASAP7_75t_R FILLER_0_146_346 ();
 DECAPx6_ASAP7_75t_R FILLER_0_146_385 ();
 DECAPx4_ASAP7_75t_R FILLER_0_146_420 ();
 FILLER_ASAP7_75t_R FILLER_0_146_430 ();
 DECAPx6_ASAP7_75t_R FILLER_0_146_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_456 ();
 FILLER_ASAP7_75t_R FILLER_0_146_460 ();
 DECAPx4_ASAP7_75t_R FILLER_0_146_464 ();
 FILLER_ASAP7_75t_R FILLER_0_146_474 ();
 DECAPx4_ASAP7_75t_R FILLER_0_146_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_489 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_493 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_515 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_537 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_559 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_581 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_603 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_647 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_669 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_691 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_713 ();
 DECAPx10_ASAP7_75t_R FILLER_0_146_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_146_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_244 ();
 DECAPx4_ASAP7_75t_R FILLER_0_147_266 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_281 ();
 FILLER_ASAP7_75t_R FILLER_0_147_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_305 ();
 FILLER_ASAP7_75t_R FILLER_0_147_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_354 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_370 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_384 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_406 ();
 FILLER_ASAP7_75t_R FILLER_0_147_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_474 ();
 DECAPx2_ASAP7_75t_R FILLER_0_147_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_487 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_491 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_513 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_535 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_557 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_579 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_601 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_623 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_645 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_667 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_689 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_711 ();
 DECAPx10_ASAP7_75t_R FILLER_0_147_733 ();
 FILLER_ASAP7_75t_R FILLER_0_147_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_147_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_222 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_244 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_280 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_315 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_325 ();
 FILLER_ASAP7_75t_R FILLER_0_148_382 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_389 ();
 DECAPx2_ASAP7_75t_R FILLER_0_148_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_433 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_440 ();
 DECAPx4_ASAP7_75t_R FILLER_0_148_447 ();
 DECAPx1_ASAP7_75t_R FILLER_0_148_492 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_499 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_521 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_543 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_565 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_587 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_609 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_631 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_653 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_675 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_697 ();
 DECAPx10_ASAP7_75t_R FILLER_0_148_719 ();
 DECAPx6_ASAP7_75t_R FILLER_0_148_741 ();
 FILLER_ASAP7_75t_R FILLER_0_148_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_148_757 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_222 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_244 ();
 DECAPx2_ASAP7_75t_R FILLER_0_149_258 ();
 FILLER_ASAP7_75t_R FILLER_0_149_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_334 ();
 FILLER_ASAP7_75t_R FILLER_0_149_356 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_409 ();
 DECAPx1_ASAP7_75t_R FILLER_0_149_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_149_419 ();
 FILLER_ASAP7_75t_R FILLER_0_149_490 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_149_722 ();
 DECAPx6_ASAP7_75t_R FILLER_0_149_744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_222 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_258 ();
 FILLER_ASAP7_75t_R FILLER_0_150_285 ();
 FILLER_ASAP7_75t_R FILLER_0_150_292 ();
 FILLER_ASAP7_75t_R FILLER_0_150_362 ();
 FILLER_ASAP7_75t_R FILLER_0_150_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_461 ();
 DECAPx1_ASAP7_75t_R FILLER_0_150_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_473 ();
 FILLER_ASAP7_75t_R FILLER_0_150_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_150_491 ();
 FILLER_ASAP7_75t_R FILLER_0_150_497 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_502 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_524 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_546 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_568 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_590 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_612 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_634 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_656 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_678 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_700 ();
 DECAPx10_ASAP7_75t_R FILLER_0_150_722 ();
 DECAPx6_ASAP7_75t_R FILLER_0_150_744 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_222 ();
 DECAPx4_ASAP7_75t_R FILLER_0_151_244 ();
 FILLER_ASAP7_75t_R FILLER_0_151_254 ();
 FILLER_ASAP7_75t_R FILLER_0_151_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_314 ();
 FILLER_ASAP7_75t_R FILLER_0_151_460 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_509 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_531 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_553 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_575 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_597 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_619 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_641 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_663 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_685 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_707 ();
 DECAPx10_ASAP7_75t_R FILLER_0_151_729 ();
 DECAPx2_ASAP7_75t_R FILLER_0_151_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_151_757 ();
endmodule
