../../nangate45/lef/fakeram45_256x95.lef