module MuxTest_width_1_inputs_1_outputs_4_pipeline_0( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [2:0] io_operation_0, // @[:@6.4]
  input  [2:0] io_operation_1, // @[:@6.4]
  input  [2:0] io_operation_2, // @[:@6.4]
  input  [2:0] io_operation_3, // @[:@6.4]
  input        io_inputs_0, // @[:@6.4]
  output       io_outputs_0, // @[:@6.4]
  output       io_outputs_1, // @[:@6.4]
  output       io_outputs_2, // @[:@6.4]
  output       io_outputs_3 // @[:@6.4]
);
  wire [1:0] _T_244; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 32:53:@8.4]
  wire  _T_245; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 32:53:@9.4]
  wire [1:0] _T_247; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 33:58:@10.4]
  wire  _T_249; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 34:56:@11.4]
  wire  _T_250; // @[Mux.scala 46:19:@12.4]
  wire  _T_251; // @[Mux.scala 46:16:@13.4]
  wire  _T_252; // @[Mux.scala 46:19:@14.4]
  wire [1:0] _T_253; // @[Mux.scala 46:16:@15.4]
  wire  _T_254; // @[Mux.scala 46:19:@16.4]
  wire [1:0] _T_255; // @[Mux.scala 46:16:@17.4]
  wire  _T_256; // @[Mux.scala 46:19:@18.4]
  wire [1:0] _T_257; // @[Mux.scala 46:16:@19.4]
  wire  _T_267; // @[Mux.scala 46:19:@24.4]
  wire  _T_268; // @[Mux.scala 46:16:@25.4]
  wire  _T_269; // @[Mux.scala 46:19:@26.4]
  wire [1:0] _T_270; // @[Mux.scala 46:16:@27.4]
  wire  _T_271; // @[Mux.scala 46:19:@28.4]
  wire [1:0] _T_272; // @[Mux.scala 46:16:@29.4]
  wire  _T_273; // @[Mux.scala 46:19:@30.4]
  wire [1:0] _T_274; // @[Mux.scala 46:16:@31.4]
  wire  _T_284; // @[Mux.scala 46:19:@36.4]
  wire  _T_285; // @[Mux.scala 46:16:@37.4]
  wire  _T_286; // @[Mux.scala 46:19:@38.4]
  wire [1:0] _T_287; // @[Mux.scala 46:16:@39.4]
  wire  _T_288; // @[Mux.scala 46:19:@40.4]
  wire [1:0] _T_289; // @[Mux.scala 46:16:@41.4]
  wire  _T_290; // @[Mux.scala 46:19:@42.4]
  wire [1:0] _T_291; // @[Mux.scala 46:16:@43.4]
  wire  _T_301; // @[Mux.scala 46:19:@48.4]
  wire  _T_302; // @[Mux.scala 46:16:@49.4]
  wire  _T_303; // @[Mux.scala 46:19:@50.4]
  wire [1:0] _T_304; // @[Mux.scala 46:16:@51.4]
  wire  _T_305; // @[Mux.scala 46:19:@52.4]
  wire [1:0] _T_306; // @[Mux.scala 46:16:@53.4]
  wire  _T_307; // @[Mux.scala 46:19:@54.4]
  wire [1:0] _T_308; // @[Mux.scala 46:16:@55.4]
  assign _T_244 = io_inputs_0 + io_inputs_0; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 32:53:@8.4]
  assign _T_245 = io_inputs_0 + io_inputs_0; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 32:53:@9.4]
  assign _T_247 = io_inputs_0 * io_inputs_0; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 33:58:@10.4]
  assign _T_249 = io_inputs_0 / io_inputs_0; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 34:56:@11.4]
  assign _T_250 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_251 = _T_250 ? _T_249 : 1'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_252 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_253 = _T_252 ? _T_247 : {{1'd0}, _T_251}; // @[Mux.scala 46:16:@15.4]
  assign _T_254 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_255 = _T_254 ? {{1'd0}, _T_245} : _T_253; // @[Mux.scala 46:16:@17.4]
  assign _T_256 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _T_257 = _T_256 ? {{1'd0}, io_inputs_0} : _T_255; // @[Mux.scala 46:16:@19.4]
  assign _T_267 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_268 = _T_267 ? _T_249 : 1'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_269 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_270 = _T_269 ? _T_247 : {{1'd0}, _T_268}; // @[Mux.scala 46:16:@27.4]
  assign _T_271 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_272 = _T_271 ? {{1'd0}, _T_245} : _T_270; // @[Mux.scala 46:16:@29.4]
  assign _T_273 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _T_274 = _T_273 ? {{1'd0}, io_inputs_0} : _T_272; // @[Mux.scala 46:16:@31.4]
  assign _T_284 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_285 = _T_284 ? _T_249 : 1'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_286 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_287 = _T_286 ? _T_247 : {{1'd0}, _T_285}; // @[Mux.scala 46:16:@39.4]
  assign _T_288 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_289 = _T_288 ? {{1'd0}, _T_245} : _T_287; // @[Mux.scala 46:16:@41.4]
  assign _T_290 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _T_291 = _T_290 ? {{1'd0}, io_inputs_0} : _T_289; // @[Mux.scala 46:16:@43.4]
  assign _T_301 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_302 = _T_301 ? _T_249 : 1'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_303 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_304 = _T_303 ? _T_247 : {{1'd0}, _T_302}; // @[Mux.scala 46:16:@51.4]
  assign _T_305 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_306 = _T_305 ? {{1'd0}, _T_245} : _T_304; // @[Mux.scala 46:16:@53.4]
  assign _T_307 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _T_308 = _T_307 ? {{1'd0}, io_inputs_0} : _T_306; // @[Mux.scala 46:16:@55.4]
  assign io_outputs_0 = _T_257[0]; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 23:14:@56.4]
  assign io_outputs_1 = _T_274[0]; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 23:14:@57.4]
  assign io_outputs_2 = _T_291[0]; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 23:14:@58.4]
  assign io_outputs_3 = _T_308[0]; // @[MuxTest_width_1_inputs_1_outputs_4_pipeline_0s.scala 23:14:@59.4]
endmodule
