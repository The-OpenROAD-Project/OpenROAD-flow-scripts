../../../../platforms/asap7/lef/fakeram7_64x21.lef