module MuxTest_width_64_inputs_1_outputs_8_pipeline_0( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [2:0]  io_operation_0, // @[:@6.4]
  input  [2:0]  io_operation_1, // @[:@6.4]
  input  [2:0]  io_operation_2, // @[:@6.4]
  input  [2:0]  io_operation_3, // @[:@6.4]
  input  [2:0]  io_operation_4, // @[:@6.4]
  input  [2:0]  io_operation_5, // @[:@6.4]
  input  [2:0]  io_operation_6, // @[:@6.4]
  input  [2:0]  io_operation_7, // @[:@6.4]
  input  [63:0] io_inputs_0, // @[:@6.4]
  output [63:0] io_outputs_0, // @[:@6.4]
  output [63:0] io_outputs_1, // @[:@6.4]
  output [63:0] io_outputs_2, // @[:@6.4]
  output [63:0] io_outputs_3, // @[:@6.4]
  output [63:0] io_outputs_4, // @[:@6.4]
  output [63:0] io_outputs_5, // @[:@6.4]
  output [63:0] io_outputs_6, // @[:@6.4]
  output [63:0] io_outputs_7 // @[:@6.4]
);
  wire [64:0] _T_404; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 32:53:@8.4]
  wire [63:0] _T_405; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 32:53:@9.4]
  wire [127:0] _T_407; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 33:58:@10.4]
  wire [63:0] _T_409; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 34:56:@11.4]
  wire  _T_410; // @[Mux.scala 46:19:@12.4]
  wire [63:0] _T_411; // @[Mux.scala 46:16:@13.4]
  wire  _T_412; // @[Mux.scala 46:19:@14.4]
  wire [127:0] _T_413; // @[Mux.scala 46:16:@15.4]
  wire  _T_414; // @[Mux.scala 46:19:@16.4]
  wire [127:0] _T_415; // @[Mux.scala 46:16:@17.4]
  wire  _T_416; // @[Mux.scala 46:19:@18.4]
  wire [127:0] _T_417; // @[Mux.scala 46:16:@19.4]
  wire  _T_427; // @[Mux.scala 46:19:@24.4]
  wire [63:0] _T_428; // @[Mux.scala 46:16:@25.4]
  wire  _T_429; // @[Mux.scala 46:19:@26.4]
  wire [127:0] _T_430; // @[Mux.scala 46:16:@27.4]
  wire  _T_431; // @[Mux.scala 46:19:@28.4]
  wire [127:0] _T_432; // @[Mux.scala 46:16:@29.4]
  wire  _T_433; // @[Mux.scala 46:19:@30.4]
  wire [127:0] _T_434; // @[Mux.scala 46:16:@31.4]
  wire  _T_444; // @[Mux.scala 46:19:@36.4]
  wire [63:0] _T_445; // @[Mux.scala 46:16:@37.4]
  wire  _T_446; // @[Mux.scala 46:19:@38.4]
  wire [127:0] _T_447; // @[Mux.scala 46:16:@39.4]
  wire  _T_448; // @[Mux.scala 46:19:@40.4]
  wire [127:0] _T_449; // @[Mux.scala 46:16:@41.4]
  wire  _T_450; // @[Mux.scala 46:19:@42.4]
  wire [127:0] _T_451; // @[Mux.scala 46:16:@43.4]
  wire  _T_461; // @[Mux.scala 46:19:@48.4]
  wire [63:0] _T_462; // @[Mux.scala 46:16:@49.4]
  wire  _T_463; // @[Mux.scala 46:19:@50.4]
  wire [127:0] _T_464; // @[Mux.scala 46:16:@51.4]
  wire  _T_465; // @[Mux.scala 46:19:@52.4]
  wire [127:0] _T_466; // @[Mux.scala 46:16:@53.4]
  wire  _T_467; // @[Mux.scala 46:19:@54.4]
  wire [127:0] _T_468; // @[Mux.scala 46:16:@55.4]
  wire  _T_478; // @[Mux.scala 46:19:@60.4]
  wire [63:0] _T_479; // @[Mux.scala 46:16:@61.4]
  wire  _T_480; // @[Mux.scala 46:19:@62.4]
  wire [127:0] _T_481; // @[Mux.scala 46:16:@63.4]
  wire  _T_482; // @[Mux.scala 46:19:@64.4]
  wire [127:0] _T_483; // @[Mux.scala 46:16:@65.4]
  wire  _T_484; // @[Mux.scala 46:19:@66.4]
  wire [127:0] _T_485; // @[Mux.scala 46:16:@67.4]
  wire  _T_495; // @[Mux.scala 46:19:@72.4]
  wire [63:0] _T_496; // @[Mux.scala 46:16:@73.4]
  wire  _T_497; // @[Mux.scala 46:19:@74.4]
  wire [127:0] _T_498; // @[Mux.scala 46:16:@75.4]
  wire  _T_499; // @[Mux.scala 46:19:@76.4]
  wire [127:0] _T_500; // @[Mux.scala 46:16:@77.4]
  wire  _T_501; // @[Mux.scala 46:19:@78.4]
  wire [127:0] _T_502; // @[Mux.scala 46:16:@79.4]
  wire  _T_512; // @[Mux.scala 46:19:@84.4]
  wire [63:0] _T_513; // @[Mux.scala 46:16:@85.4]
  wire  _T_514; // @[Mux.scala 46:19:@86.4]
  wire [127:0] _T_515; // @[Mux.scala 46:16:@87.4]
  wire  _T_516; // @[Mux.scala 46:19:@88.4]
  wire [127:0] _T_517; // @[Mux.scala 46:16:@89.4]
  wire  _T_518; // @[Mux.scala 46:19:@90.4]
  wire [127:0] _T_519; // @[Mux.scala 46:16:@91.4]
  wire  _T_529; // @[Mux.scala 46:19:@96.4]
  wire [63:0] _T_530; // @[Mux.scala 46:16:@97.4]
  wire  _T_531; // @[Mux.scala 46:19:@98.4]
  wire [127:0] _T_532; // @[Mux.scala 46:16:@99.4]
  wire  _T_533; // @[Mux.scala 46:19:@100.4]
  wire [127:0] _T_534; // @[Mux.scala 46:16:@101.4]
  wire  _T_535; // @[Mux.scala 46:19:@102.4]
  wire [127:0] _T_536; // @[Mux.scala 46:16:@103.4]
  assign _T_404 = io_inputs_0 + io_inputs_0; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 32:53:@8.4]
  assign _T_405 = io_inputs_0 + io_inputs_0; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 32:53:@9.4]
  assign _T_407 = io_inputs_0 * io_inputs_0; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 33:58:@10.4]
  assign _T_409 = io_inputs_0 / io_inputs_0; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 34:56:@11.4]
  assign _T_410 = 3'h3 == io_operation_0; // @[Mux.scala 46:19:@12.4]
  assign _T_411 = _T_410 ? _T_409 : 64'h0; // @[Mux.scala 46:16:@13.4]
  assign _T_412 = 3'h2 == io_operation_0; // @[Mux.scala 46:19:@14.4]
  assign _T_413 = _T_412 ? _T_407 : {{64'd0}, _T_411}; // @[Mux.scala 46:16:@15.4]
  assign _T_414 = 3'h1 == io_operation_0; // @[Mux.scala 46:19:@16.4]
  assign _T_415 = _T_414 ? {{64'd0}, _T_405} : _T_413; // @[Mux.scala 46:16:@17.4]
  assign _T_416 = 3'h0 == io_operation_0; // @[Mux.scala 46:19:@18.4]
  assign _T_417 = _T_416 ? {{64'd0}, io_inputs_0} : _T_415; // @[Mux.scala 46:16:@19.4]
  assign _T_427 = 3'h3 == io_operation_1; // @[Mux.scala 46:19:@24.4]
  assign _T_428 = _T_427 ? _T_409 : 64'h0; // @[Mux.scala 46:16:@25.4]
  assign _T_429 = 3'h2 == io_operation_1; // @[Mux.scala 46:19:@26.4]
  assign _T_430 = _T_429 ? _T_407 : {{64'd0}, _T_428}; // @[Mux.scala 46:16:@27.4]
  assign _T_431 = 3'h1 == io_operation_1; // @[Mux.scala 46:19:@28.4]
  assign _T_432 = _T_431 ? {{64'd0}, _T_405} : _T_430; // @[Mux.scala 46:16:@29.4]
  assign _T_433 = 3'h0 == io_operation_1; // @[Mux.scala 46:19:@30.4]
  assign _T_434 = _T_433 ? {{64'd0}, io_inputs_0} : _T_432; // @[Mux.scala 46:16:@31.4]
  assign _T_444 = 3'h3 == io_operation_2; // @[Mux.scala 46:19:@36.4]
  assign _T_445 = _T_444 ? _T_409 : 64'h0; // @[Mux.scala 46:16:@37.4]
  assign _T_446 = 3'h2 == io_operation_2; // @[Mux.scala 46:19:@38.4]
  assign _T_447 = _T_446 ? _T_407 : {{64'd0}, _T_445}; // @[Mux.scala 46:16:@39.4]
  assign _T_448 = 3'h1 == io_operation_2; // @[Mux.scala 46:19:@40.4]
  assign _T_449 = _T_448 ? {{64'd0}, _T_405} : _T_447; // @[Mux.scala 46:16:@41.4]
  assign _T_450 = 3'h0 == io_operation_2; // @[Mux.scala 46:19:@42.4]
  assign _T_451 = _T_450 ? {{64'd0}, io_inputs_0} : _T_449; // @[Mux.scala 46:16:@43.4]
  assign _T_461 = 3'h3 == io_operation_3; // @[Mux.scala 46:19:@48.4]
  assign _T_462 = _T_461 ? _T_409 : 64'h0; // @[Mux.scala 46:16:@49.4]
  assign _T_463 = 3'h2 == io_operation_3; // @[Mux.scala 46:19:@50.4]
  assign _T_464 = _T_463 ? _T_407 : {{64'd0}, _T_462}; // @[Mux.scala 46:16:@51.4]
  assign _T_465 = 3'h1 == io_operation_3; // @[Mux.scala 46:19:@52.4]
  assign _T_466 = _T_465 ? {{64'd0}, _T_405} : _T_464; // @[Mux.scala 46:16:@53.4]
  assign _T_467 = 3'h0 == io_operation_3; // @[Mux.scala 46:19:@54.4]
  assign _T_468 = _T_467 ? {{64'd0}, io_inputs_0} : _T_466; // @[Mux.scala 46:16:@55.4]
  assign _T_478 = 3'h3 == io_operation_4; // @[Mux.scala 46:19:@60.4]
  assign _T_479 = _T_478 ? _T_409 : 64'h0; // @[Mux.scala 46:16:@61.4]
  assign _T_480 = 3'h2 == io_operation_4; // @[Mux.scala 46:19:@62.4]
  assign _T_481 = _T_480 ? _T_407 : {{64'd0}, _T_479}; // @[Mux.scala 46:16:@63.4]
  assign _T_482 = 3'h1 == io_operation_4; // @[Mux.scala 46:19:@64.4]
  assign _T_483 = _T_482 ? {{64'd0}, _T_405} : _T_481; // @[Mux.scala 46:16:@65.4]
  assign _T_484 = 3'h0 == io_operation_4; // @[Mux.scala 46:19:@66.4]
  assign _T_485 = _T_484 ? {{64'd0}, io_inputs_0} : _T_483; // @[Mux.scala 46:16:@67.4]
  assign _T_495 = 3'h3 == io_operation_5; // @[Mux.scala 46:19:@72.4]
  assign _T_496 = _T_495 ? _T_409 : 64'h0; // @[Mux.scala 46:16:@73.4]
  assign _T_497 = 3'h2 == io_operation_5; // @[Mux.scala 46:19:@74.4]
  assign _T_498 = _T_497 ? _T_407 : {{64'd0}, _T_496}; // @[Mux.scala 46:16:@75.4]
  assign _T_499 = 3'h1 == io_operation_5; // @[Mux.scala 46:19:@76.4]
  assign _T_500 = _T_499 ? {{64'd0}, _T_405} : _T_498; // @[Mux.scala 46:16:@77.4]
  assign _T_501 = 3'h0 == io_operation_5; // @[Mux.scala 46:19:@78.4]
  assign _T_502 = _T_501 ? {{64'd0}, io_inputs_0} : _T_500; // @[Mux.scala 46:16:@79.4]
  assign _T_512 = 3'h3 == io_operation_6; // @[Mux.scala 46:19:@84.4]
  assign _T_513 = _T_512 ? _T_409 : 64'h0; // @[Mux.scala 46:16:@85.4]
  assign _T_514 = 3'h2 == io_operation_6; // @[Mux.scala 46:19:@86.4]
  assign _T_515 = _T_514 ? _T_407 : {{64'd0}, _T_513}; // @[Mux.scala 46:16:@87.4]
  assign _T_516 = 3'h1 == io_operation_6; // @[Mux.scala 46:19:@88.4]
  assign _T_517 = _T_516 ? {{64'd0}, _T_405} : _T_515; // @[Mux.scala 46:16:@89.4]
  assign _T_518 = 3'h0 == io_operation_6; // @[Mux.scala 46:19:@90.4]
  assign _T_519 = _T_518 ? {{64'd0}, io_inputs_0} : _T_517; // @[Mux.scala 46:16:@91.4]
  assign _T_529 = 3'h3 == io_operation_7; // @[Mux.scala 46:19:@96.4]
  assign _T_530 = _T_529 ? _T_409 : 64'h0; // @[Mux.scala 46:16:@97.4]
  assign _T_531 = 3'h2 == io_operation_7; // @[Mux.scala 46:19:@98.4]
  assign _T_532 = _T_531 ? _T_407 : {{64'd0}, _T_530}; // @[Mux.scala 46:16:@99.4]
  assign _T_533 = 3'h1 == io_operation_7; // @[Mux.scala 46:19:@100.4]
  assign _T_534 = _T_533 ? {{64'd0}, _T_405} : _T_532; // @[Mux.scala 46:16:@101.4]
  assign _T_535 = 3'h0 == io_operation_7; // @[Mux.scala 46:19:@102.4]
  assign _T_536 = _T_535 ? {{64'd0}, io_inputs_0} : _T_534; // @[Mux.scala 46:16:@103.4]
  assign io_outputs_0 = _T_417[63:0]; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 23:14:@104.4]
  assign io_outputs_1 = _T_434[63:0]; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 23:14:@105.4]
  assign io_outputs_2 = _T_451[63:0]; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 23:14:@106.4]
  assign io_outputs_3 = _T_468[63:0]; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 23:14:@107.4]
  assign io_outputs_4 = _T_485[63:0]; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 23:14:@108.4]
  assign io_outputs_5 = _T_502[63:0]; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 23:14:@109.4]
  assign io_outputs_6 = _T_519[63:0]; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 23:14:@110.4]
  assign io_outputs_7 = _T_536[63:0]; // @[MuxTest_width_64_inputs_1_outputs_8_pipeline_0s.scala 23:14:@111.4]
endmodule
