VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram_32x46
  FOREIGN fakeram_32x46 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 6.080 BY 8.400 ;
  CLASS BLOCK ;
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.048 0.024 0.072 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.096 0.024 0.120 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.144 0.024 0.168 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.192 0.024 0.216 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.240 0.024 0.264 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.288 0.024 0.312 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.336 0.024 0.360 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.384 0.024 0.408 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.432 0.024 0.456 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.480 0.024 0.504 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.528 0.024 0.552 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.576 0.024 0.600 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.624 0.024 0.648 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.672 0.024 0.696 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.720 0.024 0.744 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.768 0.024 0.792 ;
    END
  END rd_out[15]
  PIN rd_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.816 0.024 0.840 ;
    END
  END rd_out[16]
  PIN rd_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.864 0.024 0.888 ;
    END
  END rd_out[17]
  PIN rd_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.912 0.024 0.936 ;
    END
  END rd_out[18]
  PIN rd_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 0.960 0.024 0.984 ;
    END
  END rd_out[19]
  PIN rd_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.008 0.024 1.032 ;
    END
  END rd_out[20]
  PIN rd_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.056 0.024 1.080 ;
    END
  END rd_out[21]
  PIN rd_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.104 0.024 1.128 ;
    END
  END rd_out[22]
  PIN rd_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.152 0.024 1.176 ;
    END
  END rd_out[23]
  PIN rd_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.200 0.024 1.224 ;
    END
  END rd_out[24]
  PIN rd_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.248 0.024 1.272 ;
    END
  END rd_out[25]
  PIN rd_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.296 0.024 1.320 ;
    END
  END rd_out[26]
  PIN rd_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.344 0.024 1.368 ;
    END
  END rd_out[27]
  PIN rd_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.392 0.024 1.416 ;
    END
  END rd_out[28]
  PIN rd_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.440 0.024 1.464 ;
    END
  END rd_out[29]
  PIN rd_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.488 0.024 1.512 ;
    END
  END rd_out[30]
  PIN rd_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.536 0.024 1.560 ;
    END
  END rd_out[31]
  PIN rd_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.584 0.024 1.608 ;
    END
  END rd_out[32]
  PIN rd_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.632 0.024 1.656 ;
    END
  END rd_out[33]
  PIN rd_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.680 0.024 1.704 ;
    END
  END rd_out[34]
  PIN rd_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.728 0.024 1.752 ;
    END
  END rd_out[35]
  PIN rd_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.776 0.024 1.800 ;
    END
  END rd_out[36]
  PIN rd_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.824 0.024 1.848 ;
    END
  END rd_out[37]
  PIN rd_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.872 0.024 1.896 ;
    END
  END rd_out[38]
  PIN rd_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.920 0.024 1.944 ;
    END
  END rd_out[39]
  PIN rd_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 1.968 0.024 1.992 ;
    END
  END rd_out[40]
  PIN rd_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.016 0.024 2.040 ;
    END
  END rd_out[41]
  PIN rd_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.064 0.024 2.088 ;
    END
  END rd_out[42]
  PIN rd_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.112 0.024 2.136 ;
    END
  END rd_out[43]
  PIN rd_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.160 0.024 2.184 ;
    END
  END rd_out[44]
  PIN rd_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 2.208 0.024 2.232 ;
    END
  END rd_out[45]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.072 0.024 3.096 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.120 0.024 3.144 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.168 0.024 3.192 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.216 0.024 3.240 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.264 0.024 3.288 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.312 0.024 3.336 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.360 0.024 3.384 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.408 0.024 3.432 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.456 0.024 3.480 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.504 0.024 3.528 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.552 0.024 3.576 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.600 0.024 3.624 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.648 0.024 3.672 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.696 0.024 3.720 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.744 0.024 3.768 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.792 0.024 3.816 ;
    END
  END wd_in[15]
  PIN wd_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.840 0.024 3.864 ;
    END
  END wd_in[16]
  PIN wd_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.888 0.024 3.912 ;
    END
  END wd_in[17]
  PIN wd_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.936 0.024 3.960 ;
    END
  END wd_in[18]
  PIN wd_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 3.984 0.024 4.008 ;
    END
  END wd_in[19]
  PIN wd_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.032 0.024 4.056 ;
    END
  END wd_in[20]
  PIN wd_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.080 0.024 4.104 ;
    END
  END wd_in[21]
  PIN wd_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.128 0.024 4.152 ;
    END
  END wd_in[22]
  PIN wd_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.176 0.024 4.200 ;
    END
  END wd_in[23]
  PIN wd_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.224 0.024 4.248 ;
    END
  END wd_in[24]
  PIN wd_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.272 0.024 4.296 ;
    END
  END wd_in[25]
  PIN wd_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.320 0.024 4.344 ;
    END
  END wd_in[26]
  PIN wd_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.368 0.024 4.392 ;
    END
  END wd_in[27]
  PIN wd_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.416 0.024 4.440 ;
    END
  END wd_in[28]
  PIN wd_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.464 0.024 4.488 ;
    END
  END wd_in[29]
  PIN wd_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.512 0.024 4.536 ;
    END
  END wd_in[30]
  PIN wd_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.560 0.024 4.584 ;
    END
  END wd_in[31]
  PIN wd_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.608 0.024 4.632 ;
    END
  END wd_in[32]
  PIN wd_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.656 0.024 4.680 ;
    END
  END wd_in[33]
  PIN wd_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.704 0.024 4.728 ;
    END
  END wd_in[34]
  PIN wd_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.752 0.024 4.776 ;
    END
  END wd_in[35]
  PIN wd_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.800 0.024 4.824 ;
    END
  END wd_in[36]
  PIN wd_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.848 0.024 4.872 ;
    END
  END wd_in[37]
  PIN wd_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.896 0.024 4.920 ;
    END
  END wd_in[38]
  PIN wd_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.944 0.024 4.968 ;
    END
  END wd_in[39]
  PIN wd_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 4.992 0.024 5.016 ;
    END
  END wd_in[40]
  PIN wd_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.040 0.024 5.064 ;
    END
  END wd_in[41]
  PIN wd_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.088 0.024 5.112 ;
    END
  END wd_in[42]
  PIN wd_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.136 0.024 5.160 ;
    END
  END wd_in[43]
  PIN wd_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.184 0.024 5.208 ;
    END
  END wd_in[44]
  PIN wd_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 5.232 0.024 5.256 ;
    END
  END wd_in[45]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.096 0.024 6.120 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.144 0.024 6.168 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.192 0.024 6.216 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.240 0.024 6.264 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 6.288 0.024 6.312 ;
    END
  END addr_in[4]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.152 0.024 7.176 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.200 0.024 7.224 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M4 ;
      RECT 0.000 7.248 0.024 7.272 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.000 6.032 0.096 ;
      RECT 0.048 0.768 6.032 0.864 ;
      RECT 0.048 1.536 6.032 1.632 ;
      RECT 0.048 2.304 6.032 2.400 ;
      RECT 0.048 3.072 6.032 3.168 ;
      RECT 0.048 3.840 6.032 3.936 ;
      RECT 0.048 4.608 6.032 4.704 ;
      RECT 0.048 5.376 6.032 5.472 ;
      RECT 0.048 6.144 6.032 6.240 ;
      RECT 0.048 6.912 6.032 7.008 ;
      RECT 0.048 7.680 6.032 7.776 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
      RECT 0.048 0.384 6.032 0.480 ;
      RECT 0.048 1.152 6.032 1.248 ;
      RECT 0.048 1.920 6.032 2.016 ;
      RECT 0.048 2.688 6.032 2.784 ;
      RECT 0.048 3.456 6.032 3.552 ;
      RECT 0.048 4.224 6.032 4.320 ;
      RECT 0.048 4.992 6.032 5.088 ;
      RECT 0.048 5.760 6.032 5.856 ;
      RECT 0.048 6.528 6.032 6.624 ;
      RECT 0.048 7.296 6.032 7.392 ;
      RECT 0.048 8.064 6.032 8.160 ;
    END
  END VDD
  OBS
    LAYER M1 ;
    RECT 0 0 6.080 8.400 ;
    LAYER M2 ;
    RECT 0 0 6.080 8.400 ;
    LAYER M3 ;
    RECT 0 0 6.080 8.400 ;
    LAYER M4 ;
    RECT 0.024 0 0.048 8.400 ;
    RECT 6.032 0 6.080 8.400 ;
    RECT 0.048 0.000 6.032 0.000 ;
    RECT 0.048 0.096 6.032 0.384 ;
    RECT 0.048 0.480 6.032 0.768 ;
    RECT 0.048 0.864 6.032 1.152 ;
    RECT 0.048 1.248 6.032 1.536 ;
    RECT 0.048 1.632 6.032 1.920 ;
    RECT 0.048 2.016 6.032 2.304 ;
    RECT 0.048 2.400 6.032 2.688 ;
    RECT 0.048 2.784 6.032 3.072 ;
    RECT 0.048 3.168 6.032 3.456 ;
    RECT 0.048 3.552 6.032 3.840 ;
    RECT 0.048 3.936 6.032 4.224 ;
    RECT 0.048 4.320 6.032 4.608 ;
    RECT 0.048 4.704 6.032 4.992 ;
    RECT 0.048 5.088 6.032 5.376 ;
    RECT 0.048 5.472 6.032 5.760 ;
    RECT 0.048 5.856 6.032 6.144 ;
    RECT 0.048 6.240 6.032 6.528 ;
    RECT 0.048 6.624 6.032 6.912 ;
    RECT 0.048 7.008 6.032 7.296 ;
    RECT 0.048 7.392 6.032 7.680 ;
    RECT 0.048 7.776 6.032 8.064 ;
    RECT 0.048 8.160 6.032 8.400 ;
    RECT 0 0.000 0.024 0.048 ;
    RECT 0 0.072 0.024 0.096 ;
    RECT 0 0.120 0.024 0.144 ;
    RECT 0 0.168 0.024 0.192 ;
    RECT 0 0.216 0.024 0.240 ;
    RECT 0 0.264 0.024 0.288 ;
    RECT 0 0.312 0.024 0.336 ;
    RECT 0 0.360 0.024 0.384 ;
    RECT 0 0.408 0.024 0.432 ;
    RECT 0 0.456 0.024 0.480 ;
    RECT 0 0.504 0.024 0.528 ;
    RECT 0 0.552 0.024 0.576 ;
    RECT 0 0.600 0.024 0.624 ;
    RECT 0 0.648 0.024 0.672 ;
    RECT 0 0.696 0.024 0.720 ;
    RECT 0 0.744 0.024 0.768 ;
    RECT 0 0.792 0.024 0.816 ;
    RECT 0 0.840 0.024 0.864 ;
    RECT 0 0.888 0.024 0.912 ;
    RECT 0 0.936 0.024 0.960 ;
    RECT 0 0.984 0.024 1.008 ;
    RECT 0 1.032 0.024 1.056 ;
    RECT 0 1.080 0.024 1.104 ;
    RECT 0 1.128 0.024 1.152 ;
    RECT 0 1.176 0.024 1.200 ;
    RECT 0 1.224 0.024 1.248 ;
    RECT 0 1.272 0.024 1.296 ;
    RECT 0 1.320 0.024 1.344 ;
    RECT 0 1.368 0.024 1.392 ;
    RECT 0 1.416 0.024 1.440 ;
    RECT 0 1.464 0.024 1.488 ;
    RECT 0 1.512 0.024 1.536 ;
    RECT 0 1.560 0.024 1.584 ;
    RECT 0 1.608 0.024 1.632 ;
    RECT 0 1.656 0.024 1.680 ;
    RECT 0 1.704 0.024 1.728 ;
    RECT 0 1.752 0.024 1.776 ;
    RECT 0 1.800 0.024 1.824 ;
    RECT 0 1.848 0.024 1.872 ;
    RECT 0 1.896 0.024 1.920 ;
    RECT 0 1.944 0.024 1.968 ;
    RECT 0 1.992 0.024 2.016 ;
    RECT 0 2.040 0.024 2.064 ;
    RECT 0 2.088 0.024 2.112 ;
    RECT 0 2.136 0.024 2.160 ;
    RECT 0 2.184 0.024 2.208 ;
    RECT 0 2.232 0.024 3.072 ;
    RECT 0 3.096 0.024 3.120 ;
    RECT 0 3.144 0.024 3.168 ;
    RECT 0 3.192 0.024 3.216 ;
    RECT 0 3.240 0.024 3.264 ;
    RECT 0 3.288 0.024 3.312 ;
    RECT 0 3.336 0.024 3.360 ;
    RECT 0 3.384 0.024 3.408 ;
    RECT 0 3.432 0.024 3.456 ;
    RECT 0 3.480 0.024 3.504 ;
    RECT 0 3.528 0.024 3.552 ;
    RECT 0 3.576 0.024 3.600 ;
    RECT 0 3.624 0.024 3.648 ;
    RECT 0 3.672 0.024 3.696 ;
    RECT 0 3.720 0.024 3.744 ;
    RECT 0 3.768 0.024 3.792 ;
    RECT 0 3.816 0.024 3.840 ;
    RECT 0 3.864 0.024 3.888 ;
    RECT 0 3.912 0.024 3.936 ;
    RECT 0 3.960 0.024 3.984 ;
    RECT 0 4.008 0.024 4.032 ;
    RECT 0 4.056 0.024 4.080 ;
    RECT 0 4.104 0.024 4.128 ;
    RECT 0 4.152 0.024 4.176 ;
    RECT 0 4.200 0.024 4.224 ;
    RECT 0 4.248 0.024 4.272 ;
    RECT 0 4.296 0.024 4.320 ;
    RECT 0 4.344 0.024 4.368 ;
    RECT 0 4.392 0.024 4.416 ;
    RECT 0 4.440 0.024 4.464 ;
    RECT 0 4.488 0.024 4.512 ;
    RECT 0 4.536 0.024 4.560 ;
    RECT 0 4.584 0.024 4.608 ;
    RECT 0 4.632 0.024 4.656 ;
    RECT 0 4.680 0.024 4.704 ;
    RECT 0 4.728 0.024 4.752 ;
    RECT 0 4.776 0.024 4.800 ;
    RECT 0 4.824 0.024 4.848 ;
    RECT 0 4.872 0.024 4.896 ;
    RECT 0 4.920 0.024 4.944 ;
    RECT 0 4.968 0.024 4.992 ;
    RECT 0 5.016 0.024 5.040 ;
    RECT 0 5.064 0.024 5.088 ;
    RECT 0 5.112 0.024 5.136 ;
    RECT 0 5.160 0.024 5.184 ;
    RECT 0 5.208 0.024 5.232 ;
    RECT 0 5.256 0.024 6.096 ;
    RECT 0 6.120 0.024 6.144 ;
    RECT 0 6.168 0.024 6.192 ;
    RECT 0 6.216 0.024 6.240 ;
    RECT 0 6.264 0.024 6.288 ;
    RECT 0 6.312 0.024 6.336 ;
    RECT 0 6.360 0.024 6.384 ;
    RECT 0 6.408 0.024 6.432 ;
    RECT 0 6.456 0.024 6.480 ;
    RECT 0 6.504 0.024 6.528 ;
    RECT 0 6.552 0.024 6.576 ;
    RECT 0 6.600 0.024 6.624 ;
    RECT 0 6.648 0.024 6.672 ;
    RECT 0 6.696 0.024 6.720 ;
    RECT 0 6.744 0.024 6.768 ;
    RECT 0 6.792 0.024 6.816 ;
    RECT 0 6.840 0.024 6.864 ;
    RECT 0 6.888 0.024 6.912 ;
    RECT 0 6.936 0.024 6.960 ;
    RECT 0 6.984 0.024 7.008 ;
    RECT 0 7.032 0.024 7.056 ;
    RECT 0 7.080 0.024 7.104 ;
    RECT 0 7.128 0.024 7.152 ;
    RECT 0 7.176 0.024 7.200 ;
    RECT 0 7.224 0.024 7.248 ;
    RECT 0 7.272 0.024 7.296 ;
    RECT 0 7.320 0.024 7.344 ;
    RECT 0 7.368 0.024 7.392 ;
    RECT 0 7.416 0.024 7.440 ;
    RECT 0 7.464 0.024 7.488 ;
    RECT 0 7.512 0.024 7.536 ;
    RECT 0 7.560 0.024 7.584 ;
    RECT 0 7.608 0.024 7.632 ;
    RECT 0 7.656 0.024 7.680 ;
    RECT 0 7.704 0.024 7.728 ;
    RECT 0 7.752 0.024 7.776 ;
    RECT 0 7.800 0.024 7.824 ;
    RECT 0 7.848 0.024 7.872 ;
    RECT 0 7.896 0.024 7.920 ;
    RECT 0 7.944 0.024 7.968 ;
    RECT 0 7.992 0.024 8.016 ;
    RECT 0 8.040 0.024 8.064 ;
    RECT 0 8.088 0.024 8.112 ;
    RECT 0 8.136 0.024 8.160 ;
    RECT 0 8.184 0.024 8.208 ;
    RECT 0 8.232 0.024 8.256 ;
    RECT 0 8.280 0.024 9.120 ;
    RECT 0 9.144 0.024 9.168 ;
    RECT 0 9.192 0.024 9.216 ;
    RECT 0 9.240 0.024 9.264 ;
    RECT 0 9.288 0.024 9.312 ;
    RECT 0 9.336 0.024 10.176 ;
    RECT 0 10.200 0.024 10.224 ;
    RECT 0 10.248 0.024 10.272 ;
    RECT 0 10.296 0.024 8.400 ;
#    LAYER OVERLAP ;
#    RECT 0 0 6.080 8.400 ;
  END
END fakeram_32x46

END LIBRARY
