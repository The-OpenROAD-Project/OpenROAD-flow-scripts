VERSION 5.7 ;
BUSBITCHARS "[]" ;
MACRO fakeram45_256x16
  FOREIGN fakeram45_256x16 0 0 ;
  SYMMETRY X Y R90 ;
  SIZE 77.710 BY 40.600 ;
  CLASS BLOCK ;
  PIN w_mask_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.400 0.070 1.470 ;
    END
  END w_mask_in[0]
  PIN w_mask_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 1.960 0.070 2.030 ;
    END
  END w_mask_in[1]
  PIN w_mask_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 2.520 0.070 2.590 ;
    END
  END w_mask_in[2]
  PIN w_mask_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.080 0.070 3.150 ;
    END
  END w_mask_in[3]
  PIN w_mask_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 3.640 0.070 3.710 ;
    END
  END w_mask_in[4]
  PIN w_mask_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.200 0.070 4.270 ;
    END
  END w_mask_in[5]
  PIN w_mask_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 4.760 0.070 4.830 ;
    END
  END w_mask_in[6]
  PIN w_mask_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.320 0.070 5.390 ;
    END
  END w_mask_in[7]
  PIN w_mask_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 5.880 0.070 5.950 ;
    END
  END w_mask_in[8]
  PIN w_mask_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 6.440 0.070 6.510 ;
    END
  END w_mask_in[9]
  PIN w_mask_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.000 0.070 7.070 ;
    END
  END w_mask_in[10]
  PIN w_mask_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 7.560 0.070 7.630 ;
    END
  END w_mask_in[11]
  PIN w_mask_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.120 0.070 8.190 ;
    END
  END w_mask_in[12]
  PIN w_mask_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 8.680 0.070 8.750 ;
    END
  END w_mask_in[13]
  PIN w_mask_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.240 0.070 9.310 ;
    END
  END w_mask_in[14]
  PIN w_mask_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 9.800 0.070 9.870 ;
    END
  END w_mask_in[15]
  PIN rd_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 10.920 0.070 10.990 ;
    END
  END rd_out[0]
  PIN rd_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 11.480 0.070 11.550 ;
    END
  END rd_out[1]
  PIN rd_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.040 0.070 12.110 ;
    END
  END rd_out[2]
  PIN rd_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 12.600 0.070 12.670 ;
    END
  END rd_out[3]
  PIN rd_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.160 0.070 13.230 ;
    END
  END rd_out[4]
  PIN rd_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 13.720 0.070 13.790 ;
    END
  END rd_out[5]
  PIN rd_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.280 0.070 14.350 ;
    END
  END rd_out[6]
  PIN rd_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 14.840 0.070 14.910 ;
    END
  END rd_out[7]
  PIN rd_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.400 0.070 15.470 ;
    END
  END rd_out[8]
  PIN rd_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 15.960 0.070 16.030 ;
    END
  END rd_out[9]
  PIN rd_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 16.520 0.070 16.590 ;
    END
  END rd_out[10]
  PIN rd_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.080 0.070 17.150 ;
    END
  END rd_out[11]
  PIN rd_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 17.640 0.070 17.710 ;
    END
  END rd_out[12]
  PIN rd_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.200 0.070 18.270 ;
    END
  END rd_out[13]
  PIN rd_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 18.760 0.070 18.830 ;
    END
  END rd_out[14]
  PIN rd_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 19.320 0.070 19.390 ;
    END
  END rd_out[15]
  PIN wd_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 20.440 0.070 20.510 ;
    END
  END wd_in[0]
  PIN wd_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.000 0.070 21.070 ;
    END
  END wd_in[1]
  PIN wd_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 21.560 0.070 21.630 ;
    END
  END wd_in[2]
  PIN wd_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.120 0.070 22.190 ;
    END
  END wd_in[3]
  PIN wd_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 22.680 0.070 22.750 ;
    END
  END wd_in[4]
  PIN wd_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.240 0.070 23.310 ;
    END
  END wd_in[5]
  PIN wd_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 23.800 0.070 23.870 ;
    END
  END wd_in[6]
  PIN wd_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.360 0.070 24.430 ;
    END
  END wd_in[7]
  PIN wd_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 24.920 0.070 24.990 ;
    END
  END wd_in[8]
  PIN wd_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 25.480 0.070 25.550 ;
    END
  END wd_in[9]
  PIN wd_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.040 0.070 26.110 ;
    END
  END wd_in[10]
  PIN wd_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 26.600 0.070 26.670 ;
    END
  END wd_in[11]
  PIN wd_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.160 0.070 27.230 ;
    END
  END wd_in[12]
  PIN wd_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 27.720 0.070 27.790 ;
    END
  END wd_in[13]
  PIN wd_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.280 0.070 28.350 ;
    END
  END wd_in[14]
  PIN wd_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 28.840 0.070 28.910 ;
    END
  END wd_in[15]
  PIN addr_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 29.960 0.070 30.030 ;
    END
  END addr_in[0]
  PIN addr_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 30.520 0.070 30.590 ;
    END
  END addr_in[1]
  PIN addr_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.080 0.070 31.150 ;
    END
  END addr_in[2]
  PIN addr_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 31.640 0.070 31.710 ;
    END
  END addr_in[3]
  PIN addr_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.200 0.070 32.270 ;
    END
  END addr_in[4]
  PIN addr_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 32.760 0.070 32.830 ;
    END
  END addr_in[5]
  PIN addr_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.320 0.070 33.390 ;
    END
  END addr_in[6]
  PIN addr_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 33.880 0.070 33.950 ;
    END
  END addr_in[7]
  PIN we_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.000 0.070 35.070 ;
    END
  END we_in
  PIN ce_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 35.560 0.070 35.630 ;
    END
  END ce_in
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal3 ;
      RECT 0.000 36.120 0.070 36.190 ;
    END
  END clk
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER metal4 ;
      RECT 1.260 1.400 1.540 39.200 ;
      RECT 3.500 1.400 3.780 39.200 ;
      RECT 5.740 1.400 6.020 39.200 ;
      RECT 7.980 1.400 8.260 39.200 ;
      RECT 10.220 1.400 10.500 39.200 ;
      RECT 12.460 1.400 12.740 39.200 ;
      RECT 14.700 1.400 14.980 39.200 ;
      RECT 16.940 1.400 17.220 39.200 ;
      RECT 19.180 1.400 19.460 39.200 ;
      RECT 21.420 1.400 21.700 39.200 ;
      RECT 23.660 1.400 23.940 39.200 ;
      RECT 25.900 1.400 26.180 39.200 ;
      RECT 28.140 1.400 28.420 39.200 ;
      RECT 30.380 1.400 30.660 39.200 ;
      RECT 32.620 1.400 32.900 39.200 ;
      RECT 34.860 1.400 35.140 39.200 ;
      RECT 37.100 1.400 37.380 39.200 ;
      RECT 39.340 1.400 39.620 39.200 ;
      RECT 41.580 1.400 41.860 39.200 ;
      RECT 43.820 1.400 44.100 39.200 ;
      RECT 46.060 1.400 46.340 39.200 ;
      RECT 48.300 1.400 48.580 39.200 ;
      RECT 50.540 1.400 50.820 39.200 ;
      RECT 52.780 1.400 53.060 39.200 ;
      RECT 55.020 1.400 55.300 39.200 ;
      RECT 57.260 1.400 57.540 39.200 ;
      RECT 59.500 1.400 59.780 39.200 ;
      RECT 61.740 1.400 62.020 39.200 ;
      RECT 63.980 1.400 64.260 39.200 ;
      RECT 66.220 1.400 66.500 39.200 ;
      RECT 68.460 1.400 68.740 39.200 ;
      RECT 70.700 1.400 70.980 39.200 ;
      RECT 72.940 1.400 73.220 39.200 ;
      RECT 75.180 1.400 75.460 39.200 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER metal4 ;
      RECT 2.380 1.400 2.660 39.200 ;
      RECT 4.620 1.400 4.900 39.200 ;
      RECT 6.860 1.400 7.140 39.200 ;
      RECT 9.100 1.400 9.380 39.200 ;
      RECT 11.340 1.400 11.620 39.200 ;
      RECT 13.580 1.400 13.860 39.200 ;
      RECT 15.820 1.400 16.100 39.200 ;
      RECT 18.060 1.400 18.340 39.200 ;
      RECT 20.300 1.400 20.580 39.200 ;
      RECT 22.540 1.400 22.820 39.200 ;
      RECT 24.780 1.400 25.060 39.200 ;
      RECT 27.020 1.400 27.300 39.200 ;
      RECT 29.260 1.400 29.540 39.200 ;
      RECT 31.500 1.400 31.780 39.200 ;
      RECT 33.740 1.400 34.020 39.200 ;
      RECT 35.980 1.400 36.260 39.200 ;
      RECT 38.220 1.400 38.500 39.200 ;
      RECT 40.460 1.400 40.740 39.200 ;
      RECT 42.700 1.400 42.980 39.200 ;
      RECT 44.940 1.400 45.220 39.200 ;
      RECT 47.180 1.400 47.460 39.200 ;
      RECT 49.420 1.400 49.700 39.200 ;
      RECT 51.660 1.400 51.940 39.200 ;
      RECT 53.900 1.400 54.180 39.200 ;
      RECT 56.140 1.400 56.420 39.200 ;
      RECT 58.380 1.400 58.660 39.200 ;
      RECT 60.620 1.400 60.900 39.200 ;
      RECT 62.860 1.400 63.140 39.200 ;
      RECT 65.100 1.400 65.380 39.200 ;
      RECT 67.340 1.400 67.620 39.200 ;
      RECT 69.580 1.400 69.860 39.200 ;
      RECT 71.820 1.400 72.100 39.200 ;
      RECT 74.060 1.400 74.340 39.200 ;
    END
  END VDD
  OBS
    LAYER metal1 ;
    RECT 0 0 77.710 40.600 ;
    LAYER metal2 ;
    RECT 0 0 77.710 40.600 ;
    LAYER metal3 ;
    RECT 0.070 0 77.710 40.600 ;
    RECT 0 0.000 0.070 1.400 ;
    RECT 0 1.470 0.070 1.960 ;
    RECT 0 2.030 0.070 2.520 ;
    RECT 0 2.590 0.070 3.080 ;
    RECT 0 3.150 0.070 3.640 ;
    RECT 0 3.710 0.070 4.200 ;
    RECT 0 4.270 0.070 4.760 ;
    RECT 0 4.830 0.070 5.320 ;
    RECT 0 5.390 0.070 5.880 ;
    RECT 0 5.950 0.070 6.440 ;
    RECT 0 6.510 0.070 7.000 ;
    RECT 0 7.070 0.070 7.560 ;
    RECT 0 7.630 0.070 8.120 ;
    RECT 0 8.190 0.070 8.680 ;
    RECT 0 8.750 0.070 9.240 ;
    RECT 0 9.310 0.070 9.800 ;
    RECT 0 9.870 0.070 10.920 ;
    RECT 0 10.990 0.070 11.480 ;
    RECT 0 11.550 0.070 12.040 ;
    RECT 0 12.110 0.070 12.600 ;
    RECT 0 12.670 0.070 13.160 ;
    RECT 0 13.230 0.070 13.720 ;
    RECT 0 13.790 0.070 14.280 ;
    RECT 0 14.350 0.070 14.840 ;
    RECT 0 14.910 0.070 15.400 ;
    RECT 0 15.470 0.070 15.960 ;
    RECT 0 16.030 0.070 16.520 ;
    RECT 0 16.590 0.070 17.080 ;
    RECT 0 17.150 0.070 17.640 ;
    RECT 0 17.710 0.070 18.200 ;
    RECT 0 18.270 0.070 18.760 ;
    RECT 0 18.830 0.070 19.320 ;
    RECT 0 19.390 0.070 20.440 ;
    RECT 0 20.510 0.070 21.000 ;
    RECT 0 21.070 0.070 21.560 ;
    RECT 0 21.630 0.070 22.120 ;
    RECT 0 22.190 0.070 22.680 ;
    RECT 0 22.750 0.070 23.240 ;
    RECT 0 23.310 0.070 23.800 ;
    RECT 0 23.870 0.070 24.360 ;
    RECT 0 24.430 0.070 24.920 ;
    RECT 0 24.990 0.070 25.480 ;
    RECT 0 25.550 0.070 26.040 ;
    RECT 0 26.110 0.070 26.600 ;
    RECT 0 26.670 0.070 27.160 ;
    RECT 0 27.230 0.070 27.720 ;
    RECT 0 27.790 0.070 28.280 ;
    RECT 0 28.350 0.070 28.840 ;
    RECT 0 28.910 0.070 29.960 ;
    RECT 0 30.030 0.070 30.520 ;
    RECT 0 30.590 0.070 31.080 ;
    RECT 0 31.150 0.070 31.640 ;
    RECT 0 31.710 0.070 32.200 ;
    RECT 0 32.270 0.070 32.760 ;
    RECT 0 32.830 0.070 33.320 ;
    RECT 0 33.390 0.070 33.880 ;
    RECT 0 33.950 0.070 35.000 ;
    RECT 0 35.070 0.070 35.560 ;
    RECT 0 35.630 0.070 36.120 ;
    RECT 0 36.190 0.070 40.600 ;
    LAYER metal4 ;
    RECT 0 0 77.710 1.400 ;
    RECT 0 39.200 77.710 40.600 ;
    RECT 0.000 1.400 1.260 39.200 ;
    RECT 1.540 1.400 2.380 39.200 ;
    RECT 2.660 1.400 3.500 39.200 ;
    RECT 3.780 1.400 4.620 39.200 ;
    RECT 4.900 1.400 5.740 39.200 ;
    RECT 6.020 1.400 6.860 39.200 ;
    RECT 7.140 1.400 7.980 39.200 ;
    RECT 8.260 1.400 9.100 39.200 ;
    RECT 9.380 1.400 10.220 39.200 ;
    RECT 10.500 1.400 11.340 39.200 ;
    RECT 11.620 1.400 12.460 39.200 ;
    RECT 12.740 1.400 13.580 39.200 ;
    RECT 13.860 1.400 14.700 39.200 ;
    RECT 14.980 1.400 15.820 39.200 ;
    RECT 16.100 1.400 16.940 39.200 ;
    RECT 17.220 1.400 18.060 39.200 ;
    RECT 18.340 1.400 19.180 39.200 ;
    RECT 19.460 1.400 20.300 39.200 ;
    RECT 20.580 1.400 21.420 39.200 ;
    RECT 21.700 1.400 22.540 39.200 ;
    RECT 22.820 1.400 23.660 39.200 ;
    RECT 23.940 1.400 24.780 39.200 ;
    RECT 25.060 1.400 25.900 39.200 ;
    RECT 26.180 1.400 27.020 39.200 ;
    RECT 27.300 1.400 28.140 39.200 ;
    RECT 28.420 1.400 29.260 39.200 ;
    RECT 29.540 1.400 30.380 39.200 ;
    RECT 30.660 1.400 31.500 39.200 ;
    RECT 31.780 1.400 32.620 39.200 ;
    RECT 32.900 1.400 33.740 39.200 ;
    RECT 34.020 1.400 34.860 39.200 ;
    RECT 35.140 1.400 35.980 39.200 ;
    RECT 36.260 1.400 37.100 39.200 ;
    RECT 37.380 1.400 38.220 39.200 ;
    RECT 38.500 1.400 39.340 39.200 ;
    RECT 39.620 1.400 40.460 39.200 ;
    RECT 40.740 1.400 41.580 39.200 ;
    RECT 41.860 1.400 42.700 39.200 ;
    RECT 42.980 1.400 43.820 39.200 ;
    RECT 44.100 1.400 44.940 39.200 ;
    RECT 45.220 1.400 46.060 39.200 ;
    RECT 46.340 1.400 47.180 39.200 ;
    RECT 47.460 1.400 48.300 39.200 ;
    RECT 48.580 1.400 49.420 39.200 ;
    RECT 49.700 1.400 50.540 39.200 ;
    RECT 50.820 1.400 51.660 39.200 ;
    RECT 51.940 1.400 52.780 39.200 ;
    RECT 53.060 1.400 53.900 39.200 ;
    RECT 54.180 1.400 55.020 39.200 ;
    RECT 55.300 1.400 56.140 39.200 ;
    RECT 56.420 1.400 57.260 39.200 ;
    RECT 57.540 1.400 58.380 39.200 ;
    RECT 58.660 1.400 59.500 39.200 ;
    RECT 59.780 1.400 60.620 39.200 ;
    RECT 60.900 1.400 61.740 39.200 ;
    RECT 62.020 1.400 62.860 39.200 ;
    RECT 63.140 1.400 63.980 39.200 ;
    RECT 64.260 1.400 65.100 39.200 ;
    RECT 65.380 1.400 66.220 39.200 ;
    RECT 66.500 1.400 67.340 39.200 ;
    RECT 67.620 1.400 68.460 39.200 ;
    RECT 68.740 1.400 69.580 39.200 ;
    RECT 69.860 1.400 70.700 39.200 ;
    RECT 70.980 1.400 71.820 39.200 ;
    RECT 72.100 1.400 72.940 39.200 ;
    RECT 73.220 1.400 74.060 39.200 ;
    RECT 74.340 1.400 75.180 39.200 ;
    RECT 75.460 1.400 77.710 39.200 ;
    LAYER OVERLAP ;
    RECT 0 0 77.710 40.600 ;
  END
END fakeram45_256x16

END LIBRARY
