VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DFHV2Xx1_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx1_ASAP7_75t_L 0 0 ;
  SIZE 1.242 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.224 0.243 ;
        RECT 1.206 0.027 1.224 0.243 ;
        RECT 1.174 0.027 1.224 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.224 0.513 ;
        RECT 1.206 0.297 1.224 0.513 ;
        RECT 1.174 0.297 1.224 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.242 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.242 0.009 ;
        RECT 0 0.531 1.242 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.242 0.008 ;
      RECT 0 0.262 1.242 0.278 ;
      RECT 0 0.532 1.242 0.548 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.175 0.162 ;
      RECT 0.936 0.378 1.175 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx1_ASAP7_75t_L

MACRO DFHV2Xx1_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx1_ASAP7_75t_R 0 0 ;
  SIZE 1.242 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.224 0.243 ;
        RECT 1.206 0.027 1.224 0.243 ;
        RECT 1.174 0.027 1.224 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.224 0.513 ;
        RECT 1.206 0.297 1.224 0.513 ;
        RECT 1.174 0.297 1.224 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.242 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.242 0.009 ;
        RECT 0 0.531 1.242 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.242 0.008 ;
      RECT 0 0.262 1.242 0.278 ;
      RECT 0 0.532 1.242 0.548 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.175 0.162 ;
      RECT 0.936 0.378 1.175 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx1_ASAP7_75t_R

MACRO DFHV2Xx1_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx1_ASAP7_75t_SL 0 0 ;
  SIZE 1.242 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.224 0.243 ;
        RECT 1.206 0.027 1.224 0.243 ;
        RECT 1.174 0.027 1.224 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.224 0.513 ;
        RECT 1.206 0.297 1.224 0.513 ;
        RECT 1.174 0.297 1.224 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.242 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.242 0.009 ;
        RECT 0 0.531 1.242 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.242 0.008 ;
      RECT 0 0.262 1.242 0.278 ;
      RECT 0 0.532 1.242 0.548 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.175 0.162 ;
      RECT 0.936 0.378 1.175 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx1_ASAP7_75t_SL

MACRO DFHV2Xx2_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx2_ASAP7_75t_L 0 0 ;
  SIZE 1.296 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.278 0.243 ;
        RECT 1.26 0.027 1.278 0.243 ;
        RECT 1.174 0.027 1.278 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.278 0.513 ;
        RECT 1.26 0.297 1.278 0.513 ;
        RECT 1.174 0.297 1.278 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.296 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.296 0.009 ;
        RECT 0 0.531 1.296 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.296 0.008 ;
      RECT 0 0.262 1.296 0.278 ;
      RECT 0 0.532 1.296 0.548 ;
      RECT 1.203 0.125 1.227 0.147 ;
      RECT 1.203 0.393 1.227 0.415 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.206 0.101 1.224 0.167 ;
      RECT 1.206 0.373 1.224 0.439 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.229 0.162 ;
      RECT 0.936 0.378 1.229 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.206 0.144 1.224 0.162 ;
      RECT 1.206 0.378 1.224 0.396 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx2_ASAP7_75t_L

MACRO DFHV2Xx2_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx2_ASAP7_75t_R 0 0 ;
  SIZE 1.296 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.278 0.243 ;
        RECT 1.26 0.027 1.278 0.243 ;
        RECT 1.174 0.027 1.278 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.278 0.513 ;
        RECT 1.26 0.297 1.278 0.513 ;
        RECT 1.174 0.297 1.278 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.296 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.296 0.009 ;
        RECT 0 0.531 1.296 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.296 0.008 ;
      RECT 0 0.262 1.296 0.278 ;
      RECT 0 0.532 1.296 0.548 ;
      RECT 1.203 0.125 1.227 0.147 ;
      RECT 1.203 0.393 1.227 0.415 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.206 0.101 1.224 0.167 ;
      RECT 1.206 0.373 1.224 0.439 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.229 0.162 ;
      RECT 0.936 0.378 1.229 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.206 0.144 1.224 0.162 ;
      RECT 1.206 0.378 1.224 0.396 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx2_ASAP7_75t_R

MACRO DFHV2Xx2_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx2_ASAP7_75t_SL 0 0 ;
  SIZE 1.296 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.278 0.243 ;
        RECT 1.26 0.027 1.278 0.243 ;
        RECT 1.174 0.027 1.278 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.278 0.513 ;
        RECT 1.26 0.297 1.278 0.513 ;
        RECT 1.174 0.297 1.278 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.296 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.296 0.009 ;
        RECT 0 0.531 1.296 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.296 0.008 ;
      RECT 0 0.262 1.296 0.278 ;
      RECT 0 0.532 1.296 0.548 ;
      RECT 1.203 0.125 1.227 0.147 ;
      RECT 1.203 0.393 1.227 0.415 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.206 0.101 1.224 0.167 ;
      RECT 1.206 0.373 1.224 0.439 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.229 0.162 ;
      RECT 0.936 0.378 1.229 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.206 0.144 1.224 0.162 ;
      RECT 1.206 0.378 1.224 0.396 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx2_ASAP7_75t_SL

MACRO DFHV2Xx3_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx3_ASAP7_75t_L 0 0 ;
  SIZE 1.35 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.332 0.243 ;
        RECT 1.314 0.027 1.332 0.243 ;
        RECT 1.174 0.027 1.332 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.332 0.513 ;
        RECT 1.314 0.297 1.332 0.513 ;
        RECT 1.174 0.297 1.332 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.35 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.35 0.009 ;
        RECT 0 0.531 1.35 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.35 0.008 ;
      RECT 0 0.262 1.35 0.278 ;
      RECT 0 0.532 1.35 0.548 ;
      RECT 1.257 0.125 1.281 0.147 ;
      RECT 1.257 0.393 1.281 0.415 ;
      RECT 1.203 0.125 1.227 0.147 ;
      RECT 1.203 0.393 1.227 0.415 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.26 0.101 1.278 0.167 ;
      RECT 1.26 0.373 1.278 0.439 ;
      RECT 1.206 0.101 1.224 0.167 ;
      RECT 1.206 0.373 1.224 0.439 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.283 0.162 ;
      RECT 0.936 0.378 1.283 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.26 0.378 1.278 0.396 ;
      RECT 1.206 0.144 1.224 0.162 ;
      RECT 1.206 0.378 1.224 0.396 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx3_ASAP7_75t_L

MACRO DFHV2Xx3_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx3_ASAP7_75t_R 0 0 ;
  SIZE 1.35 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.332 0.243 ;
        RECT 1.314 0.027 1.332 0.243 ;
        RECT 1.174 0.027 1.332 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.332 0.513 ;
        RECT 1.314 0.297 1.332 0.513 ;
        RECT 1.174 0.297 1.332 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.35 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.35 0.009 ;
        RECT 0 0.531 1.35 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.35 0.008 ;
      RECT 0 0.262 1.35 0.278 ;
      RECT 0 0.532 1.35 0.548 ;
      RECT 1.257 0.125 1.281 0.147 ;
      RECT 1.257 0.393 1.281 0.415 ;
      RECT 1.203 0.125 1.227 0.147 ;
      RECT 1.203 0.393 1.227 0.415 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.26 0.101 1.278 0.167 ;
      RECT 1.26 0.373 1.278 0.439 ;
      RECT 1.206 0.101 1.224 0.167 ;
      RECT 1.206 0.373 1.224 0.439 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.283 0.162 ;
      RECT 0.936 0.378 1.283 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.26 0.378 1.278 0.396 ;
      RECT 1.206 0.144 1.224 0.162 ;
      RECT 1.206 0.378 1.224 0.396 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx3_ASAP7_75t_R

MACRO DFHV2Xx3_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx3_ASAP7_75t_SL 0 0 ;
  SIZE 1.35 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.332 0.243 ;
        RECT 1.314 0.027 1.332 0.243 ;
        RECT 1.174 0.027 1.332 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.332 0.513 ;
        RECT 1.314 0.297 1.332 0.513 ;
        RECT 1.174 0.297 1.332 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.35 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.35 0.009 ;
        RECT 0 0.531 1.35 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.35 0.008 ;
      RECT 0 0.262 1.35 0.278 ;
      RECT 0 0.532 1.35 0.548 ;
      RECT 1.257 0.125 1.281 0.147 ;
      RECT 1.257 0.393 1.281 0.415 ;
      RECT 1.203 0.125 1.227 0.147 ;
      RECT 1.203 0.393 1.227 0.415 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.26 0.101 1.278 0.167 ;
      RECT 1.26 0.373 1.278 0.439 ;
      RECT 1.206 0.101 1.224 0.167 ;
      RECT 1.206 0.373 1.224 0.439 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.283 0.162 ;
      RECT 0.936 0.378 1.283 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.26 0.378 1.278 0.396 ;
      RECT 1.206 0.144 1.224 0.162 ;
      RECT 1.206 0.378 1.224 0.396 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx3_ASAP7_75t_SL

MACRO DFHV2Xx4_ASAP7_75t_L
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx4_ASAP7_75t_L 0 0 ;
  SIZE 1.404 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.386 0.243 ;
        RECT 1.368 0.027 1.386 0.243 ;
        RECT 1.174 0.027 1.386 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.386 0.513 ;
        RECT 1.368 0.297 1.386 0.513 ;
        RECT 1.174 0.297 1.386 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.404 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
        RECT 0 0.531 1.404 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.404 0.008 ;
      RECT 0 0.262 1.404 0.278 ;
      RECT 0 0.532 1.404 0.548 ;
      RECT 1.311 0.125 1.335 0.147 ;
      RECT 1.311 0.393 1.335 0.415 ;
      RECT 1.257 0.125 1.281 0.147 ;
      RECT 1.257 0.393 1.281 0.415 ;
      RECT 1.203 0.125 1.227 0.147 ;
      RECT 1.203 0.393 1.227 0.415 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.314 0.101 1.332 0.167 ;
      RECT 1.314 0.373 1.332 0.439 ;
      RECT 1.26 0.101 1.278 0.167 ;
      RECT 1.26 0.373 1.278 0.439 ;
      RECT 1.206 0.101 1.224 0.167 ;
      RECT 1.206 0.373 1.224 0.439 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.337 0.162 ;
      RECT 0.936 0.378 1.337 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.314 0.144 1.332 0.162 ;
      RECT 1.314 0.378 1.332 0.396 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.26 0.378 1.278 0.396 ;
      RECT 1.206 0.144 1.224 0.162 ;
      RECT 1.206 0.378 1.224 0.396 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx4_ASAP7_75t_L

MACRO DFHV2Xx4_ASAP7_75t_R
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx4_ASAP7_75t_R 0 0 ;
  SIZE 1.404 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.386 0.243 ;
        RECT 1.368 0.027 1.386 0.243 ;
        RECT 1.174 0.027 1.386 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.386 0.513 ;
        RECT 1.368 0.297 1.386 0.513 ;
        RECT 1.174 0.297 1.386 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.404 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
        RECT 0 0.531 1.404 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.404 0.008 ;
      RECT 0 0.262 1.404 0.278 ;
      RECT 0 0.532 1.404 0.548 ;
      RECT 1.311 0.125 1.335 0.147 ;
      RECT 1.311 0.393 1.335 0.415 ;
      RECT 1.257 0.125 1.281 0.147 ;
      RECT 1.257 0.393 1.281 0.415 ;
      RECT 1.203 0.125 1.227 0.147 ;
      RECT 1.203 0.393 1.227 0.415 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.314 0.101 1.332 0.167 ;
      RECT 1.314 0.373 1.332 0.439 ;
      RECT 1.26 0.101 1.278 0.167 ;
      RECT 1.26 0.373 1.278 0.439 ;
      RECT 1.206 0.101 1.224 0.167 ;
      RECT 1.206 0.373 1.224 0.439 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.337 0.162 ;
      RECT 0.936 0.378 1.337 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.314 0.144 1.332 0.162 ;
      RECT 1.314 0.378 1.332 0.396 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.26 0.378 1.278 0.396 ;
      RECT 1.206 0.144 1.224 0.162 ;
      RECT 1.206 0.378 1.224 0.396 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx4_ASAP7_75t_R

MACRO DFHV2Xx4_ASAP7_75t_SL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFHV2Xx4_ASAP7_75t_SL 0 0 ;
  SIZE 1.404 BY 0.54 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.099 0.185 0.117 0.236 ;
        RECT 0.072 0.081 0.117 0.099 ;
        RECT 0.099 0.034 0.117 0.099 ;
        RECT 0.072 0.185 0.117 0.203 ;
        RECT 0.072 0.081 0.09 0.203 ;
    END
  END CLK
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.225 1.386 0.243 ;
        RECT 1.368 0.027 1.386 0.243 ;
        RECT 1.174 0.027 1.386 0.045 ;
    END
  END QN0
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.174 0.495 1.386 0.513 ;
        RECT 1.368 0.297 1.386 0.513 ;
        RECT 1.174 0.297 1.386 0.315 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 0.261 1.404 0.279 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.009 1.404 0.009 ;
        RECT 0 0.531 1.404 0.549 ;
    END
  END VSS
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.108 0.436 0.126 ;
      LAYER M1 ;
        RECT 0.396 0.106 0.414 0.164 ;
      LAYER V1 ;
        RECT 0.396 0.108 0.414 0.126 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.284 0.414 0.436 0.432 ;
      LAYER M1 ;
        RECT 0.396 0.376 0.414 0.434 ;
      LAYER V1 ;
        RECT 0.396 0.414 0.414 0.432 ;
    END
  END D1
  OBS
    LAYER LIG ;
      RECT 0 -0.008 1.404 0.008 ;
      RECT 0 0.262 1.404 0.278 ;
      RECT 0 0.532 1.404 0.548 ;
      RECT 1.311 0.125 1.335 0.147 ;
      RECT 1.311 0.393 1.335 0.415 ;
      RECT 1.257 0.125 1.281 0.147 ;
      RECT 1.257 0.393 1.281 0.415 ;
      RECT 1.203 0.125 1.227 0.147 ;
      RECT 1.203 0.393 1.227 0.415 ;
      RECT 1.149 0.125 1.173 0.147 ;
      RECT 1.149 0.393 1.173 0.415 ;
      RECT 1.041 0.129 1.065 0.151 ;
      RECT 1.041 0.389 1.065 0.411 ;
      RECT 0.987 0.094 1.011 0.117 ;
      RECT 0.987 0.423 1.011 0.446 ;
      RECT 0.933 0.165 0.957 0.191 ;
      RECT 0.933 0.349 0.957 0.375 ;
      RECT 0.879 0.124 0.903 0.146 ;
      RECT 0.879 0.394 0.903 0.416 ;
      RECT 0.825 0.165 0.849 0.191 ;
      RECT 0.825 0.349 0.849 0.375 ;
      RECT 0.772 0.12 0.795 0.142 ;
      RECT 0.772 0.398 0.795 0.42 ;
      RECT 0.717 0.079 0.756 0.101 ;
      RECT 0.717 0.439 0.756 0.461 ;
      RECT 0.663 0.165 0.687 0.191 ;
      RECT 0.663 0.349 0.687 0.375 ;
      RECT 0.61 0.124 0.633 0.146 ;
      RECT 0.61 0.394 0.633 0.416 ;
      RECT 0.556 0.125 0.579 0.146 ;
      RECT 0.556 0.394 0.579 0.415 ;
      RECT 0.394 0.124 0.416 0.146 ;
      RECT 0.394 0.394 0.416 0.416 ;
      RECT 0.124 0.124 0.146 0.146 ;
      RECT 0.07 0.124 0.092 0.146 ;
    LAYER M1 ;
      RECT 1.066 0.225 1.116 0.243 ;
      RECT 1.098 0.027 1.116 0.243 ;
      RECT 0.99 0.027 1.008 0.119 ;
      RECT 0.99 0.027 1.116 0.045 ;
      RECT 0.99 0.495 1.116 0.513 ;
      RECT 1.098 0.297 1.116 0.513 ;
      RECT 0.99 0.421 1.008 0.513 ;
      RECT 1.066 0.297 1.116 0.315 ;
      RECT 0.904 0.225 0.954 0.243 ;
      RECT 0.936 0.027 0.954 0.243 ;
      RECT 0.936 0.153 1.062 0.171 ;
      RECT 1.044 0.117 1.062 0.171 ;
      RECT 0.85 0.027 0.954 0.045 ;
      RECT 0.85 0.495 0.954 0.513 ;
      RECT 0.936 0.297 0.954 0.513 ;
      RECT 1.044 0.369 1.062 0.423 ;
      RECT 0.936 0.369 1.062 0.387 ;
      RECT 0.904 0.297 0.954 0.315 ;
      RECT 0.792 0.225 0.846 0.243 ;
      RECT 0.828 0.081 0.846 0.243 ;
      RECT 0.72 0.081 0.846 0.099 ;
      RECT 0.801 0.045 0.819 0.099 ;
      RECT 0.72 0.062 0.738 0.099 ;
      RECT 0.801 0.441 0.819 0.495 ;
      RECT 0.72 0.441 0.738 0.478 ;
      RECT 0.72 0.441 0.846 0.459 ;
      RECT 0.828 0.297 0.846 0.459 ;
      RECT 0.792 0.297 0.846 0.315 ;
      RECT 0.58 0.225 0.702 0.243 ;
      RECT 0.684 0.027 0.702 0.243 ;
      RECT 0.684 0.122 0.797 0.14 ;
      RECT 0.634 0.027 0.702 0.045 ;
      RECT 0.634 0.495 0.702 0.513 ;
      RECT 0.684 0.297 0.702 0.513 ;
      RECT 0.684 0.4 0.797 0.418 ;
      RECT 0.58 0.297 0.702 0.315 ;
      RECT 0.612 0.153 0.649 0.171 ;
      RECT 0.612 0.106 0.63 0.171 ;
      RECT 0.612 0.369 0.63 0.434 ;
      RECT 0.612 0.369 0.649 0.387 ;
      RECT 0.558 0.189 0.595 0.207 ;
      RECT 0.558 0.106 0.576 0.207 ;
      RECT 0.558 0.333 0.576 0.434 ;
      RECT 0.558 0.333 0.595 0.351 ;
      RECT 0.261 0.081 0.306 0.099 ;
      RECT 0.288 0.027 0.306 0.099 ;
      RECT 0.288 0.027 0.5 0.045 ;
      RECT 0.288 0.495 0.5 0.513 ;
      RECT 0.288 0.441 0.306 0.513 ;
      RECT 0.261 0.441 0.306 0.459 ;
      RECT 0.148 0.225 0.198 0.243 ;
      RECT 0.18 0.027 0.198 0.243 ;
      RECT 0.148 0.027 0.198 0.045 ;
      RECT 0.018 0.225 0.068 0.243 ;
      RECT 0.018 0.027 0.036 0.243 ;
      RECT 0.018 0.027 0.068 0.045 ;
      RECT 1.314 0.101 1.332 0.167 ;
      RECT 1.314 0.373 1.332 0.439 ;
      RECT 1.26 0.101 1.278 0.167 ;
      RECT 1.26 0.373 1.278 0.439 ;
      RECT 1.206 0.101 1.224 0.167 ;
      RECT 1.206 0.373 1.224 0.439 ;
      RECT 1.152 0.09 1.17 0.2 ;
      RECT 1.152 0.34 1.17 0.45 ;
      RECT 0.882 0.101 0.9 0.167 ;
      RECT 0.882 0.373 0.9 0.439 ;
      RECT 0.72 0.165 0.738 0.207 ;
      RECT 0.72 0.333 0.738 0.375 ;
      RECT 0.418 0.063 0.609 0.081 ;
      RECT 0.418 0.459 0.609 0.477 ;
      RECT 0.255 0.225 0.5 0.243 ;
      RECT 0.255 0.297 0.5 0.315 ;
      RECT 0.309 0.189 0.447 0.207 ;
      RECT 0.309 0.333 0.447 0.351 ;
      RECT 0.126 0.121 0.144 0.167 ;
    LAYER M2 ;
      RECT 0.936 0.144 1.337 0.162 ;
      RECT 0.936 0.378 1.337 0.396 ;
      RECT 0.013 0.144 0.9 0.162 ;
      RECT 0.607 0.378 0.9 0.396 ;
      RECT 0.175 0.18 0.743 0.198 ;
      RECT 0.553 0.342 0.743 0.36 ;
    LAYER V1 ;
      RECT 1.314 0.144 1.332 0.162 ;
      RECT 1.314 0.378 1.332 0.396 ;
      RECT 1.26 0.144 1.278 0.162 ;
      RECT 1.26 0.378 1.278 0.396 ;
      RECT 1.206 0.144 1.224 0.162 ;
      RECT 1.206 0.378 1.224 0.396 ;
      RECT 1.152 0.144 1.17 0.162 ;
      RECT 1.152 0.378 1.17 0.396 ;
      RECT 0.936 0.144 0.954 0.162 ;
      RECT 0.936 0.378 0.954 0.396 ;
      RECT 0.882 0.144 0.9 0.162 ;
      RECT 0.882 0.378 0.9 0.396 ;
      RECT 0.72 0.18 0.738 0.198 ;
      RECT 0.72 0.342 0.738 0.36 ;
      RECT 0.612 0.144 0.63 0.162 ;
      RECT 0.612 0.378 0.63 0.396 ;
      RECT 0.558 0.18 0.576 0.198 ;
      RECT 0.558 0.342 0.576 0.36 ;
      RECT 0.18 0.18 0.198 0.198 ;
      RECT 0.126 0.144 0.144 0.162 ;
      RECT 0.018 0.144 0.036 0.162 ;
    LAYER V2 ;
      RECT 0.828 0.144 0.846 0.162 ;
      RECT 0.828 0.378 0.846 0.396 ;
      RECT 0.612 0.18 0.63 0.198 ;
      RECT 0.612 0.342 0.63 0.36 ;
    LAYER M3 ;
      RECT 0.828 0.139 0.846 0.401 ;
      RECT 0.612 0.175 0.63 0.365 ;
  END
END DFHV2Xx4_ASAP7_75t_SL

END LIBRARY
