../../../../platforms/asap7/lef/fakeram7_256x34.lef