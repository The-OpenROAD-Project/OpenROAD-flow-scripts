VERSION 5.8 ;

MACRO bondpad_70x70
  CLASS COVER ;
  ORIGIN 0 0 ;
  FOREIGN bondpad_70x70 0 0 ;
  SIZE 70.0 BY 70.0 ;
  SYMMETRY X Y R90 ;
  SITE sg13g2_ioSite ;
  PIN pad
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0 0 70.0 70.0 ;
      LAYER Metal3 ;
        RECT 0 0 70.0 70.0 ;
      LAYER Metal4 ;
        RECT 0 0 70.0 70.0 ;
      LAYER Metal5 ;
        RECT 0 0 70.0 70.0 ;
      LAYER TopMetal1 ;
        RECT 0 0 70.0 70.0 ;
      LAYER TopMetal2 ;
        RECT 0 0 70.0 70.0 ;
    END
  END pad

  OBS
    LAYER Metal1 ;
      RECT 0 0 70.0 70.0 ;
    LAYER Metal2 ;
      RECT 0 0 70.0 70.0 ;
    LAYER Metal3 ;
      RECT 0 0 70.0 70.0 ;
    LAYER Metal4 ;
      RECT 0 0 70.0 70.0 ;
    LAYER Metal5 ;
      RECT 0 0 70.0 70.0 ;
    LAYER TopMetal1 ;
      RECT 0 0 70.0 70.0 ;
    LAYER TopMetal2 ;
      RECT 0 0 70.0 70.0 ;
  END
END bondpad_70x70
