../../../platforms/nangate45/lef/fakeram45_256x96.lef