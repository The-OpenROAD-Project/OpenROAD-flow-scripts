../../nangate45/lef/fakeram45_256x34.lef